
module dff_203 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_202 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_185 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_186 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_187 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_188 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_189 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_190 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_191 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_192 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_193 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_194 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_195 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_196 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_197 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_169 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_170 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_171 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_172 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_173 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_174 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_175 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_176 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_177 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_178 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_179 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_180 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_181 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_182 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_183 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_184 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_161 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_162 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_163 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_164 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_165 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_166 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_167 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_168 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_201 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_200 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_199 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_198 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX2 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module memc_Size16_7 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n214, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1162), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1161), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1160), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1159), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1158), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1157), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1156), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1155), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1154), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1153), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1152), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1151), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1150), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1149), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1148), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1147), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1146), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1145), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1144), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1143), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1142), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1141), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1140), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1139), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1138), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1137), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1136), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1135), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1134), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1133), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1132), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1131), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1130), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1129), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1128), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1127), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1126), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1125), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1124), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1123), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1122), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1121), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1120), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1119), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1118), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1117), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1116), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1115), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1114), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1113), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1112), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1111), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1110), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1109), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1108), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1107), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1106), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1105), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1104), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1103), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1102), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1101), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1100), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1099), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1098), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1097), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1096), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1095), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1094), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1093), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1092), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1091), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1090), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1089), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1088), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1087), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1086), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1085), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1083), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1082), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1081), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1080), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1079), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1078), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1077), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1076), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1075), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1074), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1073), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1072), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1071), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1070), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1069), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1068), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1067), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1066), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1065), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1064), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1063), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1062), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1061), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1060), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1059), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1058), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1057), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1056), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1055), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1054), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1053), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1052), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1051), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1050), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1049), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1048), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1047), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1046), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1045), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1044), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1043), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1042), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1041), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1040), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1039), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1038), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1037), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1036), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1035), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1034), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1033), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1032), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1031), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1030), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1029), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1028), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1027), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1026), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1025), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1024), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1023), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1022), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1021), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1020), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1019), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1018), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1017), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1016), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1015), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1014), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1013), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1012), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1011), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1010), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1009), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1008), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1007), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1006), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1005), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1004), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1003), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1002), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1001), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1000), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n999), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n998), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n997), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n996), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n995), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n994), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n993), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n992), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n991), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n990), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n989), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n988), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n987), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n986), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n985), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n984), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n983), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n982), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n981), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n980), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n979), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n978), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n977), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n976), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n975), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n974), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n973), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n972), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n971), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n970), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n969), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n968), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n967), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n966), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n965), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n964), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n963), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n962), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n961), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n960), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n959), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n958), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n957), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n956), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n955), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n954), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n953), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n952), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n951), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n950), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n949), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n948), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n947), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n946), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n945), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n944), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n943), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n942), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n941), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n940), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n939), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n938), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n937), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n936), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n935), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n934), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n933), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n932), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n931), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n930), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n929), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n928), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n927), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n926), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n925), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n924), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n923), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n922), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n921), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n920), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n919), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n918), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n917), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n916), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n915), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n914), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n913), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n912), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n911), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n910), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n909), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n908), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n907), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n906), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n905), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n904), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n903), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n902), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n901), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n900), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n899), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n898), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n897), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n896), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n895), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n894), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n893), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n892), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n891), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n890), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n889), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n888), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n887), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n886), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n885), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n884), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n883), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n882), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n881), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n880), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n879), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n878), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n877), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n876), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n875), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n874), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n873), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n872), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n871), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n870), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n869), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n868), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n867), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n866), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n865), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n864), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n863), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n862), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n861), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n860), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n859), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n858), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n857), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n856), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n855), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n854), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n853), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n852), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n851), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n850), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n849), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n848), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n847), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n846), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n845), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n844), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n843), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n842), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n841), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n840), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n839), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n838), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n837), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n836), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n835), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n834), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n833), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n832), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n831), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n830), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n829), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n828), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n827), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n826), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n825), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n824), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n823), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n822), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n821), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n820), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n819), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n818), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n817), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n816), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n815), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n814), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n813), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n812), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n811), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n810), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n809), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n808), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n807), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n806), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n805), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n804), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n803), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n802), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n801), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n800), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n799), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n798), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n797), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n796), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n795), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n794), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n793), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n792), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n791), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n790), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n789), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n788), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n787), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n786), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n785), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n784), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n783), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n782), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n781), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n780), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n779), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n778), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n777), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n776), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n775), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n774), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n773), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n772), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n771), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n770), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n769), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n768), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n767), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n766), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n765), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n764), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n763), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n762), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n761), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n760), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n759), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n758), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n757), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n756), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n755), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n754), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n753), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n752), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n751), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n750), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n749), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n748), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n747), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n746), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n745), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n744), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n743), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n742), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n741), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n740), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n739), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n738), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n737), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n736), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n735), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n734), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n733), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n732), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n731), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n730), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n729), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n728), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n727), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n726), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n725), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n724), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n723), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n722), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n721), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n720), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n719), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n718), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n717), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n716), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n715), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n714), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n713), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n712), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n711), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n710), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n709), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n708), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n707), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n706), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n705), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n704), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n703), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n702), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n701), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n700), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n699), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n698), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n697), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n696), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n695), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n694), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n693), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n692), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n691), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n690), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n689), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n688), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n687), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n686), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n685), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n684), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n683), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n682), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n681), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n680), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n679), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n678), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n677), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n676), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n675), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n674), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n673), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n672), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n671), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n670), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n669), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n668), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n667), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n666), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n665), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n664), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n663), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n662), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n661), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n660), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n659), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n658), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n657), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n656), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n655), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n654), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n653), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n652), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n651), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n214) );
  INVX4 U2 ( .A(n66), .Y(n67) );
  INVX4 U3 ( .A(n64), .Y(n65) );
  INVX4 U4 ( .A(n16), .Y(n17) );
  INVX4 U5 ( .A(n14), .Y(n15) );
  INVX4 U6 ( .A(n12), .Y(n13) );
  INVX4 U7 ( .A(n62), .Y(n63) );
  INVX4 U8 ( .A(n58), .Y(n59) );
  INVX4 U9 ( .A(n56), .Y(n57) );
  INVX4 U10 ( .A(n54), .Y(n55) );
  INVX4 U11 ( .A(n50), .Y(n51) );
  INVX4 U12 ( .A(n48), .Y(n49) );
  INVX4 U13 ( .A(n24), .Y(n25) );
  INVX4 U14 ( .A(n44), .Y(n45) );
  INVX4 U15 ( .A(n42), .Y(n43) );
  INVX4 U16 ( .A(n40), .Y(n41) );
  INVX4 U17 ( .A(n38), .Y(n39) );
  INVX4 U18 ( .A(n36), .Y(n37) );
  INVX4 U19 ( .A(n34), .Y(n35) );
  INVX4 U20 ( .A(n32), .Y(n33) );
  INVX4 U21 ( .A(n30), .Y(n31) );
  INVX4 U22 ( .A(n28), .Y(n29) );
  INVX4 U23 ( .A(n26), .Y(n27) );
  INVX4 U24 ( .A(n20), .Y(n21) );
  INVX4 U25 ( .A(n18), .Y(n19) );
  INVX4 U26 ( .A(n60), .Y(n61) );
  INVX4 U27 ( .A(n71), .Y(n1309) );
  INVX4 U28 ( .A(n68), .Y(n69) );
  INVX4 U29 ( .A(n52), .Y(n53) );
  INVX4 U30 ( .A(n46), .Y(n47) );
  INVX4 U31 ( .A(n22), .Y(n23) );
  BUFX4 U32 ( .A(n97), .Y(n1242) );
  AND2X2 U33 ( .A(\data_in<7> ), .B(n1308), .Y(n96) );
  INVX1 U34 ( .A(n1193), .Y(n1182) );
  INVX1 U35 ( .A(n1193), .Y(n1183) );
  INVX2 U36 ( .A(n1193), .Y(n1184) );
  INVX1 U37 ( .A(n1181), .Y(n1185) );
  INVX1 U38 ( .A(n1181), .Y(n1186) );
  INVX2 U39 ( .A(n1181), .Y(n1187) );
  INVX1 U40 ( .A(n1180), .Y(n1188) );
  INVX1 U41 ( .A(n1180), .Y(n1189) );
  INVX2 U42 ( .A(n1180), .Y(n1190) );
  INVX2 U43 ( .A(n1181), .Y(n1191) );
  INVX2 U44 ( .A(n1180), .Y(n1192) );
  INVX1 U45 ( .A(n645), .Y(N32) );
  INVX1 U46 ( .A(n646), .Y(N31) );
  INVX1 U47 ( .A(n647), .Y(N30) );
  INVX1 U48 ( .A(n648), .Y(N29) );
  INVX1 U49 ( .A(n649), .Y(N28) );
  INVX1 U50 ( .A(n650), .Y(N27) );
  INVX1 U51 ( .A(n1163), .Y(N26) );
  INVX1 U52 ( .A(n1164), .Y(N25) );
  INVX1 U53 ( .A(n1165), .Y(N24) );
  INVX1 U54 ( .A(n1166), .Y(N23) );
  INVX1 U55 ( .A(n1167), .Y(N22) );
  INVX1 U56 ( .A(n1168), .Y(N21) );
  INVX1 U57 ( .A(n1169), .Y(N20) );
  INVX1 U58 ( .A(n1170), .Y(N19) );
  INVX1 U59 ( .A(n1171), .Y(N18) );
  INVX1 U60 ( .A(n1172), .Y(N17) );
  BUFX2 U61 ( .A(n107), .Y(n1246) );
  BUFX2 U62 ( .A(n109), .Y(n1248) );
  BUFX2 U63 ( .A(n111), .Y(n1250) );
  BUFX2 U64 ( .A(n113), .Y(n1252) );
  BUFX2 U65 ( .A(n115), .Y(n1254) );
  BUFX2 U66 ( .A(n117), .Y(n1256) );
  BUFX2 U67 ( .A(n119), .Y(n1258) );
  BUFX2 U68 ( .A(n121), .Y(n1261) );
  BUFX2 U69 ( .A(n123), .Y(n1263) );
  BUFX2 U70 ( .A(n125), .Y(n1265) );
  BUFX2 U71 ( .A(n127), .Y(n1267) );
  BUFX2 U72 ( .A(n129), .Y(n1269) );
  BUFX2 U73 ( .A(n131), .Y(n1271) );
  BUFX2 U74 ( .A(n133), .Y(n1273) );
  BUFX2 U75 ( .A(n135), .Y(n1276) );
  BUFX2 U76 ( .A(n137), .Y(n1278) );
  BUFX2 U77 ( .A(n139), .Y(n1280) );
  BUFX2 U78 ( .A(n141), .Y(n1282) );
  BUFX2 U79 ( .A(n143), .Y(n1284) );
  BUFX2 U80 ( .A(n145), .Y(n1286) );
  BUFX2 U81 ( .A(n147), .Y(n1288) );
  BUFX2 U82 ( .A(n149), .Y(n1291) );
  BUFX2 U83 ( .A(n151), .Y(n1293) );
  BUFX2 U84 ( .A(n153), .Y(n1295) );
  BUFX2 U85 ( .A(n155), .Y(n1297) );
  BUFX2 U86 ( .A(n157), .Y(n1299) );
  BUFX2 U87 ( .A(n159), .Y(n1301) );
  BUFX2 U88 ( .A(n161), .Y(n1303) );
  INVX4 U89 ( .A(n1197), .Y(n1201) );
  INVX4 U90 ( .A(n1194), .Y(n1214) );
  INVX4 U91 ( .A(n1194), .Y(n1213) );
  INVX1 U92 ( .A(n1344), .Y(n1179) );
  INVX1 U93 ( .A(n1344), .Y(n1178) );
  INVX4 U94 ( .A(n1219), .Y(n1195) );
  INVX2 U95 ( .A(n1220), .Y(n1196) );
  INVX1 U96 ( .A(n1342), .Y(n1193) );
  INVX1 U97 ( .A(n1346), .Y(n1175) );
  INVX1 U98 ( .A(n1346), .Y(n1174) );
  INVX1 U99 ( .A(n1348), .Y(n1347) );
  INVX1 U100 ( .A(N14), .Y(n1348) );
  INVX1 U101 ( .A(N12), .Y(n1344) );
  INVX1 U102 ( .A(n1344), .Y(n1176) );
  INVX1 U103 ( .A(n1344), .Y(n1177) );
  INVX8 U104 ( .A(n1309), .Y(n1307) );
  INVX8 U105 ( .A(n1309), .Y(n1306) );
  INVX1 U106 ( .A(n103), .Y(n1275) );
  INVX1 U107 ( .A(n104), .Y(n1290) );
  INVX1 U108 ( .A(n105), .Y(n1305) );
  BUFX2 U109 ( .A(n107), .Y(n1247) );
  BUFX2 U110 ( .A(n121), .Y(n1262) );
  BUFX2 U111 ( .A(n135), .Y(n1277) );
  BUFX2 U112 ( .A(n149), .Y(n1292) );
  INVX1 U113 ( .A(n1346), .Y(n1345) );
  INVX1 U114 ( .A(N13), .Y(n1346) );
  INVX2 U115 ( .A(n1340), .Y(n1218) );
  INVX2 U116 ( .A(n1194), .Y(n1212) );
  INVX2 U117 ( .A(n1197), .Y(n1202) );
  INVX1 U118 ( .A(rst), .Y(n1339) );
  BUFX2 U119 ( .A(n157), .Y(n1300) );
  BUFX2 U120 ( .A(n159), .Y(n1302) );
  BUFX2 U121 ( .A(n161), .Y(n1304) );
  BUFX2 U122 ( .A(n151), .Y(n1294) );
  BUFX2 U123 ( .A(n153), .Y(n1296) );
  BUFX2 U124 ( .A(n155), .Y(n1298) );
  BUFX2 U125 ( .A(n123), .Y(n1264) );
  BUFX2 U126 ( .A(n127), .Y(n1268) );
  BUFX2 U127 ( .A(n143), .Y(n1285) );
  BUFX2 U128 ( .A(n147), .Y(n1289) );
  BUFX2 U129 ( .A(n109), .Y(n1249) );
  BUFX2 U130 ( .A(n111), .Y(n1251) );
  BUFX2 U131 ( .A(n113), .Y(n1253) );
  BUFX2 U132 ( .A(n115), .Y(n1255) );
  BUFX2 U133 ( .A(n117), .Y(n1257) );
  BUFX2 U134 ( .A(n119), .Y(n1259) );
  BUFX2 U135 ( .A(n125), .Y(n1266) );
  BUFX2 U136 ( .A(n129), .Y(n1270) );
  BUFX2 U137 ( .A(n131), .Y(n1272) );
  BUFX2 U138 ( .A(n133), .Y(n1274) );
  BUFX2 U139 ( .A(n137), .Y(n1279) );
  BUFX2 U140 ( .A(n139), .Y(n1281) );
  BUFX2 U141 ( .A(n141), .Y(n1283) );
  BUFX2 U142 ( .A(n145), .Y(n1287) );
  INVX1 U143 ( .A(n102), .Y(n1260) );
  INVX1 U144 ( .A(n1220), .Y(n1198) );
  INVX2 U145 ( .A(n1197), .Y(n1217) );
  INVX1 U146 ( .A(n1342), .Y(n1180) );
  INVX1 U147 ( .A(n1342), .Y(n1181) );
  INVX1 U148 ( .A(n1348), .Y(n1173) );
  INVX4 U149 ( .A(n7), .Y(n100) );
  INVX4 U150 ( .A(n6), .Y(n99) );
  INVX4 U151 ( .A(n5), .Y(n98) );
  INVX2 U152 ( .A(n4), .Y(n1) );
  BUFX2 U153 ( .A(write), .Y(n2) );
  INVX2 U154 ( .A(n4), .Y(n3) );
  INVX2 U155 ( .A(n4), .Y(n82) );
  OR2X2 U156 ( .A(write), .B(rst), .Y(n4) );
  AND2X2 U157 ( .A(n1307), .B(n156), .Y(n5) );
  AND2X2 U158 ( .A(n1307), .B(n158), .Y(n6) );
  AND2X2 U159 ( .A(n1307), .B(n160), .Y(n7) );
  AND2X2 U160 ( .A(\data_in<11> ), .B(n1307), .Y(n8) );
  AND2X2 U161 ( .A(\data_in<12> ), .B(n1307), .Y(n9) );
  AND2X2 U162 ( .A(\data_in<13> ), .B(n1307), .Y(n10) );
  AND2X2 U163 ( .A(\data_in<15> ), .B(n1307), .Y(n11) );
  AND2X2 U164 ( .A(n162), .B(n150), .Y(n12) );
  AND2X2 U165 ( .A(n162), .B(n152), .Y(n14) );
  AND2X2 U166 ( .A(n162), .B(n154), .Y(n16) );
  AND2X2 U167 ( .A(n1306), .B(n122), .Y(n18) );
  AND2X2 U168 ( .A(n1306), .B(n126), .Y(n20) );
  AND2X2 U169 ( .A(n163), .B(n142), .Y(n22) );
  AND2X2 U170 ( .A(n1307), .B(n146), .Y(n24) );
  AND2X2 U171 ( .A(n1306), .B(n106), .Y(n26) );
  AND2X2 U172 ( .A(n1306), .B(n108), .Y(n28) );
  AND2X2 U173 ( .A(n1306), .B(n110), .Y(n30) );
  AND2X2 U174 ( .A(n1306), .B(n112), .Y(n32) );
  AND2X2 U175 ( .A(n1306), .B(n114), .Y(n34) );
  AND2X2 U176 ( .A(n1306), .B(n116), .Y(n36) );
  AND2X2 U177 ( .A(n1306), .B(n118), .Y(n38) );
  AND2X2 U178 ( .A(n1306), .B(n102), .Y(n40) );
  AND2X2 U179 ( .A(n1306), .B(n120), .Y(n42) );
  AND2X2 U180 ( .A(n1306), .B(n124), .Y(n44) );
  AND2X2 U181 ( .A(n163), .B(n128), .Y(n46) );
  AND2X2 U182 ( .A(n1307), .B(n130), .Y(n48) );
  AND2X2 U183 ( .A(n1307), .B(n132), .Y(n50) );
  AND2X2 U184 ( .A(n163), .B(n103), .Y(n52) );
  AND2X2 U185 ( .A(n1307), .B(n134), .Y(n54) );
  AND2X2 U186 ( .A(n1307), .B(n136), .Y(n56) );
  AND2X2 U187 ( .A(n1307), .B(n138), .Y(n58) );
  AND2X2 U188 ( .A(n1306), .B(n140), .Y(n60) );
  AND2X2 U189 ( .A(n1307), .B(n144), .Y(n62) );
  AND2X2 U190 ( .A(n162), .B(n104), .Y(n64) );
  AND2X2 U191 ( .A(n162), .B(n148), .Y(n66) );
  AND2X2 U192 ( .A(n163), .B(n105), .Y(n68) );
  AND2X2 U193 ( .A(\data_in<14> ), .B(n163), .Y(n70) );
  AND2X2 U194 ( .A(n2), .B(n1339), .Y(n71) );
  AND2X2 U195 ( .A(\data_in<0> ), .B(n1308), .Y(n72) );
  AND2X2 U196 ( .A(\data_in<1> ), .B(n1308), .Y(n73) );
  AND2X2 U197 ( .A(\data_in<2> ), .B(n1308), .Y(n74) );
  AND2X2 U198 ( .A(\data_in<3> ), .B(n1308), .Y(n75) );
  AND2X2 U199 ( .A(\data_in<4> ), .B(n1308), .Y(n76) );
  AND2X2 U200 ( .A(\data_in<5> ), .B(n1308), .Y(n77) );
  AND2X2 U201 ( .A(\data_in<6> ), .B(n1308), .Y(n78) );
  AND2X2 U202 ( .A(\data_in<8> ), .B(n1308), .Y(n79) );
  AND2X2 U203 ( .A(\data_in<9> ), .B(n1308), .Y(n80) );
  AND2X2 U204 ( .A(\data_in<10> ), .B(n1308), .Y(n81) );
  INVX1 U205 ( .A(n1309), .Y(n162) );
  INVX1 U206 ( .A(n1341), .Y(n1340) );
  AND2X1 U207 ( .A(n1178), .B(n1342), .Y(n83) );
  INVX1 U208 ( .A(n1343), .Y(n1342) );
  AND2X1 U209 ( .A(n214), .B(n1347), .Y(n84) );
  INVX2 U210 ( .A(n1309), .Y(n1308) );
  BUFX2 U211 ( .A(n1381), .Y(n85) );
  INVX1 U212 ( .A(n85), .Y(n1773) );
  BUFX2 U213 ( .A(n1398), .Y(n86) );
  INVX1 U214 ( .A(n86), .Y(n1790) );
  BUFX2 U215 ( .A(n1415), .Y(n87) );
  INVX1 U216 ( .A(n87), .Y(n1807) );
  BUFX2 U217 ( .A(n1432), .Y(n88) );
  INVX1 U218 ( .A(n88), .Y(n1824) );
  BUFX2 U219 ( .A(n1449), .Y(n89) );
  INVX1 U220 ( .A(n89), .Y(n1841) );
  BUFX2 U221 ( .A(n1610), .Y(n90) );
  INVX1 U222 ( .A(n90), .Y(n1723) );
  BUFX2 U223 ( .A(n1740), .Y(n91) );
  INVX1 U224 ( .A(n91), .Y(n1858) );
  AND2X1 U225 ( .A(n1340), .B(n83), .Y(n92) );
  AND2X1 U226 ( .A(n1345), .B(n84), .Y(n93) );
  AND2X1 U227 ( .A(n1341), .B(n83), .Y(n94) );
  AND2X1 U228 ( .A(n1346), .B(n84), .Y(n95) );
  INVX1 U229 ( .A(n96), .Y(n97) );
  BUFX2 U230 ( .A(n101), .Y(n1243) );
  INVX1 U231 ( .A(n96), .Y(n101) );
  AND2X1 U232 ( .A(n93), .B(n1859), .Y(n102) );
  AND2X1 U233 ( .A(n1859), .B(n95), .Y(n103) );
  AND2X1 U234 ( .A(n1859), .B(n1723), .Y(n104) );
  AND2X1 U235 ( .A(n1859), .B(n1858), .Y(n105) );
  AND2X1 U236 ( .A(n92), .B(n93), .Y(n106) );
  INVX1 U237 ( .A(n106), .Y(n107) );
  AND2X1 U238 ( .A(n93), .B(n94), .Y(n108) );
  INVX1 U239 ( .A(n108), .Y(n109) );
  AND2X1 U240 ( .A(n93), .B(n1773), .Y(n110) );
  INVX1 U241 ( .A(n110), .Y(n111) );
  AND2X1 U242 ( .A(n93), .B(n1790), .Y(n112) );
  INVX1 U243 ( .A(n112), .Y(n113) );
  AND2X1 U244 ( .A(n93), .B(n1807), .Y(n114) );
  INVX1 U245 ( .A(n114), .Y(n115) );
  AND2X1 U246 ( .A(n93), .B(n1824), .Y(n116) );
  INVX1 U247 ( .A(n116), .Y(n117) );
  AND2X1 U248 ( .A(n93), .B(n1841), .Y(n118) );
  INVX1 U249 ( .A(n118), .Y(n119) );
  AND2X1 U250 ( .A(n92), .B(n95), .Y(n120) );
  INVX1 U251 ( .A(n120), .Y(n121) );
  AND2X1 U252 ( .A(n94), .B(n95), .Y(n122) );
  INVX1 U253 ( .A(n122), .Y(n123) );
  AND2X1 U254 ( .A(n1773), .B(n95), .Y(n124) );
  INVX1 U255 ( .A(n124), .Y(n125) );
  AND2X1 U256 ( .A(n1790), .B(n95), .Y(n126) );
  INVX1 U257 ( .A(n126), .Y(n127) );
  AND2X1 U258 ( .A(n1807), .B(n95), .Y(n128) );
  INVX1 U259 ( .A(n128), .Y(n129) );
  AND2X1 U260 ( .A(n1824), .B(n95), .Y(n130) );
  INVX1 U261 ( .A(n130), .Y(n131) );
  AND2X1 U262 ( .A(n1841), .B(n95), .Y(n132) );
  INVX1 U263 ( .A(n132), .Y(n133) );
  AND2X1 U264 ( .A(n92), .B(n1723), .Y(n134) );
  INVX1 U265 ( .A(n134), .Y(n135) );
  AND2X1 U266 ( .A(n94), .B(n1723), .Y(n136) );
  INVX1 U267 ( .A(n136), .Y(n137) );
  AND2X1 U268 ( .A(n1773), .B(n1723), .Y(n138) );
  INVX1 U269 ( .A(n138), .Y(n139) );
  AND2X1 U270 ( .A(n1790), .B(n1723), .Y(n140) );
  INVX1 U271 ( .A(n140), .Y(n141) );
  AND2X1 U272 ( .A(n1807), .B(n1723), .Y(n142) );
  INVX1 U273 ( .A(n142), .Y(n143) );
  AND2X1 U274 ( .A(n1824), .B(n1723), .Y(n144) );
  INVX1 U275 ( .A(n144), .Y(n145) );
  AND2X1 U276 ( .A(n1841), .B(n1723), .Y(n146) );
  INVX1 U277 ( .A(n146), .Y(n147) );
  AND2X1 U278 ( .A(n92), .B(n1858), .Y(n148) );
  INVX1 U279 ( .A(n148), .Y(n149) );
  AND2X1 U280 ( .A(n94), .B(n1858), .Y(n150) );
  INVX1 U281 ( .A(n150), .Y(n151) );
  AND2X1 U282 ( .A(n1773), .B(n1858), .Y(n152) );
  INVX1 U283 ( .A(n152), .Y(n153) );
  AND2X1 U284 ( .A(n1790), .B(n1858), .Y(n154) );
  INVX1 U285 ( .A(n154), .Y(n155) );
  AND2X1 U286 ( .A(n1807), .B(n1858), .Y(n156) );
  INVX1 U287 ( .A(n156), .Y(n157) );
  AND2X1 U288 ( .A(n1824), .B(n1858), .Y(n158) );
  INVX1 U289 ( .A(n158), .Y(n159) );
  AND2X1 U290 ( .A(n1841), .B(n1858), .Y(n160) );
  INVX1 U291 ( .A(n160), .Y(n161) );
  INVX1 U292 ( .A(n1309), .Y(n163) );
  MUX2X1 U293 ( .B(n165), .A(n166), .S(n1182), .Y(n164) );
  MUX2X1 U294 ( .B(n168), .A(n169), .S(n1182), .Y(n167) );
  MUX2X1 U295 ( .B(n171), .A(n172), .S(n1182), .Y(n170) );
  MUX2X1 U296 ( .B(n174), .A(n175), .S(n1182), .Y(n173) );
  MUX2X1 U297 ( .B(n177), .A(n178), .S(n1175), .Y(n176) );
  MUX2X1 U298 ( .B(n180), .A(n181), .S(n1182), .Y(n179) );
  MUX2X1 U299 ( .B(n183), .A(n184), .S(n1182), .Y(n182) );
  MUX2X1 U300 ( .B(n186), .A(n187), .S(n1182), .Y(n185) );
  MUX2X1 U301 ( .B(n189), .A(n190), .S(n1182), .Y(n188) );
  MUX2X1 U302 ( .B(n192), .A(n193), .S(n1175), .Y(n191) );
  MUX2X1 U303 ( .B(n195), .A(n196), .S(n1183), .Y(n194) );
  MUX2X1 U304 ( .B(n198), .A(n199), .S(n1183), .Y(n197) );
  MUX2X1 U305 ( .B(n201), .A(n202), .S(n1183), .Y(n200) );
  MUX2X1 U306 ( .B(n204), .A(n205), .S(n1183), .Y(n203) );
  MUX2X1 U307 ( .B(n207), .A(n208), .S(n1175), .Y(n206) );
  MUX2X1 U308 ( .B(n210), .A(n211), .S(n1183), .Y(n209) );
  MUX2X1 U309 ( .B(n213), .A(n215), .S(n1183), .Y(n212) );
  MUX2X1 U310 ( .B(n217), .A(n218), .S(n1183), .Y(n216) );
  MUX2X1 U311 ( .B(n220), .A(n221), .S(n1183), .Y(n219) );
  MUX2X1 U312 ( .B(n223), .A(n224), .S(n1175), .Y(n222) );
  MUX2X1 U313 ( .B(n226), .A(n227), .S(n1183), .Y(n225) );
  MUX2X1 U314 ( .B(n229), .A(n230), .S(n1183), .Y(n228) );
  MUX2X1 U315 ( .B(n232), .A(n233), .S(n1183), .Y(n231) );
  MUX2X1 U316 ( .B(n235), .A(n236), .S(n1183), .Y(n234) );
  MUX2X1 U317 ( .B(n238), .A(n239), .S(n1175), .Y(n237) );
  MUX2X1 U318 ( .B(n241), .A(n242), .S(n1184), .Y(n240) );
  MUX2X1 U319 ( .B(n244), .A(n245), .S(n1184), .Y(n243) );
  MUX2X1 U320 ( .B(n247), .A(n248), .S(n1184), .Y(n246) );
  MUX2X1 U321 ( .B(n250), .A(n251), .S(n1184), .Y(n249) );
  MUX2X1 U322 ( .B(n253), .A(n254), .S(n1175), .Y(n252) );
  MUX2X1 U323 ( .B(n256), .A(n257), .S(n1184), .Y(n255) );
  MUX2X1 U324 ( .B(n259), .A(n260), .S(n1184), .Y(n258) );
  MUX2X1 U325 ( .B(n262), .A(n263), .S(n1184), .Y(n261) );
  MUX2X1 U326 ( .B(n265), .A(n266), .S(n1184), .Y(n264) );
  MUX2X1 U327 ( .B(n268), .A(n269), .S(n1175), .Y(n267) );
  MUX2X1 U328 ( .B(n271), .A(n272), .S(n1184), .Y(n270) );
  MUX2X1 U329 ( .B(n274), .A(n275), .S(n1184), .Y(n273) );
  MUX2X1 U330 ( .B(n277), .A(n278), .S(n1184), .Y(n276) );
  MUX2X1 U331 ( .B(n280), .A(n281), .S(n1184), .Y(n279) );
  MUX2X1 U332 ( .B(n283), .A(n284), .S(n1175), .Y(n282) );
  MUX2X1 U333 ( .B(n286), .A(n287), .S(n1185), .Y(n285) );
  MUX2X1 U334 ( .B(n289), .A(n290), .S(n1185), .Y(n288) );
  MUX2X1 U335 ( .B(n292), .A(n293), .S(n1185), .Y(n291) );
  MUX2X1 U336 ( .B(n295), .A(n296), .S(n1185), .Y(n294) );
  MUX2X1 U337 ( .B(n298), .A(n299), .S(n1175), .Y(n297) );
  MUX2X1 U338 ( .B(n301), .A(n302), .S(n1185), .Y(n300) );
  MUX2X1 U339 ( .B(n304), .A(n305), .S(n1185), .Y(n303) );
  MUX2X1 U340 ( .B(n307), .A(n308), .S(n1185), .Y(n306) );
  MUX2X1 U341 ( .B(n310), .A(n311), .S(n1185), .Y(n309) );
  MUX2X1 U342 ( .B(n313), .A(n314), .S(n1175), .Y(n312) );
  MUX2X1 U343 ( .B(n316), .A(n317), .S(n1185), .Y(n315) );
  MUX2X1 U344 ( .B(n319), .A(n320), .S(n1185), .Y(n318) );
  MUX2X1 U345 ( .B(n322), .A(n323), .S(n1185), .Y(n321) );
  MUX2X1 U346 ( .B(n325), .A(n326), .S(n1185), .Y(n324) );
  MUX2X1 U347 ( .B(n328), .A(n329), .S(n1175), .Y(n327) );
  MUX2X1 U348 ( .B(n331), .A(n332), .S(n1186), .Y(n330) );
  MUX2X1 U349 ( .B(n334), .A(n335), .S(n1186), .Y(n333) );
  MUX2X1 U350 ( .B(n337), .A(n338), .S(n1186), .Y(n336) );
  MUX2X1 U351 ( .B(n340), .A(n341), .S(n1186), .Y(n339) );
  MUX2X1 U352 ( .B(n343), .A(n344), .S(n1175), .Y(n342) );
  MUX2X1 U353 ( .B(n346), .A(n347), .S(n1186), .Y(n345) );
  MUX2X1 U354 ( .B(n349), .A(n350), .S(n1186), .Y(n348) );
  MUX2X1 U355 ( .B(n352), .A(n353), .S(n1186), .Y(n351) );
  MUX2X1 U356 ( .B(n355), .A(n356), .S(n1186), .Y(n354) );
  MUX2X1 U357 ( .B(n358), .A(n359), .S(n1174), .Y(n357) );
  MUX2X1 U358 ( .B(n361), .A(n362), .S(n1186), .Y(n360) );
  MUX2X1 U359 ( .B(n364), .A(n365), .S(n1186), .Y(n363) );
  MUX2X1 U360 ( .B(n367), .A(n368), .S(n1186), .Y(n366) );
  MUX2X1 U361 ( .B(n370), .A(n371), .S(n1186), .Y(n369) );
  MUX2X1 U362 ( .B(n373), .A(n374), .S(n1174), .Y(n372) );
  MUX2X1 U363 ( .B(n376), .A(n377), .S(n1187), .Y(n375) );
  MUX2X1 U364 ( .B(n379), .A(n380), .S(n1187), .Y(n378) );
  MUX2X1 U365 ( .B(n382), .A(n383), .S(n1187), .Y(n381) );
  MUX2X1 U366 ( .B(n385), .A(n386), .S(n1187), .Y(n384) );
  MUX2X1 U367 ( .B(n388), .A(n389), .S(n1174), .Y(n387) );
  MUX2X1 U368 ( .B(n391), .A(n392), .S(n1187), .Y(n390) );
  MUX2X1 U369 ( .B(n394), .A(n395), .S(n1187), .Y(n393) );
  MUX2X1 U370 ( .B(n397), .A(n398), .S(n1187), .Y(n396) );
  MUX2X1 U371 ( .B(n400), .A(n401), .S(n1187), .Y(n399) );
  MUX2X1 U372 ( .B(n403), .A(n404), .S(n1174), .Y(n402) );
  MUX2X1 U373 ( .B(n406), .A(n407), .S(n1187), .Y(n405) );
  MUX2X1 U374 ( .B(n409), .A(n410), .S(n1187), .Y(n408) );
  MUX2X1 U375 ( .B(n412), .A(n413), .S(n1187), .Y(n411) );
  MUX2X1 U376 ( .B(n415), .A(n416), .S(n1187), .Y(n414) );
  MUX2X1 U377 ( .B(n418), .A(n419), .S(n1174), .Y(n417) );
  MUX2X1 U378 ( .B(n421), .A(n422), .S(n1188), .Y(n420) );
  MUX2X1 U379 ( .B(n424), .A(n425), .S(n1188), .Y(n423) );
  MUX2X1 U380 ( .B(n427), .A(n428), .S(n1188), .Y(n426) );
  MUX2X1 U381 ( .B(n430), .A(n431), .S(n1188), .Y(n429) );
  MUX2X1 U382 ( .B(n433), .A(n434), .S(n1174), .Y(n432) );
  MUX2X1 U383 ( .B(n436), .A(n437), .S(n1188), .Y(n435) );
  MUX2X1 U384 ( .B(n439), .A(n440), .S(n1188), .Y(n438) );
  MUX2X1 U385 ( .B(n442), .A(n443), .S(n1188), .Y(n441) );
  MUX2X1 U386 ( .B(n445), .A(n446), .S(n1188), .Y(n444) );
  MUX2X1 U387 ( .B(n448), .A(n449), .S(n1174), .Y(n447) );
  MUX2X1 U388 ( .B(n451), .A(n452), .S(n1188), .Y(n450) );
  MUX2X1 U389 ( .B(n454), .A(n455), .S(n1188), .Y(n453) );
  MUX2X1 U390 ( .B(n457), .A(n458), .S(n1188), .Y(n456) );
  MUX2X1 U391 ( .B(n460), .A(n461), .S(n1188), .Y(n459) );
  MUX2X1 U392 ( .B(n463), .A(n464), .S(n1174), .Y(n462) );
  MUX2X1 U393 ( .B(n466), .A(n467), .S(n1189), .Y(n465) );
  MUX2X1 U394 ( .B(n469), .A(n470), .S(n1189), .Y(n468) );
  MUX2X1 U395 ( .B(n472), .A(n473), .S(n1189), .Y(n471) );
  MUX2X1 U396 ( .B(n475), .A(n476), .S(n1189), .Y(n474) );
  MUX2X1 U397 ( .B(n478), .A(n479), .S(n1174), .Y(n477) );
  MUX2X1 U398 ( .B(n481), .A(n482), .S(n1189), .Y(n480) );
  MUX2X1 U399 ( .B(n484), .A(n485), .S(n1189), .Y(n483) );
  MUX2X1 U400 ( .B(n487), .A(n488), .S(n1189), .Y(n486) );
  MUX2X1 U401 ( .B(n490), .A(n491), .S(n1189), .Y(n489) );
  MUX2X1 U402 ( .B(n493), .A(n494), .S(n1174), .Y(n492) );
  MUX2X1 U403 ( .B(n496), .A(n497), .S(n1189), .Y(n495) );
  MUX2X1 U404 ( .B(n499), .A(n500), .S(n1189), .Y(n498) );
  MUX2X1 U405 ( .B(n502), .A(n503), .S(n1189), .Y(n501) );
  MUX2X1 U406 ( .B(n505), .A(n506), .S(n1189), .Y(n504) );
  MUX2X1 U407 ( .B(n508), .A(n509), .S(n1174), .Y(n507) );
  MUX2X1 U408 ( .B(n511), .A(n512), .S(n1190), .Y(n510) );
  MUX2X1 U409 ( .B(n514), .A(n515), .S(n1190), .Y(n513) );
  MUX2X1 U410 ( .B(n517), .A(n518), .S(n1190), .Y(n516) );
  MUX2X1 U411 ( .B(n520), .A(n521), .S(n1190), .Y(n519) );
  MUX2X1 U412 ( .B(n523), .A(n524), .S(n1174), .Y(n522) );
  MUX2X1 U413 ( .B(n526), .A(n527), .S(n1190), .Y(n525) );
  MUX2X1 U414 ( .B(n529), .A(n530), .S(n1190), .Y(n528) );
  MUX2X1 U415 ( .B(n532), .A(n533), .S(n1190), .Y(n531) );
  MUX2X1 U416 ( .B(n535), .A(n536), .S(n1190), .Y(n534) );
  MUX2X1 U417 ( .B(n538), .A(n539), .S(n1175), .Y(n537) );
  MUX2X1 U418 ( .B(n541), .A(n542), .S(n1190), .Y(n540) );
  MUX2X1 U419 ( .B(n544), .A(n545), .S(n1190), .Y(n543) );
  MUX2X1 U420 ( .B(n547), .A(n548), .S(n1190), .Y(n546) );
  MUX2X1 U421 ( .B(n550), .A(n551), .S(n1190), .Y(n549) );
  MUX2X1 U422 ( .B(n553), .A(n554), .S(n1175), .Y(n552) );
  MUX2X1 U423 ( .B(n556), .A(n557), .S(n1191), .Y(n555) );
  MUX2X1 U424 ( .B(n559), .A(n560), .S(n1191), .Y(n558) );
  MUX2X1 U425 ( .B(n562), .A(n563), .S(n1191), .Y(n561) );
  MUX2X1 U426 ( .B(n565), .A(n566), .S(n1191), .Y(n564) );
  MUX2X1 U427 ( .B(n568), .A(n569), .S(n1174), .Y(n567) );
  MUX2X1 U428 ( .B(n571), .A(n572), .S(n1191), .Y(n570) );
  MUX2X1 U429 ( .B(n574), .A(n575), .S(n1191), .Y(n573) );
  MUX2X1 U430 ( .B(n577), .A(n578), .S(n1191), .Y(n576) );
  MUX2X1 U431 ( .B(n580), .A(n581), .S(n1191), .Y(n579) );
  MUX2X1 U432 ( .B(n583), .A(n584), .S(n1174), .Y(n582) );
  MUX2X1 U433 ( .B(n586), .A(n587), .S(n1191), .Y(n585) );
  MUX2X1 U434 ( .B(n589), .A(n590), .S(n1191), .Y(n588) );
  MUX2X1 U435 ( .B(n592), .A(n593), .S(n1191), .Y(n591) );
  MUX2X1 U436 ( .B(n595), .A(n596), .S(n1191), .Y(n594) );
  MUX2X1 U437 ( .B(n598), .A(n599), .S(n1174), .Y(n597) );
  MUX2X1 U438 ( .B(n601), .A(n602), .S(n1192), .Y(n600) );
  MUX2X1 U439 ( .B(n604), .A(n605), .S(n1192), .Y(n603) );
  MUX2X1 U440 ( .B(n607), .A(n608), .S(n1192), .Y(n606) );
  MUX2X1 U441 ( .B(n610), .A(n611), .S(n1192), .Y(n609) );
  MUX2X1 U442 ( .B(n613), .A(n614), .S(n1174), .Y(n612) );
  MUX2X1 U443 ( .B(n616), .A(n617), .S(n1192), .Y(n615) );
  MUX2X1 U444 ( .B(n619), .A(n620), .S(n1192), .Y(n618) );
  MUX2X1 U445 ( .B(n622), .A(n623), .S(n1192), .Y(n621) );
  MUX2X1 U446 ( .B(n625), .A(n626), .S(n1192), .Y(n624) );
  MUX2X1 U447 ( .B(n628), .A(n629), .S(n1175), .Y(n627) );
  MUX2X1 U448 ( .B(n631), .A(n632), .S(n1192), .Y(n630) );
  MUX2X1 U449 ( .B(n634), .A(n635), .S(n1192), .Y(n633) );
  MUX2X1 U450 ( .B(n637), .A(n638), .S(n1192), .Y(n636) );
  MUX2X1 U451 ( .B(n640), .A(n641), .S(n1192), .Y(n639) );
  MUX2X1 U452 ( .B(n643), .A(n644), .S(n1175), .Y(n642) );
  MUX2X1 U453 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1201), .Y(n166) );
  MUX2X1 U454 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1217), .Y(n165) );
  MUX2X1 U455 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1205), .Y(n169) );
  MUX2X1 U456 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1217), .Y(n168) );
  MUX2X1 U457 ( .B(n167), .A(n164), .S(n1179), .Y(n178) );
  MUX2X1 U458 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1199), .Y(n172) );
  MUX2X1 U459 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1199), .Y(n171) );
  MUX2X1 U460 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1199), .Y(n175) );
  MUX2X1 U461 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1199), .Y(n174) );
  MUX2X1 U462 ( .B(n173), .A(n170), .S(n1179), .Y(n177) );
  MUX2X1 U463 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1199), .Y(n181) );
  MUX2X1 U464 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1199), .Y(n180) );
  MUX2X1 U465 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1199), .Y(n184) );
  MUX2X1 U466 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1199), .Y(n183) );
  MUX2X1 U467 ( .B(n182), .A(n179), .S(n1179), .Y(n193) );
  MUX2X1 U468 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1199), .Y(n187) );
  MUX2X1 U469 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1199), .Y(n186) );
  MUX2X1 U470 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1199), .Y(n190) );
  MUX2X1 U471 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1199), .Y(n189) );
  MUX2X1 U472 ( .B(n188), .A(n185), .S(n1179), .Y(n192) );
  MUX2X1 U473 ( .B(n191), .A(n176), .S(n1173), .Y(n645) );
  MUX2X1 U474 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1200), .Y(n196) );
  MUX2X1 U475 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1200), .Y(n195) );
  MUX2X1 U476 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1200), .Y(n199) );
  MUX2X1 U477 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1200), .Y(n198) );
  MUX2X1 U478 ( .B(n197), .A(n194), .S(n1179), .Y(n208) );
  MUX2X1 U479 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1200), .Y(n202) );
  MUX2X1 U480 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1200), .Y(n201) );
  MUX2X1 U481 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1200), .Y(n205) );
  MUX2X1 U482 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1200), .Y(n204) );
  MUX2X1 U483 ( .B(n203), .A(n200), .S(n1179), .Y(n207) );
  MUX2X1 U484 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1200), .Y(n211) );
  MUX2X1 U485 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1200), .Y(n210) );
  MUX2X1 U486 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1200), .Y(n215) );
  MUX2X1 U487 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1200), .Y(n213) );
  MUX2X1 U488 ( .B(n212), .A(n209), .S(n1179), .Y(n224) );
  MUX2X1 U489 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1201), .Y(n218) );
  MUX2X1 U490 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1214), .Y(n217) );
  MUX2X1 U491 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1201), .Y(n221) );
  MUX2X1 U492 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1201), .Y(n220) );
  MUX2X1 U493 ( .B(n219), .A(n216), .S(n1179), .Y(n223) );
  MUX2X1 U494 ( .B(n222), .A(n206), .S(n1173), .Y(n646) );
  MUX2X1 U495 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1213), .Y(n227) );
  MUX2X1 U496 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1214), .Y(n226) );
  MUX2X1 U497 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1201), .Y(n230) );
  MUX2X1 U498 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1201), .Y(n229) );
  MUX2X1 U499 ( .B(n228), .A(n225), .S(n1179), .Y(n239) );
  MUX2X1 U500 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1201), .Y(n233) );
  MUX2X1 U501 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1213), .Y(n232) );
  MUX2X1 U502 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1213), .Y(n236) );
  MUX2X1 U503 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1214), .Y(n235) );
  MUX2X1 U504 ( .B(n234), .A(n231), .S(n1179), .Y(n238) );
  MUX2X1 U505 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1201), .Y(n242) );
  MUX2X1 U506 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1201), .Y(n241) );
  MUX2X1 U507 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1201), .Y(n245) );
  MUX2X1 U508 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1201), .Y(n244) );
  MUX2X1 U509 ( .B(n243), .A(n240), .S(n1179), .Y(n254) );
  MUX2X1 U510 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1201), .Y(n248) );
  MUX2X1 U511 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1201), .Y(n247) );
  MUX2X1 U512 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1201), .Y(n251) );
  MUX2X1 U513 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1201), .Y(n250) );
  MUX2X1 U514 ( .B(n249), .A(n246), .S(n1179), .Y(n253) );
  MUX2X1 U515 ( .B(n252), .A(n237), .S(n1173), .Y(n647) );
  MUX2X1 U516 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1201), .Y(n257) );
  MUX2X1 U517 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1201), .Y(n256) );
  MUX2X1 U518 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1201), .Y(n260) );
  MUX2X1 U519 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1201), .Y(n259) );
  MUX2X1 U520 ( .B(n258), .A(n255), .S(n1178), .Y(n269) );
  MUX2X1 U521 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1202), .Y(n263) );
  MUX2X1 U522 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1202), .Y(n262) );
  MUX2X1 U523 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1202), .Y(n266) );
  MUX2X1 U524 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1202), .Y(n265) );
  MUX2X1 U525 ( .B(n264), .A(n261), .S(n1178), .Y(n268) );
  MUX2X1 U526 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1202), .Y(n272) );
  MUX2X1 U527 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1202), .Y(n271) );
  MUX2X1 U528 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1202), .Y(n275) );
  MUX2X1 U529 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1202), .Y(n274) );
  MUX2X1 U530 ( .B(n273), .A(n270), .S(n1178), .Y(n284) );
  MUX2X1 U531 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1202), .Y(n278) );
  MUX2X1 U532 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1202), .Y(n277) );
  MUX2X1 U533 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1202), .Y(n281) );
  MUX2X1 U534 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1202), .Y(n280) );
  MUX2X1 U535 ( .B(n279), .A(n276), .S(n1178), .Y(n283) );
  MUX2X1 U536 ( .B(n282), .A(n267), .S(n1173), .Y(n648) );
  MUX2X1 U537 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1203), .Y(n287) );
  MUX2X1 U538 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1203), .Y(n286) );
  MUX2X1 U539 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1203), .Y(n290) );
  MUX2X1 U540 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1203), .Y(n289) );
  MUX2X1 U541 ( .B(n288), .A(n285), .S(n1178), .Y(n299) );
  MUX2X1 U542 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1203), .Y(n293) );
  MUX2X1 U543 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1203), .Y(n292) );
  MUX2X1 U544 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1203), .Y(n296) );
  MUX2X1 U545 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1203), .Y(n295) );
  MUX2X1 U546 ( .B(n294), .A(n291), .S(n1178), .Y(n298) );
  MUX2X1 U547 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1203), .Y(n302) );
  MUX2X1 U548 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1203), .Y(n301) );
  MUX2X1 U549 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1203), .Y(n305) );
  MUX2X1 U550 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1203), .Y(n304) );
  MUX2X1 U551 ( .B(n303), .A(n300), .S(n1178), .Y(n314) );
  MUX2X1 U552 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1204), .Y(n308) );
  MUX2X1 U553 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1204), .Y(n307) );
  MUX2X1 U554 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1204), .Y(n311) );
  MUX2X1 U555 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1204), .Y(n310) );
  MUX2X1 U556 ( .B(n309), .A(n306), .S(n1178), .Y(n313) );
  MUX2X1 U557 ( .B(n312), .A(n297), .S(n1173), .Y(n649) );
  MUX2X1 U558 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1204), .Y(n317) );
  MUX2X1 U559 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1204), .Y(n316) );
  MUX2X1 U560 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1204), .Y(n320) );
  MUX2X1 U561 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1204), .Y(n319) );
  MUX2X1 U562 ( .B(n318), .A(n315), .S(n1178), .Y(n329) );
  MUX2X1 U563 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1204), .Y(n323) );
  MUX2X1 U564 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1204), .Y(n322) );
  MUX2X1 U565 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1204), .Y(n326) );
  MUX2X1 U566 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1204), .Y(n325) );
  MUX2X1 U567 ( .B(n324), .A(n321), .S(n1178), .Y(n328) );
  MUX2X1 U568 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1205), .Y(n332) );
  MUX2X1 U569 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1205), .Y(n331) );
  MUX2X1 U570 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1205), .Y(n335) );
  MUX2X1 U571 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1205), .Y(n334) );
  MUX2X1 U572 ( .B(n333), .A(n330), .S(n1178), .Y(n344) );
  MUX2X1 U573 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1205), .Y(n338) );
  MUX2X1 U574 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1205), .Y(n337) );
  MUX2X1 U575 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1205), .Y(n341) );
  MUX2X1 U576 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1205), .Y(n340) );
  MUX2X1 U577 ( .B(n339), .A(n336), .S(n1178), .Y(n343) );
  MUX2X1 U578 ( .B(n342), .A(n327), .S(n1173), .Y(n650) );
  MUX2X1 U579 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1205), .Y(n347) );
  MUX2X1 U580 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1205), .Y(n346) );
  MUX2X1 U581 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1205), .Y(n350) );
  MUX2X1 U582 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1205), .Y(n349) );
  MUX2X1 U583 ( .B(n348), .A(n345), .S(n1178), .Y(n359) );
  MUX2X1 U584 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1206), .Y(n353) );
  MUX2X1 U585 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1206), .Y(n352) );
  MUX2X1 U586 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1206), .Y(n356) );
  MUX2X1 U587 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1206), .Y(n355) );
  MUX2X1 U588 ( .B(n354), .A(n351), .S(n1178), .Y(n358) );
  MUX2X1 U589 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1206), .Y(n362) );
  MUX2X1 U590 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1206), .Y(n361) );
  MUX2X1 U591 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1206), .Y(n365) );
  MUX2X1 U592 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1206), .Y(n364) );
  MUX2X1 U593 ( .B(n363), .A(n360), .S(n1178), .Y(n374) );
  MUX2X1 U594 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1206), .Y(n368) );
  MUX2X1 U595 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1206), .Y(n367) );
  MUX2X1 U596 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1206), .Y(n371) );
  MUX2X1 U597 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1206), .Y(n370) );
  MUX2X1 U598 ( .B(n369), .A(n366), .S(n1178), .Y(n373) );
  MUX2X1 U599 ( .B(n372), .A(n357), .S(n1173), .Y(n1163) );
  MUX2X1 U600 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1207), .Y(n377) );
  MUX2X1 U601 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1207), .Y(n376) );
  MUX2X1 U602 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1207), .Y(n380) );
  MUX2X1 U603 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1207), .Y(n379) );
  MUX2X1 U604 ( .B(n378), .A(n375), .S(n1179), .Y(n389) );
  MUX2X1 U605 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1207), .Y(n383) );
  MUX2X1 U606 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1207), .Y(n382) );
  MUX2X1 U607 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1207), .Y(n386) );
  MUX2X1 U608 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1207), .Y(n385) );
  MUX2X1 U609 ( .B(n384), .A(n381), .S(n1179), .Y(n388) );
  MUX2X1 U610 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1207), .Y(n392) );
  MUX2X1 U611 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1207), .Y(n391) );
  MUX2X1 U612 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1207), .Y(n395) );
  MUX2X1 U613 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1207), .Y(n394) );
  MUX2X1 U614 ( .B(n393), .A(n390), .S(n1179), .Y(n404) );
  MUX2X1 U615 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1208), .Y(n398) );
  MUX2X1 U616 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1208), .Y(n397) );
  MUX2X1 U617 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1208), .Y(n401) );
  MUX2X1 U618 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1208), .Y(n400) );
  MUX2X1 U619 ( .B(n399), .A(n396), .S(n1179), .Y(n403) );
  MUX2X1 U620 ( .B(n402), .A(n387), .S(n1173), .Y(n1164) );
  MUX2X1 U621 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1208), .Y(n407) );
  MUX2X1 U622 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1208), .Y(n406) );
  MUX2X1 U623 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1208), .Y(n410) );
  MUX2X1 U624 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1208), .Y(n409) );
  MUX2X1 U625 ( .B(n408), .A(n405), .S(n1179), .Y(n419) );
  MUX2X1 U626 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1208), .Y(n413) );
  MUX2X1 U627 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1208), .Y(n412) );
  MUX2X1 U628 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1208), .Y(n416) );
  MUX2X1 U629 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1208), .Y(n415) );
  MUX2X1 U630 ( .B(n414), .A(n411), .S(n1178), .Y(n418) );
  MUX2X1 U631 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1209), .Y(n422) );
  MUX2X1 U632 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1209), .Y(n421) );
  MUX2X1 U633 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1209), .Y(n425) );
  MUX2X1 U634 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1209), .Y(n424) );
  MUX2X1 U635 ( .B(n423), .A(n420), .S(n1179), .Y(n434) );
  MUX2X1 U636 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1209), .Y(n428) );
  MUX2X1 U637 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1209), .Y(n427) );
  MUX2X1 U638 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1209), .Y(n431) );
  MUX2X1 U639 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1209), .Y(n430) );
  MUX2X1 U640 ( .B(n429), .A(n426), .S(n1178), .Y(n433) );
  MUX2X1 U641 ( .B(n432), .A(n417), .S(n1173), .Y(n1165) );
  MUX2X1 U642 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1209), .Y(n437) );
  MUX2X1 U643 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1209), .Y(n436) );
  MUX2X1 U644 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1209), .Y(n440) );
  MUX2X1 U645 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1209), .Y(n439) );
  MUX2X1 U646 ( .B(n438), .A(n435), .S(n1177), .Y(n449) );
  MUX2X1 U647 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1210), .Y(n443) );
  MUX2X1 U648 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1210), .Y(n442) );
  MUX2X1 U649 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1210), .Y(n446) );
  MUX2X1 U650 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1210), .Y(n445) );
  MUX2X1 U651 ( .B(n444), .A(n441), .S(n1177), .Y(n448) );
  MUX2X1 U652 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1210), .Y(n452) );
  MUX2X1 U653 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1210), .Y(n451) );
  MUX2X1 U654 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1210), .Y(n455) );
  MUX2X1 U655 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1210), .Y(n454) );
  MUX2X1 U656 ( .B(n453), .A(n450), .S(n1177), .Y(n464) );
  MUX2X1 U657 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1210), .Y(n458) );
  MUX2X1 U658 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1210), .Y(n457) );
  MUX2X1 U659 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1210), .Y(n461) );
  MUX2X1 U660 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1210), .Y(n460) );
  MUX2X1 U661 ( .B(n459), .A(n456), .S(n1177), .Y(n463) );
  MUX2X1 U662 ( .B(n462), .A(n447), .S(n1173), .Y(n1166) );
  MUX2X1 U663 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1211), .Y(n467) );
  MUX2X1 U664 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1211), .Y(n466) );
  MUX2X1 U665 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1211), .Y(n470) );
  MUX2X1 U666 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1211), .Y(n469) );
  MUX2X1 U667 ( .B(n468), .A(n465), .S(n1177), .Y(n479) );
  MUX2X1 U668 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1211), .Y(n473) );
  MUX2X1 U669 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1211), .Y(n472) );
  MUX2X1 U670 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1211), .Y(n476) );
  MUX2X1 U671 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1211), .Y(n475) );
  MUX2X1 U672 ( .B(n474), .A(n471), .S(n1177), .Y(n478) );
  MUX2X1 U673 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1211), .Y(n482) );
  MUX2X1 U674 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1211), .Y(n481) );
  MUX2X1 U675 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1211), .Y(n485) );
  MUX2X1 U676 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1211), .Y(n484) );
  MUX2X1 U677 ( .B(n483), .A(n480), .S(n1177), .Y(n494) );
  MUX2X1 U678 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1212), .Y(n488) );
  MUX2X1 U679 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1212), .Y(n487) );
  MUX2X1 U680 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1212), .Y(n491) );
  MUX2X1 U681 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1212), .Y(n490) );
  MUX2X1 U682 ( .B(n489), .A(n486), .S(n1177), .Y(n493) );
  MUX2X1 U683 ( .B(n492), .A(n477), .S(n1173), .Y(n1167) );
  MUX2X1 U684 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1212), .Y(n497) );
  MUX2X1 U685 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1212), .Y(n496) );
  MUX2X1 U686 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1212), .Y(n500) );
  MUX2X1 U687 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1212), .Y(n499) );
  MUX2X1 U688 ( .B(n498), .A(n495), .S(n1177), .Y(n509) );
  MUX2X1 U689 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1212), .Y(n503) );
  MUX2X1 U690 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1212), .Y(n502) );
  MUX2X1 U691 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1212), .Y(n506) );
  MUX2X1 U692 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1212), .Y(n505) );
  MUX2X1 U693 ( .B(n504), .A(n501), .S(n1177), .Y(n508) );
  MUX2X1 U694 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1213), .Y(n512) );
  MUX2X1 U695 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1213), .Y(n511) );
  MUX2X1 U696 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1213), .Y(n515) );
  MUX2X1 U697 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1213), .Y(n514) );
  MUX2X1 U698 ( .B(n513), .A(n510), .S(n1177), .Y(n524) );
  MUX2X1 U699 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1213), .Y(n518) );
  MUX2X1 U700 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1213), .Y(n517) );
  MUX2X1 U701 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1213), .Y(n521) );
  MUX2X1 U702 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1213), .Y(n520) );
  MUX2X1 U703 ( .B(n519), .A(n516), .S(n1177), .Y(n523) );
  MUX2X1 U704 ( .B(n522), .A(n507), .S(n1173), .Y(n1168) );
  MUX2X1 U705 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1213), .Y(n527) );
  MUX2X1 U706 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1213), .Y(n526) );
  MUX2X1 U707 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1213), .Y(n530) );
  MUX2X1 U708 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1213), .Y(n529) );
  MUX2X1 U709 ( .B(n528), .A(n525), .S(n1176), .Y(n539) );
  MUX2X1 U710 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1214), .Y(n533) );
  MUX2X1 U711 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1214), .Y(n532) );
  MUX2X1 U712 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1214), .Y(n536) );
  MUX2X1 U713 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1214), .Y(n535) );
  MUX2X1 U714 ( .B(n534), .A(n531), .S(n1176), .Y(n538) );
  MUX2X1 U715 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1214), .Y(n542) );
  MUX2X1 U716 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1214), .Y(n541) );
  MUX2X1 U717 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1214), .Y(n545) );
  MUX2X1 U718 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1214), .Y(n544) );
  MUX2X1 U719 ( .B(n543), .A(n540), .S(n1176), .Y(n554) );
  MUX2X1 U720 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1214), .Y(n548) );
  MUX2X1 U721 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1214), .Y(n547) );
  MUX2X1 U722 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1214), .Y(n551) );
  MUX2X1 U723 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1214), .Y(n550) );
  MUX2X1 U724 ( .B(n549), .A(n546), .S(n1176), .Y(n553) );
  MUX2X1 U725 ( .B(n552), .A(n537), .S(n1173), .Y(n1169) );
  MUX2X1 U726 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1215), .Y(n557) );
  MUX2X1 U727 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1215), .Y(n556) );
  MUX2X1 U728 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1215), .Y(n560) );
  MUX2X1 U729 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1215), .Y(n559) );
  MUX2X1 U730 ( .B(n558), .A(n555), .S(n1176), .Y(n569) );
  MUX2X1 U731 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1215), .Y(n563) );
  MUX2X1 U732 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1215), .Y(n562) );
  MUX2X1 U733 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1215), .Y(n566) );
  MUX2X1 U734 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1215), .Y(n565) );
  MUX2X1 U735 ( .B(n564), .A(n561), .S(n1176), .Y(n568) );
  MUX2X1 U736 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1215), .Y(n572) );
  MUX2X1 U737 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1215), .Y(n571) );
  MUX2X1 U738 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1215), .Y(n575) );
  MUX2X1 U739 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1215), .Y(n574) );
  MUX2X1 U740 ( .B(n573), .A(n570), .S(n1176), .Y(n584) );
  MUX2X1 U741 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1216), .Y(n578) );
  MUX2X1 U742 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1216), .Y(n577) );
  MUX2X1 U743 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1216), .Y(n581) );
  MUX2X1 U744 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1216), .Y(n580) );
  MUX2X1 U745 ( .B(n579), .A(n576), .S(n1176), .Y(n583) );
  MUX2X1 U746 ( .B(n582), .A(n567), .S(n1173), .Y(n1170) );
  MUX2X1 U747 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1216), .Y(n587) );
  MUX2X1 U748 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1216), .Y(n586) );
  MUX2X1 U749 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1216), .Y(n590) );
  MUX2X1 U750 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1216), .Y(n589) );
  MUX2X1 U751 ( .B(n588), .A(n585), .S(n1176), .Y(n599) );
  MUX2X1 U752 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1216), .Y(n593) );
  MUX2X1 U753 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1216), .Y(n592) );
  MUX2X1 U754 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1216), .Y(n596) );
  MUX2X1 U755 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1216), .Y(n595) );
  MUX2X1 U756 ( .B(n594), .A(n591), .S(n1176), .Y(n598) );
  MUX2X1 U757 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1217), .Y(n602) );
  MUX2X1 U758 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1217), .Y(n601) );
  MUX2X1 U759 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1217), .Y(n605) );
  MUX2X1 U760 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1217), .Y(n604) );
  MUX2X1 U761 ( .B(n603), .A(n600), .S(n1176), .Y(n614) );
  MUX2X1 U762 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1217), .Y(n608) );
  MUX2X1 U763 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1217), .Y(n607) );
  MUX2X1 U764 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1217), .Y(n611) );
  MUX2X1 U765 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1217), .Y(n610) );
  MUX2X1 U766 ( .B(n609), .A(n606), .S(n1176), .Y(n613) );
  MUX2X1 U767 ( .B(n612), .A(n597), .S(n1173), .Y(n1171) );
  MUX2X1 U768 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1217), .Y(n617) );
  MUX2X1 U769 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1217), .Y(n616) );
  MUX2X1 U770 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1217), .Y(n620) );
  MUX2X1 U771 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1217), .Y(n619) );
  MUX2X1 U772 ( .B(n618), .A(n615), .S(n1176), .Y(n629) );
  MUX2X1 U773 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1204), .Y(n623) );
  MUX2X1 U774 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1212), .Y(n622) );
  MUX2X1 U775 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1204), .Y(n626) );
  MUX2X1 U776 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1201), .Y(n625) );
  MUX2X1 U777 ( .B(n624), .A(n621), .S(n1177), .Y(n628) );
  MUX2X1 U778 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1202), .Y(n632) );
  MUX2X1 U779 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1201), .Y(n631) );
  MUX2X1 U780 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1219), .Y(n635) );
  MUX2X1 U781 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1219), .Y(n634) );
  MUX2X1 U782 ( .B(n633), .A(n630), .S(n1176), .Y(n644) );
  MUX2X1 U783 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1203), .Y(n638) );
  MUX2X1 U784 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1201), .Y(n637) );
  MUX2X1 U785 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1219), .Y(n641) );
  MUX2X1 U786 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1219), .Y(n640) );
  MUX2X1 U787 ( .B(n639), .A(n636), .S(n1177), .Y(n643) );
  MUX2X1 U788 ( .B(n642), .A(n627), .S(n1173), .Y(n1172) );
  INVX8 U789 ( .A(n1219), .Y(n1194) );
  INVX8 U790 ( .A(n1220), .Y(n1197) );
  INVX8 U791 ( .A(n1198), .Y(n1199) );
  INVX8 U792 ( .A(n1198), .Y(n1200) );
  INVX8 U793 ( .A(n1196), .Y(n1203) );
  INVX8 U794 ( .A(n1196), .Y(n1204) );
  INVX8 U795 ( .A(n1196), .Y(n1205) );
  INVX8 U796 ( .A(n1195), .Y(n1206) );
  INVX8 U797 ( .A(n1195), .Y(n1207) );
  INVX8 U798 ( .A(n1195), .Y(n1208) );
  INVX8 U799 ( .A(n1195), .Y(n1209) );
  INVX8 U800 ( .A(n1195), .Y(n1210) );
  INVX8 U801 ( .A(n1195), .Y(n1211) );
  INVX8 U802 ( .A(n1196), .Y(n1215) );
  INVX8 U803 ( .A(n1196), .Y(n1216) );
  INVX8 U804 ( .A(n1218), .Y(n1219) );
  INVX8 U805 ( .A(n1218), .Y(n1220) );
  INVX1 U806 ( .A(n1245), .Y(n1221) );
  INVX1 U807 ( .A(n1245), .Y(n1222) );
  INVX1 U808 ( .A(n1245), .Y(n1223) );
  INVX1 U809 ( .A(n70), .Y(n1224) );
  INVX1 U810 ( .A(n70), .Y(n1225) );
  INVX1 U811 ( .A(n70), .Y(n1226) );
  INVX1 U812 ( .A(n70), .Y(n1227) );
  INVX1 U813 ( .A(n70), .Y(n1228) );
  INVX1 U814 ( .A(n70), .Y(n1229) );
  INVX1 U815 ( .A(n1336), .Y(n1230) );
  INVX1 U816 ( .A(n1336), .Y(n1231) );
  INVX1 U817 ( .A(n1336), .Y(n1232) );
  INVX1 U818 ( .A(n1336), .Y(n1233) );
  INVX1 U819 ( .A(n1336), .Y(n1234) );
  INVX1 U820 ( .A(n1336), .Y(n1235) );
  INVX1 U821 ( .A(n1245), .Y(n1236) );
  INVX1 U822 ( .A(n1336), .Y(n1237) );
  INVX1 U823 ( .A(n1228), .Y(n1336) );
  INVX1 U824 ( .A(n96), .Y(n1238) );
  INVX1 U825 ( .A(n96), .Y(n1239) );
  INVX1 U826 ( .A(n96), .Y(n1240) );
  INVX1 U827 ( .A(n96), .Y(n1241) );
  BUFX2 U828 ( .A(n101), .Y(n1244) );
  INVX1 U829 ( .A(n1229), .Y(n1245) );
  INVX1 U830 ( .A(N11), .Y(n1343) );
  INVX1 U831 ( .A(N10), .Y(n1341) );
  INVX8 U832 ( .A(n72), .Y(n1310) );
  INVX8 U833 ( .A(n72), .Y(n1311) );
  INVX8 U834 ( .A(n73), .Y(n1312) );
  INVX8 U835 ( .A(n73), .Y(n1313) );
  INVX8 U836 ( .A(n74), .Y(n1314) );
  INVX8 U837 ( .A(n74), .Y(n1315) );
  INVX8 U838 ( .A(n75), .Y(n1316) );
  INVX8 U839 ( .A(n75), .Y(n1317) );
  INVX8 U840 ( .A(n76), .Y(n1318) );
  INVX8 U841 ( .A(n76), .Y(n1319) );
  INVX8 U842 ( .A(n77), .Y(n1320) );
  INVX8 U843 ( .A(n77), .Y(n1321) );
  INVX8 U844 ( .A(n78), .Y(n1322) );
  INVX8 U845 ( .A(n78), .Y(n1323) );
  INVX8 U846 ( .A(n79), .Y(n1324) );
  INVX8 U847 ( .A(n79), .Y(n1325) );
  INVX8 U848 ( .A(n80), .Y(n1326) );
  INVX8 U849 ( .A(n80), .Y(n1327) );
  INVX8 U850 ( .A(n81), .Y(n1328) );
  INVX8 U851 ( .A(n81), .Y(n1329) );
  INVX8 U852 ( .A(n8), .Y(n1330) );
  INVX8 U853 ( .A(n8), .Y(n1331) );
  INVX8 U854 ( .A(n9), .Y(n1332) );
  INVX8 U855 ( .A(n9), .Y(n1333) );
  INVX8 U856 ( .A(n10), .Y(n1334) );
  INVX8 U857 ( .A(n10), .Y(n1335) );
  INVX8 U858 ( .A(n11), .Y(n1337) );
  INVX8 U859 ( .A(n11), .Y(n1338) );
  AND2X2 U860 ( .A(n82), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U861 ( .A(n1), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U862 ( .A(N30), .B(n3), .Y(\data_out<2> ) );
  AND2X2 U863 ( .A(n82), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U864 ( .A(n82), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U865 ( .A(n82), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U866 ( .A(n1), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U867 ( .A(n1), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U868 ( .A(N24), .B(n3), .Y(\data_out<8> ) );
  AND2X2 U869 ( .A(n82), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U870 ( .A(N22), .B(n3), .Y(\data_out<10> ) );
  AND2X2 U871 ( .A(n82), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U872 ( .A(n1), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U873 ( .A(n1), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U874 ( .A(N18), .B(n3), .Y(\data_out<14> ) );
  AND2X2 U875 ( .A(n1), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U876 ( .A(\mem<31><0> ), .B(n27), .Y(n1349) );
  OAI21X1 U877 ( .A(n1247), .B(n1310), .C(n1349), .Y(n651) );
  NAND2X1 U878 ( .A(\mem<31><1> ), .B(n27), .Y(n1350) );
  OAI21X1 U879 ( .A(n1313), .B(n1246), .C(n1350), .Y(n652) );
  NAND2X1 U880 ( .A(\mem<31><2> ), .B(n27), .Y(n1351) );
  OAI21X1 U881 ( .A(n1315), .B(n1246), .C(n1351), .Y(n653) );
  NAND2X1 U882 ( .A(\mem<31><3> ), .B(n27), .Y(n1352) );
  OAI21X1 U883 ( .A(n1317), .B(n1246), .C(n1352), .Y(n654) );
  NAND2X1 U884 ( .A(\mem<31><4> ), .B(n27), .Y(n1353) );
  OAI21X1 U885 ( .A(n1319), .B(n1246), .C(n1353), .Y(n655) );
  NAND2X1 U886 ( .A(\mem<31><5> ), .B(n27), .Y(n1354) );
  OAI21X1 U887 ( .A(n1321), .B(n1246), .C(n1354), .Y(n656) );
  NAND2X1 U888 ( .A(\mem<31><6> ), .B(n27), .Y(n1355) );
  OAI21X1 U889 ( .A(n1323), .B(n1246), .C(n1355), .Y(n657) );
  NAND2X1 U890 ( .A(\mem<31><7> ), .B(n27), .Y(n1356) );
  OAI21X1 U891 ( .A(n1243), .B(n1246), .C(n1356), .Y(n658) );
  NAND2X1 U892 ( .A(\mem<31><8> ), .B(n27), .Y(n1357) );
  OAI21X1 U893 ( .A(n1325), .B(n1246), .C(n1357), .Y(n659) );
  NAND2X1 U894 ( .A(\mem<31><9> ), .B(n27), .Y(n1358) );
  OAI21X1 U895 ( .A(n1327), .B(n1247), .C(n1358), .Y(n660) );
  NAND2X1 U896 ( .A(\mem<31><10> ), .B(n27), .Y(n1359) );
  OAI21X1 U897 ( .A(n1329), .B(n1247), .C(n1359), .Y(n661) );
  NAND2X1 U898 ( .A(\mem<31><11> ), .B(n27), .Y(n1360) );
  OAI21X1 U899 ( .A(n1331), .B(n1247), .C(n1360), .Y(n662) );
  NAND2X1 U900 ( .A(\mem<31><12> ), .B(n27), .Y(n1361) );
  OAI21X1 U901 ( .A(n1333), .B(n1247), .C(n1361), .Y(n663) );
  NAND2X1 U902 ( .A(\mem<31><13> ), .B(n27), .Y(n1362) );
  OAI21X1 U903 ( .A(n1335), .B(n1247), .C(n1362), .Y(n664) );
  NAND2X1 U904 ( .A(\mem<31><14> ), .B(n27), .Y(n1363) );
  OAI21X1 U905 ( .A(n1221), .B(n1247), .C(n1363), .Y(n665) );
  NAND2X1 U906 ( .A(\mem<31><15> ), .B(n27), .Y(n1364) );
  OAI21X1 U907 ( .A(n1338), .B(n1247), .C(n1364), .Y(n666) );
  NAND2X1 U908 ( .A(\mem<30><0> ), .B(n29), .Y(n1365) );
  OAI21X1 U909 ( .A(n1248), .B(n1310), .C(n1365), .Y(n667) );
  NAND2X1 U910 ( .A(\mem<30><1> ), .B(n29), .Y(n1366) );
  OAI21X1 U911 ( .A(n1248), .B(n1313), .C(n1366), .Y(n668) );
  NAND2X1 U912 ( .A(\mem<30><2> ), .B(n29), .Y(n1367) );
  OAI21X1 U913 ( .A(n1248), .B(n1315), .C(n1367), .Y(n669) );
  NAND2X1 U914 ( .A(\mem<30><3> ), .B(n29), .Y(n1368) );
  OAI21X1 U915 ( .A(n1248), .B(n1317), .C(n1368), .Y(n670) );
  NAND2X1 U916 ( .A(\mem<30><4> ), .B(n29), .Y(n1369) );
  OAI21X1 U917 ( .A(n1248), .B(n1319), .C(n1369), .Y(n671) );
  NAND2X1 U918 ( .A(\mem<30><5> ), .B(n29), .Y(n1370) );
  OAI21X1 U919 ( .A(n1248), .B(n1321), .C(n1370), .Y(n672) );
  NAND2X1 U920 ( .A(\mem<30><6> ), .B(n29), .Y(n1371) );
  OAI21X1 U921 ( .A(n1248), .B(n1323), .C(n1371), .Y(n673) );
  NAND2X1 U922 ( .A(\mem<30><7> ), .B(n29), .Y(n1372) );
  OAI21X1 U923 ( .A(n1248), .B(n1239), .C(n1372), .Y(n674) );
  NAND2X1 U924 ( .A(\mem<30><8> ), .B(n29), .Y(n1373) );
  OAI21X1 U925 ( .A(n1249), .B(n1325), .C(n1373), .Y(n675) );
  NAND2X1 U926 ( .A(\mem<30><9> ), .B(n29), .Y(n1374) );
  OAI21X1 U927 ( .A(n1249), .B(n1327), .C(n1374), .Y(n676) );
  NAND2X1 U928 ( .A(\mem<30><10> ), .B(n29), .Y(n1375) );
  OAI21X1 U929 ( .A(n1249), .B(n1329), .C(n1375), .Y(n677) );
  NAND2X1 U930 ( .A(\mem<30><11> ), .B(n29), .Y(n1376) );
  OAI21X1 U931 ( .A(n1249), .B(n1331), .C(n1376), .Y(n678) );
  NAND2X1 U932 ( .A(\mem<30><12> ), .B(n29), .Y(n1377) );
  OAI21X1 U933 ( .A(n1249), .B(n1333), .C(n1377), .Y(n679) );
  NAND2X1 U934 ( .A(\mem<30><13> ), .B(n29), .Y(n1378) );
  OAI21X1 U935 ( .A(n1249), .B(n1335), .C(n1378), .Y(n680) );
  NAND2X1 U936 ( .A(\mem<30><14> ), .B(n29), .Y(n1379) );
  OAI21X1 U937 ( .A(n1249), .B(n1230), .C(n1379), .Y(n681) );
  NAND2X1 U938 ( .A(\mem<30><15> ), .B(n29), .Y(n1380) );
  OAI21X1 U939 ( .A(n1249), .B(n1338), .C(n1380), .Y(n682) );
  NAND3X1 U940 ( .A(n1340), .B(n1179), .C(n1343), .Y(n1381) );
  NAND2X1 U941 ( .A(\mem<29><0> ), .B(n31), .Y(n1382) );
  OAI21X1 U942 ( .A(n1250), .B(n1310), .C(n1382), .Y(n683) );
  NAND2X1 U943 ( .A(\mem<29><1> ), .B(n31), .Y(n1383) );
  OAI21X1 U944 ( .A(n1250), .B(n1313), .C(n1383), .Y(n684) );
  NAND2X1 U945 ( .A(\mem<29><2> ), .B(n31), .Y(n1384) );
  OAI21X1 U946 ( .A(n1250), .B(n1315), .C(n1384), .Y(n685) );
  NAND2X1 U947 ( .A(\mem<29><3> ), .B(n31), .Y(n1385) );
  OAI21X1 U948 ( .A(n1250), .B(n1317), .C(n1385), .Y(n686) );
  NAND2X1 U949 ( .A(\mem<29><4> ), .B(n31), .Y(n1386) );
  OAI21X1 U950 ( .A(n1250), .B(n1319), .C(n1386), .Y(n687) );
  NAND2X1 U951 ( .A(\mem<29><5> ), .B(n31), .Y(n1387) );
  OAI21X1 U952 ( .A(n1250), .B(n1321), .C(n1387), .Y(n688) );
  NAND2X1 U953 ( .A(\mem<29><6> ), .B(n31), .Y(n1388) );
  OAI21X1 U954 ( .A(n1250), .B(n1323), .C(n1388), .Y(n689) );
  NAND2X1 U955 ( .A(\mem<29><7> ), .B(n31), .Y(n1389) );
  OAI21X1 U956 ( .A(n1250), .B(n1240), .C(n1389), .Y(n690) );
  NAND2X1 U957 ( .A(\mem<29><8> ), .B(n31), .Y(n1390) );
  OAI21X1 U958 ( .A(n1251), .B(n1325), .C(n1390), .Y(n691) );
  NAND2X1 U959 ( .A(\mem<29><9> ), .B(n31), .Y(n1391) );
  OAI21X1 U960 ( .A(n1251), .B(n1327), .C(n1391), .Y(n692) );
  NAND2X1 U961 ( .A(\mem<29><10> ), .B(n31), .Y(n1392) );
  OAI21X1 U962 ( .A(n1251), .B(n1329), .C(n1392), .Y(n693) );
  NAND2X1 U963 ( .A(\mem<29><11> ), .B(n31), .Y(n1393) );
  OAI21X1 U964 ( .A(n1251), .B(n1331), .C(n1393), .Y(n694) );
  NAND2X1 U965 ( .A(\mem<29><12> ), .B(n31), .Y(n1394) );
  OAI21X1 U966 ( .A(n1251), .B(n1333), .C(n1394), .Y(n695) );
  NAND2X1 U967 ( .A(\mem<29><13> ), .B(n31), .Y(n1395) );
  OAI21X1 U968 ( .A(n1251), .B(n1335), .C(n1395), .Y(n696) );
  NAND2X1 U969 ( .A(\mem<29><14> ), .B(n31), .Y(n1396) );
  OAI21X1 U970 ( .A(n1251), .B(n1227), .C(n1396), .Y(n697) );
  NAND2X1 U971 ( .A(\mem<29><15> ), .B(n31), .Y(n1397) );
  OAI21X1 U972 ( .A(n1251), .B(n1338), .C(n1397), .Y(n698) );
  NAND3X1 U973 ( .A(n1178), .B(n1343), .C(n1341), .Y(n1398) );
  NAND2X1 U974 ( .A(\mem<28><0> ), .B(n33), .Y(n1399) );
  OAI21X1 U975 ( .A(n1252), .B(n1310), .C(n1399), .Y(n699) );
  NAND2X1 U976 ( .A(\mem<28><1> ), .B(n33), .Y(n1400) );
  OAI21X1 U977 ( .A(n1252), .B(n1313), .C(n1400), .Y(n700) );
  NAND2X1 U978 ( .A(\mem<28><2> ), .B(n33), .Y(n1401) );
  OAI21X1 U979 ( .A(n1252), .B(n1315), .C(n1401), .Y(n701) );
  NAND2X1 U980 ( .A(\mem<28><3> ), .B(n33), .Y(n1402) );
  OAI21X1 U981 ( .A(n1252), .B(n1317), .C(n1402), .Y(n702) );
  NAND2X1 U982 ( .A(\mem<28><4> ), .B(n33), .Y(n1403) );
  OAI21X1 U983 ( .A(n1252), .B(n1319), .C(n1403), .Y(n703) );
  NAND2X1 U984 ( .A(\mem<28><5> ), .B(n33), .Y(n1404) );
  OAI21X1 U985 ( .A(n1252), .B(n1321), .C(n1404), .Y(n704) );
  NAND2X1 U986 ( .A(\mem<28><6> ), .B(n33), .Y(n1405) );
  OAI21X1 U987 ( .A(n1252), .B(n1323), .C(n1405), .Y(n705) );
  NAND2X1 U988 ( .A(\mem<28><7> ), .B(n33), .Y(n1406) );
  OAI21X1 U989 ( .A(n1252), .B(n1241), .C(n1406), .Y(n706) );
  NAND2X1 U990 ( .A(\mem<28><8> ), .B(n33), .Y(n1407) );
  OAI21X1 U991 ( .A(n1253), .B(n1325), .C(n1407), .Y(n707) );
  NAND2X1 U992 ( .A(\mem<28><9> ), .B(n33), .Y(n1408) );
  OAI21X1 U993 ( .A(n1253), .B(n1327), .C(n1408), .Y(n708) );
  NAND2X1 U994 ( .A(\mem<28><10> ), .B(n33), .Y(n1409) );
  OAI21X1 U995 ( .A(n1253), .B(n1329), .C(n1409), .Y(n709) );
  NAND2X1 U996 ( .A(\mem<28><11> ), .B(n33), .Y(n1410) );
  OAI21X1 U997 ( .A(n1253), .B(n1331), .C(n1410), .Y(n710) );
  NAND2X1 U998 ( .A(\mem<28><12> ), .B(n33), .Y(n1411) );
  OAI21X1 U999 ( .A(n1253), .B(n1333), .C(n1411), .Y(n711) );
  NAND2X1 U1000 ( .A(\mem<28><13> ), .B(n33), .Y(n1412) );
  OAI21X1 U1001 ( .A(n1253), .B(n1335), .C(n1412), .Y(n712) );
  NAND2X1 U1002 ( .A(\mem<28><14> ), .B(n33), .Y(n1413) );
  OAI21X1 U1003 ( .A(n1253), .B(n1228), .C(n1413), .Y(n713) );
  NAND2X1 U1004 ( .A(\mem<28><15> ), .B(n33), .Y(n1414) );
  OAI21X1 U1005 ( .A(n1253), .B(n1338), .C(n1414), .Y(n714) );
  NAND3X1 U1006 ( .A(n1340), .B(n1342), .C(n1344), .Y(n1415) );
  NAND2X1 U1007 ( .A(\mem<27><0> ), .B(n35), .Y(n1416) );
  OAI21X1 U1008 ( .A(n1254), .B(n1310), .C(n1416), .Y(n715) );
  NAND2X1 U1009 ( .A(\mem<27><1> ), .B(n35), .Y(n1417) );
  OAI21X1 U1010 ( .A(n1254), .B(n1313), .C(n1417), .Y(n716) );
  NAND2X1 U1011 ( .A(\mem<27><2> ), .B(n35), .Y(n1418) );
  OAI21X1 U1012 ( .A(n1254), .B(n1315), .C(n1418), .Y(n717) );
  NAND2X1 U1013 ( .A(\mem<27><3> ), .B(n35), .Y(n1419) );
  OAI21X1 U1014 ( .A(n1254), .B(n1317), .C(n1419), .Y(n718) );
  NAND2X1 U1015 ( .A(\mem<27><4> ), .B(n35), .Y(n1420) );
  OAI21X1 U1016 ( .A(n1254), .B(n1319), .C(n1420), .Y(n719) );
  NAND2X1 U1017 ( .A(\mem<27><5> ), .B(n35), .Y(n1421) );
  OAI21X1 U1018 ( .A(n1254), .B(n1321), .C(n1421), .Y(n720) );
  NAND2X1 U1019 ( .A(\mem<27><6> ), .B(n35), .Y(n1422) );
  OAI21X1 U1020 ( .A(n1254), .B(n1323), .C(n1422), .Y(n721) );
  NAND2X1 U1021 ( .A(\mem<27><7> ), .B(n35), .Y(n1423) );
  OAI21X1 U1022 ( .A(n1254), .B(n1241), .C(n1423), .Y(n722) );
  NAND2X1 U1023 ( .A(\mem<27><8> ), .B(n35), .Y(n1424) );
  OAI21X1 U1024 ( .A(n1255), .B(n1325), .C(n1424), .Y(n723) );
  NAND2X1 U1025 ( .A(\mem<27><9> ), .B(n35), .Y(n1425) );
  OAI21X1 U1026 ( .A(n1255), .B(n1327), .C(n1425), .Y(n724) );
  NAND2X1 U1027 ( .A(\mem<27><10> ), .B(n35), .Y(n1426) );
  OAI21X1 U1028 ( .A(n1255), .B(n1329), .C(n1426), .Y(n725) );
  NAND2X1 U1029 ( .A(\mem<27><11> ), .B(n35), .Y(n1427) );
  OAI21X1 U1030 ( .A(n1255), .B(n1331), .C(n1427), .Y(n726) );
  NAND2X1 U1031 ( .A(\mem<27><12> ), .B(n35), .Y(n1428) );
  OAI21X1 U1032 ( .A(n1255), .B(n1333), .C(n1428), .Y(n727) );
  NAND2X1 U1033 ( .A(\mem<27><13> ), .B(n35), .Y(n1429) );
  OAI21X1 U1034 ( .A(n1255), .B(n1335), .C(n1429), .Y(n728) );
  NAND2X1 U1035 ( .A(\mem<27><14> ), .B(n35), .Y(n1430) );
  OAI21X1 U1036 ( .A(n1255), .B(n1229), .C(n1430), .Y(n729) );
  NAND2X1 U1037 ( .A(\mem<27><15> ), .B(n35), .Y(n1431) );
  OAI21X1 U1038 ( .A(n1255), .B(n1338), .C(n1431), .Y(n730) );
  NAND3X1 U1039 ( .A(n1344), .B(n1342), .C(n1341), .Y(n1432) );
  NAND2X1 U1040 ( .A(\mem<26><0> ), .B(n37), .Y(n1433) );
  OAI21X1 U1041 ( .A(n1256), .B(n1310), .C(n1433), .Y(n731) );
  NAND2X1 U1042 ( .A(\mem<26><1> ), .B(n37), .Y(n1434) );
  OAI21X1 U1043 ( .A(n1256), .B(n1313), .C(n1434), .Y(n732) );
  NAND2X1 U1044 ( .A(\mem<26><2> ), .B(n37), .Y(n1435) );
  OAI21X1 U1045 ( .A(n1256), .B(n1315), .C(n1435), .Y(n733) );
  NAND2X1 U1046 ( .A(\mem<26><3> ), .B(n37), .Y(n1436) );
  OAI21X1 U1047 ( .A(n1256), .B(n1317), .C(n1436), .Y(n734) );
  NAND2X1 U1048 ( .A(\mem<26><4> ), .B(n37), .Y(n1437) );
  OAI21X1 U1049 ( .A(n1256), .B(n1319), .C(n1437), .Y(n735) );
  NAND2X1 U1050 ( .A(\mem<26><5> ), .B(n37), .Y(n1438) );
  OAI21X1 U1051 ( .A(n1256), .B(n1321), .C(n1438), .Y(n736) );
  NAND2X1 U1052 ( .A(\mem<26><6> ), .B(n37), .Y(n1439) );
  OAI21X1 U1053 ( .A(n1256), .B(n1323), .C(n1439), .Y(n737) );
  NAND2X1 U1054 ( .A(\mem<26><7> ), .B(n37), .Y(n1440) );
  OAI21X1 U1055 ( .A(n1256), .B(n1244), .C(n1440), .Y(n738) );
  NAND2X1 U1056 ( .A(\mem<26><8> ), .B(n37), .Y(n1441) );
  OAI21X1 U1057 ( .A(n1257), .B(n1325), .C(n1441), .Y(n739) );
  NAND2X1 U1058 ( .A(\mem<26><9> ), .B(n37), .Y(n1442) );
  OAI21X1 U1059 ( .A(n1257), .B(n1327), .C(n1442), .Y(n740) );
  NAND2X1 U1060 ( .A(\mem<26><10> ), .B(n37), .Y(n1443) );
  OAI21X1 U1061 ( .A(n1257), .B(n1329), .C(n1443), .Y(n741) );
  NAND2X1 U1062 ( .A(\mem<26><11> ), .B(n37), .Y(n1444) );
  OAI21X1 U1063 ( .A(n1257), .B(n1331), .C(n1444), .Y(n742) );
  NAND2X1 U1064 ( .A(\mem<26><12> ), .B(n37), .Y(n1445) );
  OAI21X1 U1065 ( .A(n1257), .B(n1333), .C(n1445), .Y(n743) );
  NAND2X1 U1066 ( .A(\mem<26><13> ), .B(n37), .Y(n1446) );
  OAI21X1 U1067 ( .A(n1257), .B(n1335), .C(n1446), .Y(n744) );
  NAND2X1 U1068 ( .A(\mem<26><14> ), .B(n37), .Y(n1447) );
  OAI21X1 U1069 ( .A(n1257), .B(n1226), .C(n1447), .Y(n745) );
  NAND2X1 U1070 ( .A(\mem<26><15> ), .B(n37), .Y(n1448) );
  OAI21X1 U1071 ( .A(n1257), .B(n1338), .C(n1448), .Y(n746) );
  NAND3X1 U1072 ( .A(n1340), .B(n1344), .C(n1343), .Y(n1449) );
  NAND2X1 U1073 ( .A(\mem<25><0> ), .B(n39), .Y(n1450) );
  OAI21X1 U1074 ( .A(n1258), .B(n1310), .C(n1450), .Y(n747) );
  NAND2X1 U1075 ( .A(\mem<25><1> ), .B(n39), .Y(n1451) );
  OAI21X1 U1076 ( .A(n1258), .B(n1313), .C(n1451), .Y(n748) );
  NAND2X1 U1077 ( .A(\mem<25><2> ), .B(n39), .Y(n1452) );
  OAI21X1 U1078 ( .A(n1258), .B(n1315), .C(n1452), .Y(n749) );
  NAND2X1 U1079 ( .A(\mem<25><3> ), .B(n39), .Y(n1453) );
  OAI21X1 U1080 ( .A(n1258), .B(n1317), .C(n1453), .Y(n750) );
  NAND2X1 U1081 ( .A(\mem<25><4> ), .B(n39), .Y(n1454) );
  OAI21X1 U1082 ( .A(n1258), .B(n1319), .C(n1454), .Y(n751) );
  NAND2X1 U1083 ( .A(\mem<25><5> ), .B(n39), .Y(n1455) );
  OAI21X1 U1084 ( .A(n1258), .B(n1321), .C(n1455), .Y(n752) );
  NAND2X1 U1085 ( .A(\mem<25><6> ), .B(n39), .Y(n1456) );
  OAI21X1 U1086 ( .A(n1258), .B(n1323), .C(n1456), .Y(n753) );
  NAND2X1 U1087 ( .A(\mem<25><7> ), .B(n39), .Y(n1457) );
  OAI21X1 U1088 ( .A(n1258), .B(n1242), .C(n1457), .Y(n754) );
  NAND2X1 U1089 ( .A(\mem<25><8> ), .B(n39), .Y(n1458) );
  OAI21X1 U1090 ( .A(n1259), .B(n1325), .C(n1458), .Y(n755) );
  NAND2X1 U1091 ( .A(\mem<25><9> ), .B(n39), .Y(n1459) );
  OAI21X1 U1092 ( .A(n1259), .B(n1327), .C(n1459), .Y(n756) );
  NAND2X1 U1093 ( .A(\mem<25><10> ), .B(n39), .Y(n1460) );
  OAI21X1 U1094 ( .A(n1259), .B(n1329), .C(n1460), .Y(n757) );
  NAND2X1 U1095 ( .A(\mem<25><11> ), .B(n39), .Y(n1461) );
  OAI21X1 U1096 ( .A(n1259), .B(n1331), .C(n1461), .Y(n758) );
  NAND2X1 U1097 ( .A(\mem<25><12> ), .B(n39), .Y(n1462) );
  OAI21X1 U1098 ( .A(n1259), .B(n1333), .C(n1462), .Y(n759) );
  NAND2X1 U1099 ( .A(\mem<25><13> ), .B(n39), .Y(n1463) );
  OAI21X1 U1100 ( .A(n1259), .B(n1335), .C(n1463), .Y(n760) );
  NAND2X1 U1101 ( .A(\mem<25><14> ), .B(n39), .Y(n1464) );
  OAI21X1 U1102 ( .A(n1259), .B(n1225), .C(n1464), .Y(n761) );
  NAND2X1 U1103 ( .A(\mem<25><15> ), .B(n39), .Y(n1465) );
  OAI21X1 U1104 ( .A(n1259), .B(n1338), .C(n1465), .Y(n762) );
  NOR3X1 U1105 ( .A(n1340), .B(n1342), .C(n1179), .Y(n1859) );
  NAND2X1 U1106 ( .A(\mem<24><0> ), .B(n41), .Y(n1466) );
  OAI21X1 U1107 ( .A(n1260), .B(n1310), .C(n1466), .Y(n763) );
  NAND2X1 U1108 ( .A(\mem<24><1> ), .B(n41), .Y(n1467) );
  OAI21X1 U1109 ( .A(n1260), .B(n1313), .C(n1467), .Y(n764) );
  NAND2X1 U1110 ( .A(\mem<24><2> ), .B(n41), .Y(n1468) );
  OAI21X1 U1111 ( .A(n1260), .B(n1315), .C(n1468), .Y(n765) );
  NAND2X1 U1112 ( .A(\mem<24><3> ), .B(n41), .Y(n1469) );
  OAI21X1 U1113 ( .A(n1260), .B(n1317), .C(n1469), .Y(n766) );
  NAND2X1 U1114 ( .A(\mem<24><4> ), .B(n41), .Y(n1470) );
  OAI21X1 U1115 ( .A(n1260), .B(n1319), .C(n1470), .Y(n767) );
  NAND2X1 U1116 ( .A(\mem<24><5> ), .B(n41), .Y(n1471) );
  OAI21X1 U1117 ( .A(n1260), .B(n1321), .C(n1471), .Y(n768) );
  NAND2X1 U1118 ( .A(\mem<24><6> ), .B(n41), .Y(n1472) );
  OAI21X1 U1119 ( .A(n1260), .B(n1323), .C(n1472), .Y(n769) );
  NAND2X1 U1120 ( .A(\mem<24><7> ), .B(n41), .Y(n1473) );
  OAI21X1 U1121 ( .A(n1260), .B(n1242), .C(n1473), .Y(n770) );
  NAND2X1 U1122 ( .A(\mem<24><8> ), .B(n41), .Y(n1474) );
  OAI21X1 U1123 ( .A(n1260), .B(n1325), .C(n1474), .Y(n771) );
  NAND2X1 U1124 ( .A(\mem<24><9> ), .B(n41), .Y(n1475) );
  OAI21X1 U1125 ( .A(n1260), .B(n1327), .C(n1475), .Y(n772) );
  NAND2X1 U1126 ( .A(\mem<24><10> ), .B(n41), .Y(n1476) );
  OAI21X1 U1127 ( .A(n1260), .B(n1329), .C(n1476), .Y(n773) );
  NAND2X1 U1128 ( .A(\mem<24><11> ), .B(n41), .Y(n1477) );
  OAI21X1 U1129 ( .A(n1260), .B(n1331), .C(n1477), .Y(n774) );
  NAND2X1 U1130 ( .A(\mem<24><12> ), .B(n41), .Y(n1478) );
  OAI21X1 U1131 ( .A(n1260), .B(n1333), .C(n1478), .Y(n775) );
  NAND2X1 U1132 ( .A(\mem<24><13> ), .B(n41), .Y(n1479) );
  OAI21X1 U1133 ( .A(n1260), .B(n1335), .C(n1479), .Y(n776) );
  NAND2X1 U1134 ( .A(\mem<24><14> ), .B(n41), .Y(n1480) );
  OAI21X1 U1135 ( .A(n1260), .B(n1227), .C(n1480), .Y(n777) );
  NAND2X1 U1136 ( .A(\mem<24><15> ), .B(n41), .Y(n1481) );
  OAI21X1 U1137 ( .A(n1260), .B(n1338), .C(n1481), .Y(n778) );
  NAND2X1 U1138 ( .A(\mem<23><0> ), .B(n43), .Y(n1482) );
  OAI21X1 U1139 ( .A(n1261), .B(n1310), .C(n1482), .Y(n779) );
  NAND2X1 U1140 ( .A(\mem<23><1> ), .B(n43), .Y(n1483) );
  OAI21X1 U1141 ( .A(n1261), .B(n1313), .C(n1483), .Y(n780) );
  NAND2X1 U1142 ( .A(\mem<23><2> ), .B(n43), .Y(n1484) );
  OAI21X1 U1143 ( .A(n1261), .B(n1315), .C(n1484), .Y(n781) );
  NAND2X1 U1144 ( .A(\mem<23><3> ), .B(n43), .Y(n1485) );
  OAI21X1 U1145 ( .A(n1261), .B(n1317), .C(n1485), .Y(n782) );
  NAND2X1 U1146 ( .A(\mem<23><4> ), .B(n43), .Y(n1486) );
  OAI21X1 U1147 ( .A(n1261), .B(n1319), .C(n1486), .Y(n783) );
  NAND2X1 U1148 ( .A(\mem<23><5> ), .B(n43), .Y(n1487) );
  OAI21X1 U1149 ( .A(n1261), .B(n1321), .C(n1487), .Y(n784) );
  NAND2X1 U1150 ( .A(\mem<23><6> ), .B(n43), .Y(n1488) );
  OAI21X1 U1151 ( .A(n1261), .B(n1323), .C(n1488), .Y(n785) );
  NAND2X1 U1152 ( .A(\mem<23><7> ), .B(n43), .Y(n1489) );
  OAI21X1 U1153 ( .A(n1261), .B(n1238), .C(n1489), .Y(n786) );
  NAND2X1 U1154 ( .A(\mem<23><8> ), .B(n43), .Y(n1490) );
  OAI21X1 U1155 ( .A(n1262), .B(n1325), .C(n1490), .Y(n787) );
  NAND2X1 U1156 ( .A(\mem<23><9> ), .B(n43), .Y(n1491) );
  OAI21X1 U1157 ( .A(n1262), .B(n1327), .C(n1491), .Y(n788) );
  NAND2X1 U1158 ( .A(\mem<23><10> ), .B(n43), .Y(n1492) );
  OAI21X1 U1159 ( .A(n1262), .B(n1329), .C(n1492), .Y(n789) );
  NAND2X1 U1160 ( .A(\mem<23><11> ), .B(n43), .Y(n1493) );
  OAI21X1 U1161 ( .A(n1262), .B(n1331), .C(n1493), .Y(n790) );
  NAND2X1 U1162 ( .A(\mem<23><12> ), .B(n43), .Y(n1494) );
  OAI21X1 U1163 ( .A(n1262), .B(n1333), .C(n1494), .Y(n791) );
  NAND2X1 U1164 ( .A(\mem<23><13> ), .B(n43), .Y(n1495) );
  OAI21X1 U1165 ( .A(n1262), .B(n1335), .C(n1495), .Y(n792) );
  NAND2X1 U1166 ( .A(\mem<23><14> ), .B(n43), .Y(n1496) );
  OAI21X1 U1167 ( .A(n1262), .B(n1222), .C(n1496), .Y(n793) );
  NAND2X1 U1168 ( .A(\mem<23><15> ), .B(n43), .Y(n1497) );
  OAI21X1 U1169 ( .A(n1262), .B(n1338), .C(n1497), .Y(n794) );
  NAND2X1 U1170 ( .A(\mem<22><0> ), .B(n19), .Y(n1498) );
  OAI21X1 U1171 ( .A(n1263), .B(n1310), .C(n1498), .Y(n795) );
  NAND2X1 U1172 ( .A(\mem<22><1> ), .B(n19), .Y(n1499) );
  OAI21X1 U1173 ( .A(n1263), .B(n1313), .C(n1499), .Y(n796) );
  NAND2X1 U1174 ( .A(\mem<22><2> ), .B(n19), .Y(n1500) );
  OAI21X1 U1175 ( .A(n1263), .B(n1315), .C(n1500), .Y(n797) );
  NAND2X1 U1177 ( .A(\mem<22><3> ), .B(n19), .Y(n1501) );
  OAI21X1 U1178 ( .A(n1263), .B(n1317), .C(n1501), .Y(n798) );
  NAND2X1 U1179 ( .A(\mem<22><4> ), .B(n19), .Y(n1502) );
  OAI21X1 U1180 ( .A(n1263), .B(n1319), .C(n1502), .Y(n799) );
  NAND2X1 U1181 ( .A(\mem<22><5> ), .B(n19), .Y(n1503) );
  OAI21X1 U1182 ( .A(n1263), .B(n1321), .C(n1503), .Y(n800) );
  NAND2X1 U1183 ( .A(\mem<22><6> ), .B(n19), .Y(n1504) );
  OAI21X1 U1184 ( .A(n1263), .B(n1323), .C(n1504), .Y(n801) );
  NAND2X1 U1185 ( .A(\mem<22><7> ), .B(n19), .Y(n1505) );
  OAI21X1 U1186 ( .A(n1263), .B(n1239), .C(n1505), .Y(n802) );
  NAND2X1 U1187 ( .A(\mem<22><8> ), .B(n19), .Y(n1506) );
  OAI21X1 U1188 ( .A(n1264), .B(n1325), .C(n1506), .Y(n803) );
  NAND2X1 U1189 ( .A(\mem<22><9> ), .B(n19), .Y(n1507) );
  OAI21X1 U1190 ( .A(n1264), .B(n1327), .C(n1507), .Y(n804) );
  NAND2X1 U1191 ( .A(\mem<22><10> ), .B(n19), .Y(n1508) );
  OAI21X1 U1192 ( .A(n1264), .B(n1329), .C(n1508), .Y(n805) );
  NAND2X1 U1193 ( .A(\mem<22><11> ), .B(n19), .Y(n1509) );
  OAI21X1 U1194 ( .A(n1264), .B(n1331), .C(n1509), .Y(n806) );
  NAND2X1 U1195 ( .A(\mem<22><12> ), .B(n19), .Y(n1510) );
  OAI21X1 U1196 ( .A(n1264), .B(n1333), .C(n1510), .Y(n807) );
  NAND2X1 U1197 ( .A(\mem<22><13> ), .B(n19), .Y(n1511) );
  OAI21X1 U1198 ( .A(n1264), .B(n1335), .C(n1511), .Y(n808) );
  NAND2X1 U1199 ( .A(\mem<22><14> ), .B(n19), .Y(n1512) );
  OAI21X1 U1200 ( .A(n1264), .B(n1223), .C(n1512), .Y(n809) );
  NAND2X1 U1201 ( .A(\mem<22><15> ), .B(n19), .Y(n1513) );
  OAI21X1 U1202 ( .A(n1264), .B(n1338), .C(n1513), .Y(n810) );
  NAND2X1 U1203 ( .A(\mem<21><0> ), .B(n45), .Y(n1514) );
  OAI21X1 U1204 ( .A(n1265), .B(n1310), .C(n1514), .Y(n811) );
  NAND2X1 U1205 ( .A(\mem<21><1> ), .B(n45), .Y(n1515) );
  OAI21X1 U1206 ( .A(n1265), .B(n1313), .C(n1515), .Y(n812) );
  NAND2X1 U1207 ( .A(\mem<21><2> ), .B(n45), .Y(n1516) );
  OAI21X1 U1208 ( .A(n1265), .B(n1315), .C(n1516), .Y(n813) );
  NAND2X1 U1209 ( .A(\mem<21><3> ), .B(n45), .Y(n1517) );
  OAI21X1 U1210 ( .A(n1265), .B(n1317), .C(n1517), .Y(n814) );
  NAND2X1 U1211 ( .A(\mem<21><4> ), .B(n45), .Y(n1518) );
  OAI21X1 U1212 ( .A(n1265), .B(n1319), .C(n1518), .Y(n815) );
  NAND2X1 U1213 ( .A(\mem<21><5> ), .B(n45), .Y(n1519) );
  OAI21X1 U1214 ( .A(n1265), .B(n1321), .C(n1519), .Y(n816) );
  NAND2X1 U1215 ( .A(\mem<21><6> ), .B(n45), .Y(n1520) );
  OAI21X1 U1216 ( .A(n1265), .B(n1323), .C(n1520), .Y(n817) );
  NAND2X1 U1217 ( .A(\mem<21><7> ), .B(n45), .Y(n1521) );
  OAI21X1 U1218 ( .A(n1265), .B(n1243), .C(n1521), .Y(n818) );
  NAND2X1 U1219 ( .A(\mem<21><8> ), .B(n45), .Y(n1522) );
  OAI21X1 U1220 ( .A(n1266), .B(n1325), .C(n1522), .Y(n819) );
  NAND2X1 U1221 ( .A(\mem<21><9> ), .B(n45), .Y(n1523) );
  OAI21X1 U1222 ( .A(n1266), .B(n1327), .C(n1523), .Y(n820) );
  NAND2X1 U1223 ( .A(\mem<21><10> ), .B(n45), .Y(n1524) );
  OAI21X1 U1224 ( .A(n1266), .B(n1329), .C(n1524), .Y(n821) );
  NAND2X1 U1225 ( .A(\mem<21><11> ), .B(n45), .Y(n1525) );
  OAI21X1 U1226 ( .A(n1266), .B(n1331), .C(n1525), .Y(n822) );
  NAND2X1 U1227 ( .A(\mem<21><12> ), .B(n45), .Y(n1526) );
  OAI21X1 U1228 ( .A(n1266), .B(n1333), .C(n1526), .Y(n823) );
  NAND2X1 U1229 ( .A(\mem<21><13> ), .B(n45), .Y(n1527) );
  OAI21X1 U1230 ( .A(n1266), .B(n1335), .C(n1527), .Y(n824) );
  NAND2X1 U1231 ( .A(\mem<21><14> ), .B(n45), .Y(n1528) );
  OAI21X1 U1232 ( .A(n1266), .B(n1224), .C(n1528), .Y(n825) );
  NAND2X1 U1233 ( .A(\mem<21><15> ), .B(n45), .Y(n1529) );
  OAI21X1 U1234 ( .A(n1266), .B(n1338), .C(n1529), .Y(n826) );
  NAND2X1 U1235 ( .A(\mem<20><0> ), .B(n21), .Y(n1530) );
  OAI21X1 U1236 ( .A(n1267), .B(n1310), .C(n1530), .Y(n827) );
  NAND2X1 U1237 ( .A(\mem<20><1> ), .B(n21), .Y(n1531) );
  OAI21X1 U1238 ( .A(n1267), .B(n1313), .C(n1531), .Y(n828) );
  NAND2X1 U1239 ( .A(\mem<20><2> ), .B(n21), .Y(n1532) );
  OAI21X1 U1240 ( .A(n1267), .B(n1315), .C(n1532), .Y(n829) );
  NAND2X1 U1241 ( .A(\mem<20><3> ), .B(n21), .Y(n1533) );
  OAI21X1 U1242 ( .A(n1267), .B(n1317), .C(n1533), .Y(n830) );
  NAND2X1 U1243 ( .A(\mem<20><4> ), .B(n21), .Y(n1534) );
  OAI21X1 U1244 ( .A(n1267), .B(n1319), .C(n1534), .Y(n831) );
  NAND2X1 U1245 ( .A(\mem<20><5> ), .B(n21), .Y(n1535) );
  OAI21X1 U1246 ( .A(n1267), .B(n1321), .C(n1535), .Y(n832) );
  NAND2X1 U1247 ( .A(\mem<20><6> ), .B(n21), .Y(n1536) );
  OAI21X1 U1248 ( .A(n1267), .B(n1323), .C(n1536), .Y(n833) );
  NAND2X1 U1249 ( .A(\mem<20><7> ), .B(n21), .Y(n1537) );
  OAI21X1 U1250 ( .A(n1267), .B(n1242), .C(n1537), .Y(n834) );
  NAND2X1 U1251 ( .A(\mem<20><8> ), .B(n21), .Y(n1538) );
  OAI21X1 U1252 ( .A(n1268), .B(n1325), .C(n1538), .Y(n835) );
  NAND2X1 U1253 ( .A(\mem<20><9> ), .B(n21), .Y(n1539) );
  OAI21X1 U1254 ( .A(n1268), .B(n1327), .C(n1539), .Y(n836) );
  NAND2X1 U1255 ( .A(\mem<20><10> ), .B(n21), .Y(n1540) );
  OAI21X1 U1256 ( .A(n1268), .B(n1329), .C(n1540), .Y(n837) );
  NAND2X1 U1257 ( .A(\mem<20><11> ), .B(n21), .Y(n1541) );
  OAI21X1 U1258 ( .A(n1268), .B(n1331), .C(n1541), .Y(n838) );
  NAND2X1 U1259 ( .A(\mem<20><12> ), .B(n21), .Y(n1542) );
  OAI21X1 U1260 ( .A(n1268), .B(n1333), .C(n1542), .Y(n839) );
  NAND2X1 U1261 ( .A(\mem<20><13> ), .B(n21), .Y(n1543) );
  OAI21X1 U1262 ( .A(n1268), .B(n1335), .C(n1543), .Y(n840) );
  NAND2X1 U1263 ( .A(\mem<20><14> ), .B(n21), .Y(n1544) );
  OAI21X1 U1264 ( .A(n1268), .B(n1226), .C(n1544), .Y(n841) );
  NAND2X1 U1265 ( .A(\mem<20><15> ), .B(n21), .Y(n1545) );
  OAI21X1 U1266 ( .A(n1268), .B(n1338), .C(n1545), .Y(n842) );
  NAND2X1 U1267 ( .A(\mem<19><0> ), .B(n47), .Y(n1546) );
  OAI21X1 U1268 ( .A(n1269), .B(n1310), .C(n1546), .Y(n843) );
  NAND2X1 U1269 ( .A(\mem<19><1> ), .B(n47), .Y(n1547) );
  OAI21X1 U1270 ( .A(n1269), .B(n1312), .C(n1547), .Y(n844) );
  NAND2X1 U1271 ( .A(\mem<19><2> ), .B(n47), .Y(n1548) );
  OAI21X1 U1272 ( .A(n1269), .B(n1314), .C(n1548), .Y(n845) );
  NAND2X1 U1273 ( .A(\mem<19><3> ), .B(n47), .Y(n1549) );
  OAI21X1 U1274 ( .A(n1269), .B(n1316), .C(n1549), .Y(n846) );
  NAND2X1 U1275 ( .A(\mem<19><4> ), .B(n47), .Y(n1550) );
  OAI21X1 U1276 ( .A(n1269), .B(n1318), .C(n1550), .Y(n847) );
  NAND2X1 U1277 ( .A(\mem<19><5> ), .B(n47), .Y(n1551) );
  OAI21X1 U1278 ( .A(n1269), .B(n1320), .C(n1551), .Y(n848) );
  NAND2X1 U1279 ( .A(\mem<19><6> ), .B(n47), .Y(n1552) );
  OAI21X1 U1280 ( .A(n1269), .B(n1322), .C(n1552), .Y(n849) );
  NAND2X1 U1281 ( .A(\mem<19><7> ), .B(n47), .Y(n1553) );
  OAI21X1 U1282 ( .A(n1269), .B(n1243), .C(n1553), .Y(n850) );
  NAND2X1 U1283 ( .A(\mem<19><8> ), .B(n47), .Y(n1554) );
  OAI21X1 U1284 ( .A(n1270), .B(n1325), .C(n1554), .Y(n851) );
  NAND2X1 U1285 ( .A(\mem<19><9> ), .B(n47), .Y(n1555) );
  OAI21X1 U1286 ( .A(n1270), .B(n1327), .C(n1555), .Y(n852) );
  NAND2X1 U1287 ( .A(\mem<19><10> ), .B(n47), .Y(n1556) );
  OAI21X1 U1288 ( .A(n1270), .B(n1329), .C(n1556), .Y(n853) );
  NAND2X1 U1289 ( .A(\mem<19><11> ), .B(n47), .Y(n1557) );
  OAI21X1 U1290 ( .A(n1270), .B(n1331), .C(n1557), .Y(n854) );
  NAND2X1 U1291 ( .A(\mem<19><12> ), .B(n47), .Y(n1558) );
  OAI21X1 U1292 ( .A(n1270), .B(n1333), .C(n1558), .Y(n855) );
  NAND2X1 U1293 ( .A(\mem<19><13> ), .B(n47), .Y(n1559) );
  OAI21X1 U1294 ( .A(n1270), .B(n1335), .C(n1559), .Y(n856) );
  NAND2X1 U1295 ( .A(\mem<19><14> ), .B(n47), .Y(n1560) );
  OAI21X1 U1296 ( .A(n1270), .B(n1226), .C(n1560), .Y(n857) );
  NAND2X1 U1297 ( .A(\mem<19><15> ), .B(n47), .Y(n1561) );
  OAI21X1 U1298 ( .A(n1270), .B(n1338), .C(n1561), .Y(n858) );
  NAND2X1 U1299 ( .A(\mem<18><0> ), .B(n49), .Y(n1562) );
  OAI21X1 U1300 ( .A(n1271), .B(n1311), .C(n1562), .Y(n859) );
  NAND2X1 U1301 ( .A(\mem<18><1> ), .B(n49), .Y(n1563) );
  OAI21X1 U1302 ( .A(n1271), .B(n1313), .C(n1563), .Y(n860) );
  NAND2X1 U1303 ( .A(\mem<18><2> ), .B(n49), .Y(n1564) );
  OAI21X1 U1304 ( .A(n1271), .B(n1315), .C(n1564), .Y(n861) );
  NAND2X1 U1305 ( .A(\mem<18><3> ), .B(n49), .Y(n1565) );
  OAI21X1 U1306 ( .A(n1271), .B(n1317), .C(n1565), .Y(n862) );
  NAND2X1 U1307 ( .A(\mem<18><4> ), .B(n49), .Y(n1566) );
  OAI21X1 U1308 ( .A(n1271), .B(n1319), .C(n1566), .Y(n863) );
  NAND2X1 U1309 ( .A(\mem<18><5> ), .B(n49), .Y(n1567) );
  OAI21X1 U1310 ( .A(n1271), .B(n1321), .C(n1567), .Y(n864) );
  NAND2X1 U1311 ( .A(\mem<18><6> ), .B(n49), .Y(n1568) );
  OAI21X1 U1312 ( .A(n1271), .B(n1323), .C(n1568), .Y(n865) );
  NAND2X1 U1313 ( .A(\mem<18><7> ), .B(n49), .Y(n1569) );
  OAI21X1 U1314 ( .A(n1271), .B(n1244), .C(n1569), .Y(n866) );
  NAND2X1 U1315 ( .A(\mem<18><8> ), .B(n49), .Y(n1570) );
  OAI21X1 U1316 ( .A(n1272), .B(n1324), .C(n1570), .Y(n867) );
  NAND2X1 U1317 ( .A(\mem<18><9> ), .B(n49), .Y(n1571) );
  OAI21X1 U1318 ( .A(n1272), .B(n1326), .C(n1571), .Y(n868) );
  NAND2X1 U1319 ( .A(\mem<18><10> ), .B(n49), .Y(n1572) );
  OAI21X1 U1320 ( .A(n1272), .B(n1328), .C(n1572), .Y(n869) );
  NAND2X1 U1321 ( .A(\mem<18><11> ), .B(n49), .Y(n1573) );
  OAI21X1 U1322 ( .A(n1272), .B(n1330), .C(n1573), .Y(n870) );
  NAND2X1 U1323 ( .A(\mem<18><12> ), .B(n49), .Y(n1574) );
  OAI21X1 U1324 ( .A(n1272), .B(n1332), .C(n1574), .Y(n871) );
  NAND2X1 U1325 ( .A(\mem<18><13> ), .B(n49), .Y(n1575) );
  OAI21X1 U1326 ( .A(n1272), .B(n1334), .C(n1575), .Y(n872) );
  NAND2X1 U1327 ( .A(\mem<18><14> ), .B(n49), .Y(n1576) );
  OAI21X1 U1328 ( .A(n1272), .B(n1226), .C(n1576), .Y(n873) );
  NAND2X1 U1329 ( .A(\mem<18><15> ), .B(n49), .Y(n1577) );
  OAI21X1 U1330 ( .A(n1272), .B(n1337), .C(n1577), .Y(n874) );
  NAND2X1 U1331 ( .A(\mem<17><0> ), .B(n51), .Y(n1578) );
  OAI21X1 U1332 ( .A(n1273), .B(n1310), .C(n1578), .Y(n875) );
  NAND2X1 U1333 ( .A(\mem<17><1> ), .B(n51), .Y(n1579) );
  OAI21X1 U1334 ( .A(n1273), .B(n1312), .C(n1579), .Y(n876) );
  NAND2X1 U1335 ( .A(\mem<17><2> ), .B(n51), .Y(n1580) );
  OAI21X1 U1336 ( .A(n1273), .B(n1314), .C(n1580), .Y(n877) );
  NAND2X1 U1337 ( .A(\mem<17><3> ), .B(n51), .Y(n1581) );
  OAI21X1 U1338 ( .A(n1273), .B(n1316), .C(n1581), .Y(n878) );
  NAND2X1 U1339 ( .A(\mem<17><4> ), .B(n51), .Y(n1582) );
  OAI21X1 U1340 ( .A(n1273), .B(n1318), .C(n1582), .Y(n879) );
  NAND2X1 U1341 ( .A(\mem<17><5> ), .B(n51), .Y(n1583) );
  OAI21X1 U1342 ( .A(n1273), .B(n1320), .C(n1583), .Y(n880) );
  NAND2X1 U1343 ( .A(\mem<17><6> ), .B(n51), .Y(n1584) );
  OAI21X1 U1344 ( .A(n1273), .B(n1322), .C(n1584), .Y(n881) );
  NAND2X1 U1345 ( .A(\mem<17><7> ), .B(n51), .Y(n1585) );
  OAI21X1 U1346 ( .A(n1273), .B(n1238), .C(n1585), .Y(n882) );
  NAND2X1 U1347 ( .A(\mem<17><8> ), .B(n51), .Y(n1586) );
  OAI21X1 U1348 ( .A(n1274), .B(n1325), .C(n1586), .Y(n883) );
  NAND2X1 U1349 ( .A(\mem<17><9> ), .B(n51), .Y(n1587) );
  OAI21X1 U1350 ( .A(n1274), .B(n1327), .C(n1587), .Y(n884) );
  NAND2X1 U1351 ( .A(\mem<17><10> ), .B(n51), .Y(n1588) );
  OAI21X1 U1352 ( .A(n1274), .B(n1329), .C(n1588), .Y(n885) );
  NAND2X1 U1353 ( .A(\mem<17><11> ), .B(n51), .Y(n1589) );
  OAI21X1 U1354 ( .A(n1274), .B(n1331), .C(n1589), .Y(n886) );
  NAND2X1 U1355 ( .A(\mem<17><12> ), .B(n51), .Y(n1590) );
  OAI21X1 U1356 ( .A(n1274), .B(n1333), .C(n1590), .Y(n887) );
  NAND2X1 U1357 ( .A(\mem<17><13> ), .B(n51), .Y(n1591) );
  OAI21X1 U1358 ( .A(n1274), .B(n1335), .C(n1591), .Y(n888) );
  NAND2X1 U1359 ( .A(\mem<17><14> ), .B(n51), .Y(n1592) );
  OAI21X1 U1360 ( .A(n1274), .B(n1225), .C(n1592), .Y(n889) );
  NAND2X1 U1361 ( .A(\mem<17><15> ), .B(n51), .Y(n1593) );
  OAI21X1 U1362 ( .A(n1274), .B(n1338), .C(n1593), .Y(n890) );
  NAND2X1 U1363 ( .A(\mem<16><0> ), .B(n53), .Y(n1594) );
  OAI21X1 U1364 ( .A(n1275), .B(n1311), .C(n1594), .Y(n891) );
  NAND2X1 U1365 ( .A(\mem<16><1> ), .B(n53), .Y(n1595) );
  OAI21X1 U1366 ( .A(n1275), .B(n1313), .C(n1595), .Y(n892) );
  NAND2X1 U1367 ( .A(\mem<16><2> ), .B(n53), .Y(n1596) );
  OAI21X1 U1368 ( .A(n1275), .B(n1315), .C(n1596), .Y(n893) );
  NAND2X1 U1369 ( .A(\mem<16><3> ), .B(n53), .Y(n1597) );
  OAI21X1 U1370 ( .A(n1275), .B(n1317), .C(n1597), .Y(n894) );
  NAND2X1 U1371 ( .A(\mem<16><4> ), .B(n53), .Y(n1598) );
  OAI21X1 U1372 ( .A(n1275), .B(n1319), .C(n1598), .Y(n895) );
  NAND2X1 U1373 ( .A(\mem<16><5> ), .B(n53), .Y(n1599) );
  OAI21X1 U1374 ( .A(n1275), .B(n1321), .C(n1599), .Y(n896) );
  NAND2X1 U1375 ( .A(\mem<16><6> ), .B(n53), .Y(n1600) );
  OAI21X1 U1376 ( .A(n1275), .B(n1323), .C(n1600), .Y(n897) );
  NAND2X1 U1377 ( .A(\mem<16><7> ), .B(n53), .Y(n1601) );
  OAI21X1 U1378 ( .A(n1275), .B(n1242), .C(n1601), .Y(n898) );
  NAND2X1 U1379 ( .A(\mem<16><8> ), .B(n53), .Y(n1602) );
  OAI21X1 U1380 ( .A(n1275), .B(n1324), .C(n1602), .Y(n899) );
  NAND2X1 U1381 ( .A(\mem<16><9> ), .B(n53), .Y(n1603) );
  OAI21X1 U1382 ( .A(n1275), .B(n1326), .C(n1603), .Y(n900) );
  NAND2X1 U1383 ( .A(\mem<16><10> ), .B(n53), .Y(n1604) );
  OAI21X1 U1384 ( .A(n1275), .B(n1328), .C(n1604), .Y(n901) );
  NAND2X1 U1385 ( .A(\mem<16><11> ), .B(n53), .Y(n1605) );
  OAI21X1 U1386 ( .A(n1275), .B(n1330), .C(n1605), .Y(n902) );
  NAND2X1 U1387 ( .A(\mem<16><12> ), .B(n53), .Y(n1606) );
  OAI21X1 U1388 ( .A(n1275), .B(n1332), .C(n1606), .Y(n903) );
  NAND2X1 U1389 ( .A(\mem<16><13> ), .B(n53), .Y(n1607) );
  OAI21X1 U1390 ( .A(n1275), .B(n1334), .C(n1607), .Y(n904) );
  NAND2X1 U1391 ( .A(\mem<16><14> ), .B(n53), .Y(n1608) );
  OAI21X1 U1392 ( .A(n1275), .B(n1236), .C(n1608), .Y(n905) );
  NAND2X1 U1393 ( .A(\mem<16><15> ), .B(n53), .Y(n1609) );
  OAI21X1 U1394 ( .A(n1275), .B(n1337), .C(n1609), .Y(n906) );
  NAND3X1 U1395 ( .A(n1345), .B(n214), .C(n1348), .Y(n1610) );
  NAND2X1 U1396 ( .A(\mem<15><0> ), .B(n55), .Y(n1611) );
  OAI21X1 U1397 ( .A(n1276), .B(n1311), .C(n1611), .Y(n907) );
  NAND2X1 U1398 ( .A(\mem<15><1> ), .B(n55), .Y(n1612) );
  OAI21X1 U1399 ( .A(n1276), .B(n1313), .C(n1612), .Y(n908) );
  NAND2X1 U1400 ( .A(\mem<15><2> ), .B(n55), .Y(n1613) );
  OAI21X1 U1401 ( .A(n1276), .B(n1315), .C(n1613), .Y(n909) );
  NAND2X1 U1402 ( .A(\mem<15><3> ), .B(n55), .Y(n1614) );
  OAI21X1 U1403 ( .A(n1276), .B(n1317), .C(n1614), .Y(n910) );
  NAND2X1 U1404 ( .A(\mem<15><4> ), .B(n55), .Y(n1615) );
  OAI21X1 U1405 ( .A(n1276), .B(n1319), .C(n1615), .Y(n911) );
  NAND2X1 U1406 ( .A(\mem<15><5> ), .B(n55), .Y(n1616) );
  OAI21X1 U1407 ( .A(n1276), .B(n1321), .C(n1616), .Y(n912) );
  NAND2X1 U1408 ( .A(\mem<15><6> ), .B(n55), .Y(n1617) );
  OAI21X1 U1409 ( .A(n1276), .B(n1323), .C(n1617), .Y(n913) );
  NAND2X1 U1410 ( .A(\mem<15><7> ), .B(n55), .Y(n1618) );
  OAI21X1 U1411 ( .A(n1276), .B(n1238), .C(n1618), .Y(n914) );
  NAND2X1 U1412 ( .A(\mem<15><8> ), .B(n55), .Y(n1619) );
  OAI21X1 U1413 ( .A(n1277), .B(n1324), .C(n1619), .Y(n915) );
  NAND2X1 U1414 ( .A(\mem<15><9> ), .B(n55), .Y(n1620) );
  OAI21X1 U1415 ( .A(n1277), .B(n1326), .C(n1620), .Y(n916) );
  NAND2X1 U1416 ( .A(\mem<15><10> ), .B(n55), .Y(n1621) );
  OAI21X1 U1417 ( .A(n1277), .B(n1328), .C(n1621), .Y(n917) );
  NAND2X1 U1418 ( .A(\mem<15><11> ), .B(n55), .Y(n1622) );
  OAI21X1 U1419 ( .A(n1277), .B(n1330), .C(n1622), .Y(n918) );
  NAND2X1 U1420 ( .A(\mem<15><12> ), .B(n55), .Y(n1623) );
  OAI21X1 U1421 ( .A(n1277), .B(n1332), .C(n1623), .Y(n919) );
  NAND2X1 U1422 ( .A(\mem<15><13> ), .B(n55), .Y(n1624) );
  OAI21X1 U1423 ( .A(n1277), .B(n1334), .C(n1624), .Y(n920) );
  NAND2X1 U1424 ( .A(\mem<15><14> ), .B(n55), .Y(n1625) );
  OAI21X1 U1425 ( .A(n1277), .B(n1223), .C(n1625), .Y(n921) );
  NAND2X1 U1426 ( .A(\mem<15><15> ), .B(n55), .Y(n1626) );
  OAI21X1 U1427 ( .A(n1277), .B(n1337), .C(n1626), .Y(n922) );
  NAND2X1 U1428 ( .A(\mem<14><0> ), .B(n57), .Y(n1627) );
  OAI21X1 U1429 ( .A(n1278), .B(n1310), .C(n1627), .Y(n923) );
  NAND2X1 U1430 ( .A(\mem<14><1> ), .B(n57), .Y(n1628) );
  OAI21X1 U1431 ( .A(n1278), .B(n1312), .C(n1628), .Y(n924) );
  NAND2X1 U1432 ( .A(\mem<14><2> ), .B(n57), .Y(n1629) );
  OAI21X1 U1433 ( .A(n1278), .B(n1314), .C(n1629), .Y(n925) );
  NAND2X1 U1434 ( .A(\mem<14><3> ), .B(n57), .Y(n1630) );
  OAI21X1 U1435 ( .A(n1278), .B(n1316), .C(n1630), .Y(n926) );
  NAND2X1 U1436 ( .A(\mem<14><4> ), .B(n57), .Y(n1631) );
  OAI21X1 U1437 ( .A(n1278), .B(n1318), .C(n1631), .Y(n927) );
  NAND2X1 U1438 ( .A(\mem<14><5> ), .B(n57), .Y(n1632) );
  OAI21X1 U1439 ( .A(n1278), .B(n1320), .C(n1632), .Y(n928) );
  NAND2X1 U1440 ( .A(\mem<14><6> ), .B(n57), .Y(n1633) );
  OAI21X1 U1441 ( .A(n1278), .B(n1322), .C(n1633), .Y(n929) );
  NAND2X1 U1442 ( .A(\mem<14><7> ), .B(n57), .Y(n1634) );
  OAI21X1 U1443 ( .A(n1278), .B(n1239), .C(n1634), .Y(n930) );
  NAND2X1 U1444 ( .A(\mem<14><8> ), .B(n57), .Y(n1635) );
  OAI21X1 U1445 ( .A(n1279), .B(n1325), .C(n1635), .Y(n931) );
  NAND2X1 U1446 ( .A(\mem<14><9> ), .B(n57), .Y(n1636) );
  OAI21X1 U1447 ( .A(n1279), .B(n1327), .C(n1636), .Y(n932) );
  NAND2X1 U1448 ( .A(\mem<14><10> ), .B(n57), .Y(n1637) );
  OAI21X1 U1449 ( .A(n1279), .B(n1329), .C(n1637), .Y(n933) );
  NAND2X1 U1450 ( .A(\mem<14><11> ), .B(n57), .Y(n1638) );
  OAI21X1 U1451 ( .A(n1279), .B(n1331), .C(n1638), .Y(n934) );
  NAND2X1 U1452 ( .A(\mem<14><12> ), .B(n57), .Y(n1639) );
  OAI21X1 U1453 ( .A(n1279), .B(n1333), .C(n1639), .Y(n935) );
  NAND2X1 U1454 ( .A(\mem<14><13> ), .B(n57), .Y(n1640) );
  OAI21X1 U1455 ( .A(n1279), .B(n1335), .C(n1640), .Y(n936) );
  NAND2X1 U1456 ( .A(\mem<14><14> ), .B(n57), .Y(n1641) );
  OAI21X1 U1457 ( .A(n1279), .B(n1224), .C(n1641), .Y(n937) );
  NAND2X1 U1458 ( .A(\mem<14><15> ), .B(n57), .Y(n1642) );
  OAI21X1 U1459 ( .A(n1279), .B(n1338), .C(n1642), .Y(n938) );
  NAND2X1 U1460 ( .A(\mem<13><0> ), .B(n59), .Y(n1643) );
  OAI21X1 U1461 ( .A(n1280), .B(n1311), .C(n1643), .Y(n939) );
  NAND2X1 U1462 ( .A(\mem<13><1> ), .B(n59), .Y(n1644) );
  OAI21X1 U1463 ( .A(n1280), .B(n1313), .C(n1644), .Y(n940) );
  NAND2X1 U1464 ( .A(\mem<13><2> ), .B(n59), .Y(n1645) );
  OAI21X1 U1465 ( .A(n1280), .B(n1315), .C(n1645), .Y(n941) );
  NAND2X1 U1466 ( .A(\mem<13><3> ), .B(n59), .Y(n1646) );
  OAI21X1 U1467 ( .A(n1280), .B(n1317), .C(n1646), .Y(n942) );
  NAND2X1 U1468 ( .A(\mem<13><4> ), .B(n59), .Y(n1647) );
  OAI21X1 U1469 ( .A(n1280), .B(n1319), .C(n1647), .Y(n943) );
  NAND2X1 U1470 ( .A(\mem<13><5> ), .B(n59), .Y(n1648) );
  OAI21X1 U1471 ( .A(n1280), .B(n1321), .C(n1648), .Y(n944) );
  NAND2X1 U1472 ( .A(\mem<13><6> ), .B(n59), .Y(n1649) );
  OAI21X1 U1473 ( .A(n1280), .B(n1323), .C(n1649), .Y(n945) );
  NAND2X1 U1474 ( .A(\mem<13><7> ), .B(n59), .Y(n1650) );
  OAI21X1 U1475 ( .A(n1280), .B(n1240), .C(n1650), .Y(n946) );
  NAND2X1 U1476 ( .A(\mem<13><8> ), .B(n59), .Y(n1651) );
  OAI21X1 U1477 ( .A(n1281), .B(n1324), .C(n1651), .Y(n947) );
  NAND2X1 U1478 ( .A(\mem<13><9> ), .B(n59), .Y(n1652) );
  OAI21X1 U1479 ( .A(n1281), .B(n1326), .C(n1652), .Y(n948) );
  NAND2X1 U1480 ( .A(\mem<13><10> ), .B(n59), .Y(n1653) );
  OAI21X1 U1481 ( .A(n1281), .B(n1328), .C(n1653), .Y(n949) );
  NAND2X1 U1482 ( .A(\mem<13><11> ), .B(n59), .Y(n1654) );
  OAI21X1 U1483 ( .A(n1281), .B(n1330), .C(n1654), .Y(n950) );
  NAND2X1 U1484 ( .A(\mem<13><12> ), .B(n59), .Y(n1655) );
  OAI21X1 U1485 ( .A(n1281), .B(n1332), .C(n1655), .Y(n951) );
  NAND2X1 U1486 ( .A(\mem<13><13> ), .B(n59), .Y(n1656) );
  OAI21X1 U1487 ( .A(n1281), .B(n1334), .C(n1656), .Y(n952) );
  NAND2X1 U1488 ( .A(\mem<13><14> ), .B(n59), .Y(n1657) );
  OAI21X1 U1489 ( .A(n1281), .B(n1224), .C(n1657), .Y(n953) );
  NAND2X1 U1490 ( .A(\mem<13><15> ), .B(n59), .Y(n1658) );
  OAI21X1 U1491 ( .A(n1281), .B(n1337), .C(n1658), .Y(n954) );
  NAND2X1 U1492 ( .A(\mem<12><0> ), .B(n61), .Y(n1659) );
  OAI21X1 U1493 ( .A(n1282), .B(n1310), .C(n1659), .Y(n955) );
  NAND2X1 U1494 ( .A(\mem<12><1> ), .B(n61), .Y(n1660) );
  OAI21X1 U1495 ( .A(n1282), .B(n1312), .C(n1660), .Y(n956) );
  NAND2X1 U1496 ( .A(\mem<12><2> ), .B(n61), .Y(n1661) );
  OAI21X1 U1497 ( .A(n1282), .B(n1314), .C(n1661), .Y(n957) );
  NAND2X1 U1498 ( .A(\mem<12><3> ), .B(n61), .Y(n1662) );
  OAI21X1 U1499 ( .A(n1282), .B(n1316), .C(n1662), .Y(n958) );
  NAND2X1 U1500 ( .A(\mem<12><4> ), .B(n61), .Y(n1663) );
  OAI21X1 U1501 ( .A(n1282), .B(n1318), .C(n1663), .Y(n959) );
  NAND2X1 U1502 ( .A(\mem<12><5> ), .B(n61), .Y(n1664) );
  OAI21X1 U1503 ( .A(n1282), .B(n1320), .C(n1664), .Y(n960) );
  NAND2X1 U1504 ( .A(\mem<12><6> ), .B(n61), .Y(n1665) );
  OAI21X1 U1505 ( .A(n1282), .B(n1322), .C(n1665), .Y(n961) );
  NAND2X1 U1506 ( .A(\mem<12><7> ), .B(n61), .Y(n1666) );
  OAI21X1 U1507 ( .A(n1282), .B(n1239), .C(n1666), .Y(n962) );
  NAND2X1 U1508 ( .A(\mem<12><8> ), .B(n61), .Y(n1667) );
  OAI21X1 U1509 ( .A(n1283), .B(n1325), .C(n1667), .Y(n963) );
  NAND2X1 U1510 ( .A(\mem<12><9> ), .B(n61), .Y(n1668) );
  OAI21X1 U1511 ( .A(n1283), .B(n1327), .C(n1668), .Y(n964) );
  NAND2X1 U1512 ( .A(\mem<12><10> ), .B(n61), .Y(n1669) );
  OAI21X1 U1513 ( .A(n1283), .B(n1329), .C(n1669), .Y(n965) );
  NAND2X1 U1514 ( .A(\mem<12><11> ), .B(n61), .Y(n1670) );
  OAI21X1 U1515 ( .A(n1283), .B(n1331), .C(n1670), .Y(n966) );
  NAND2X1 U1516 ( .A(\mem<12><12> ), .B(n61), .Y(n1671) );
  OAI21X1 U1517 ( .A(n1283), .B(n1333), .C(n1671), .Y(n967) );
  NAND2X1 U1518 ( .A(\mem<12><13> ), .B(n61), .Y(n1672) );
  OAI21X1 U1519 ( .A(n1283), .B(n1335), .C(n1672), .Y(n968) );
  NAND2X1 U1520 ( .A(\mem<12><14> ), .B(n61), .Y(n1673) );
  OAI21X1 U1521 ( .A(n1283), .B(n1225), .C(n1673), .Y(n969) );
  NAND2X1 U1522 ( .A(\mem<12><15> ), .B(n61), .Y(n1674) );
  OAI21X1 U1523 ( .A(n1283), .B(n1338), .C(n1674), .Y(n970) );
  NAND2X1 U1524 ( .A(\mem<11><0> ), .B(n23), .Y(n1675) );
  OAI21X1 U1525 ( .A(n1284), .B(n1311), .C(n1675), .Y(n971) );
  NAND2X1 U1526 ( .A(\mem<11><1> ), .B(n23), .Y(n1676) );
  OAI21X1 U1527 ( .A(n1284), .B(n1312), .C(n1676), .Y(n972) );
  NAND2X1 U1528 ( .A(\mem<11><2> ), .B(n23), .Y(n1677) );
  OAI21X1 U1529 ( .A(n1284), .B(n1314), .C(n1677), .Y(n973) );
  NAND2X1 U1530 ( .A(\mem<11><3> ), .B(n23), .Y(n1678) );
  OAI21X1 U1531 ( .A(n1284), .B(n1316), .C(n1678), .Y(n974) );
  NAND2X1 U1532 ( .A(\mem<11><4> ), .B(n23), .Y(n1679) );
  OAI21X1 U1533 ( .A(n1284), .B(n1318), .C(n1679), .Y(n975) );
  NAND2X1 U1534 ( .A(\mem<11><5> ), .B(n23), .Y(n1680) );
  OAI21X1 U1535 ( .A(n1284), .B(n1320), .C(n1680), .Y(n976) );
  NAND2X1 U1536 ( .A(\mem<11><6> ), .B(n23), .Y(n1681) );
  OAI21X1 U1537 ( .A(n1284), .B(n1322), .C(n1681), .Y(n977) );
  NAND2X1 U1538 ( .A(\mem<11><7> ), .B(n23), .Y(n1682) );
  OAI21X1 U1539 ( .A(n1284), .B(n1241), .C(n1682), .Y(n978) );
  NAND2X1 U1540 ( .A(\mem<11><8> ), .B(n23), .Y(n1683) );
  OAI21X1 U1541 ( .A(n1285), .B(n1324), .C(n1683), .Y(n979) );
  NAND2X1 U1542 ( .A(\mem<11><9> ), .B(n23), .Y(n1684) );
  OAI21X1 U1543 ( .A(n1285), .B(n1326), .C(n1684), .Y(n980) );
  NAND2X1 U1544 ( .A(\mem<11><10> ), .B(n23), .Y(n1685) );
  OAI21X1 U1545 ( .A(n1285), .B(n1328), .C(n1685), .Y(n981) );
  NAND2X1 U1546 ( .A(\mem<11><11> ), .B(n23), .Y(n1686) );
  OAI21X1 U1547 ( .A(n1285), .B(n1330), .C(n1686), .Y(n982) );
  NAND2X1 U1548 ( .A(\mem<11><12> ), .B(n23), .Y(n1687) );
  OAI21X1 U1549 ( .A(n1285), .B(n1332), .C(n1687), .Y(n983) );
  NAND2X1 U1550 ( .A(\mem<11><13> ), .B(n23), .Y(n1688) );
  OAI21X1 U1551 ( .A(n1285), .B(n1334), .C(n1688), .Y(n984) );
  NAND2X1 U1552 ( .A(\mem<11><14> ), .B(n23), .Y(n1689) );
  OAI21X1 U1553 ( .A(n1285), .B(n1225), .C(n1689), .Y(n985) );
  NAND2X1 U1554 ( .A(\mem<11><15> ), .B(n23), .Y(n1690) );
  OAI21X1 U1555 ( .A(n1285), .B(n1337), .C(n1690), .Y(n986) );
  NAND2X1 U1556 ( .A(\mem<10><0> ), .B(n63), .Y(n1691) );
  OAI21X1 U1557 ( .A(n1286), .B(n1311), .C(n1691), .Y(n987) );
  NAND2X1 U1558 ( .A(\mem<10><1> ), .B(n63), .Y(n1692) );
  OAI21X1 U1559 ( .A(n1286), .B(n1312), .C(n1692), .Y(n988) );
  NAND2X1 U1560 ( .A(\mem<10><2> ), .B(n63), .Y(n1693) );
  OAI21X1 U1561 ( .A(n1286), .B(n1314), .C(n1693), .Y(n989) );
  NAND2X1 U1562 ( .A(\mem<10><3> ), .B(n63), .Y(n1694) );
  OAI21X1 U1563 ( .A(n1286), .B(n1316), .C(n1694), .Y(n990) );
  NAND2X1 U1564 ( .A(\mem<10><4> ), .B(n63), .Y(n1695) );
  OAI21X1 U1565 ( .A(n1286), .B(n1318), .C(n1695), .Y(n991) );
  NAND2X1 U1566 ( .A(\mem<10><5> ), .B(n63), .Y(n1696) );
  OAI21X1 U1567 ( .A(n1286), .B(n1320), .C(n1696), .Y(n992) );
  NAND2X1 U1568 ( .A(\mem<10><6> ), .B(n63), .Y(n1697) );
  OAI21X1 U1569 ( .A(n1286), .B(n1322), .C(n1697), .Y(n993) );
  NAND2X1 U1570 ( .A(\mem<10><7> ), .B(n63), .Y(n1698) );
  OAI21X1 U1571 ( .A(n1286), .B(n1244), .C(n1698), .Y(n994) );
  NAND2X1 U1572 ( .A(\mem<10><8> ), .B(n63), .Y(n1699) );
  OAI21X1 U1573 ( .A(n1287), .B(n1324), .C(n1699), .Y(n995) );
  NAND2X1 U1574 ( .A(\mem<10><9> ), .B(n63), .Y(n1700) );
  OAI21X1 U1575 ( .A(n1287), .B(n1326), .C(n1700), .Y(n996) );
  NAND2X1 U1576 ( .A(\mem<10><10> ), .B(n63), .Y(n1701) );
  OAI21X1 U1577 ( .A(n1287), .B(n1328), .C(n1701), .Y(n997) );
  NAND2X1 U1578 ( .A(\mem<10><11> ), .B(n63), .Y(n1702) );
  OAI21X1 U1579 ( .A(n1287), .B(n1330), .C(n1702), .Y(n998) );
  NAND2X1 U1580 ( .A(\mem<10><12> ), .B(n63), .Y(n1703) );
  OAI21X1 U1581 ( .A(n1287), .B(n1332), .C(n1703), .Y(n999) );
  NAND2X1 U1582 ( .A(\mem<10><13> ), .B(n63), .Y(n1704) );
  OAI21X1 U1583 ( .A(n1287), .B(n1334), .C(n1704), .Y(n1000) );
  NAND2X1 U1584 ( .A(\mem<10><14> ), .B(n63), .Y(n1705) );
  OAI21X1 U1585 ( .A(n1287), .B(n1231), .C(n1705), .Y(n1001) );
  NAND2X1 U1586 ( .A(\mem<10><15> ), .B(n63), .Y(n1706) );
  OAI21X1 U1587 ( .A(n1287), .B(n1337), .C(n1706), .Y(n1002) );
  NAND2X1 U1588 ( .A(\mem<9><0> ), .B(n25), .Y(n1707) );
  OAI21X1 U1589 ( .A(n1288), .B(n1311), .C(n1707), .Y(n1003) );
  NAND2X1 U1590 ( .A(\mem<9><1> ), .B(n25), .Y(n1708) );
  OAI21X1 U1591 ( .A(n1288), .B(n1312), .C(n1708), .Y(n1004) );
  NAND2X1 U1592 ( .A(\mem<9><2> ), .B(n25), .Y(n1709) );
  OAI21X1 U1593 ( .A(n1288), .B(n1314), .C(n1709), .Y(n1005) );
  NAND2X1 U1594 ( .A(\mem<9><3> ), .B(n25), .Y(n1710) );
  OAI21X1 U1595 ( .A(n1288), .B(n1316), .C(n1710), .Y(n1006) );
  NAND2X1 U1596 ( .A(\mem<9><4> ), .B(n25), .Y(n1711) );
  OAI21X1 U1597 ( .A(n1288), .B(n1318), .C(n1711), .Y(n1007) );
  NAND2X1 U1598 ( .A(\mem<9><5> ), .B(n25), .Y(n1712) );
  OAI21X1 U1599 ( .A(n1288), .B(n1320), .C(n1712), .Y(n1008) );
  NAND2X1 U1600 ( .A(\mem<9><6> ), .B(n25), .Y(n1713) );
  OAI21X1 U1601 ( .A(n1288), .B(n1322), .C(n1713), .Y(n1009) );
  NAND2X1 U1602 ( .A(\mem<9><7> ), .B(n25), .Y(n1714) );
  OAI21X1 U1603 ( .A(n1288), .B(n1240), .C(n1714), .Y(n1010) );
  NAND2X1 U1604 ( .A(\mem<9><8> ), .B(n25), .Y(n1715) );
  OAI21X1 U1605 ( .A(n1289), .B(n1324), .C(n1715), .Y(n1011) );
  NAND2X1 U1606 ( .A(\mem<9><9> ), .B(n25), .Y(n1716) );
  OAI21X1 U1607 ( .A(n1289), .B(n1326), .C(n1716), .Y(n1012) );
  NAND2X1 U1608 ( .A(\mem<9><10> ), .B(n25), .Y(n1717) );
  OAI21X1 U1609 ( .A(n1289), .B(n1328), .C(n1717), .Y(n1013) );
  NAND2X1 U1610 ( .A(\mem<9><11> ), .B(n25), .Y(n1718) );
  OAI21X1 U1611 ( .A(n1289), .B(n1330), .C(n1718), .Y(n1014) );
  NAND2X1 U1612 ( .A(\mem<9><12> ), .B(n25), .Y(n1719) );
  OAI21X1 U1613 ( .A(n1289), .B(n1332), .C(n1719), .Y(n1015) );
  NAND2X1 U1614 ( .A(\mem<9><13> ), .B(n25), .Y(n1720) );
  OAI21X1 U1615 ( .A(n1289), .B(n1334), .C(n1720), .Y(n1016) );
  NAND2X1 U1616 ( .A(\mem<9><14> ), .B(n25), .Y(n1721) );
  OAI21X1 U1617 ( .A(n1289), .B(n1232), .C(n1721), .Y(n1017) );
  NAND2X1 U1618 ( .A(\mem<9><15> ), .B(n25), .Y(n1722) );
  OAI21X1 U1619 ( .A(n1289), .B(n1337), .C(n1722), .Y(n1018) );
  NAND2X1 U1620 ( .A(\mem<8><0> ), .B(n65), .Y(n1724) );
  OAI21X1 U1621 ( .A(n1290), .B(n1311), .C(n1724), .Y(n1019) );
  NAND2X1 U1622 ( .A(\mem<8><1> ), .B(n65), .Y(n1725) );
  OAI21X1 U1623 ( .A(n1290), .B(n1312), .C(n1725), .Y(n1020) );
  NAND2X1 U1624 ( .A(\mem<8><2> ), .B(n65), .Y(n1726) );
  OAI21X1 U1625 ( .A(n1290), .B(n1314), .C(n1726), .Y(n1021) );
  NAND2X1 U1626 ( .A(\mem<8><3> ), .B(n65), .Y(n1727) );
  OAI21X1 U1627 ( .A(n1290), .B(n1316), .C(n1727), .Y(n1022) );
  NAND2X1 U1628 ( .A(\mem<8><4> ), .B(n65), .Y(n1728) );
  OAI21X1 U1629 ( .A(n1290), .B(n1318), .C(n1728), .Y(n1023) );
  NAND2X1 U1630 ( .A(\mem<8><5> ), .B(n65), .Y(n1729) );
  OAI21X1 U1631 ( .A(n1290), .B(n1320), .C(n1729), .Y(n1024) );
  NAND2X1 U1632 ( .A(\mem<8><6> ), .B(n65), .Y(n1730) );
  OAI21X1 U1633 ( .A(n1290), .B(n1322), .C(n1730), .Y(n1025) );
  NAND2X1 U1634 ( .A(\mem<8><7> ), .B(n65), .Y(n1731) );
  OAI21X1 U1635 ( .A(n1290), .B(n1238), .C(n1731), .Y(n1026) );
  NAND2X1 U1636 ( .A(\mem<8><8> ), .B(n65), .Y(n1732) );
  OAI21X1 U1637 ( .A(n1290), .B(n1324), .C(n1732), .Y(n1027) );
  NAND2X1 U1638 ( .A(\mem<8><9> ), .B(n65), .Y(n1733) );
  OAI21X1 U1639 ( .A(n1290), .B(n1326), .C(n1733), .Y(n1028) );
  NAND2X1 U1640 ( .A(\mem<8><10> ), .B(n65), .Y(n1734) );
  OAI21X1 U1641 ( .A(n1290), .B(n1328), .C(n1734), .Y(n1029) );
  NAND2X1 U1642 ( .A(\mem<8><11> ), .B(n65), .Y(n1735) );
  OAI21X1 U1643 ( .A(n1290), .B(n1330), .C(n1735), .Y(n1030) );
  NAND2X1 U1644 ( .A(\mem<8><12> ), .B(n65), .Y(n1736) );
  OAI21X1 U1645 ( .A(n1290), .B(n1332), .C(n1736), .Y(n1031) );
  NAND2X1 U1646 ( .A(\mem<8><13> ), .B(n65), .Y(n1737) );
  OAI21X1 U1647 ( .A(n1290), .B(n1334), .C(n1737), .Y(n1032) );
  NAND2X1 U1648 ( .A(\mem<8><14> ), .B(n65), .Y(n1738) );
  OAI21X1 U1649 ( .A(n1290), .B(n1237), .C(n1738), .Y(n1033) );
  NAND2X1 U1650 ( .A(\mem<8><15> ), .B(n65), .Y(n1739) );
  OAI21X1 U1651 ( .A(n1290), .B(n1337), .C(n1739), .Y(n1034) );
  NAND3X1 U1652 ( .A(n1346), .B(n214), .C(n1348), .Y(n1740) );
  NAND2X1 U1653 ( .A(\mem<7><0> ), .B(n67), .Y(n1741) );
  OAI21X1 U1654 ( .A(n1291), .B(n1311), .C(n1741), .Y(n1035) );
  NAND2X1 U1655 ( .A(\mem<7><1> ), .B(n67), .Y(n1742) );
  OAI21X1 U1656 ( .A(n1291), .B(n1312), .C(n1742), .Y(n1036) );
  NAND2X1 U1657 ( .A(\mem<7><2> ), .B(n67), .Y(n1743) );
  OAI21X1 U1658 ( .A(n1291), .B(n1314), .C(n1743), .Y(n1037) );
  NAND2X1 U1659 ( .A(\mem<7><3> ), .B(n67), .Y(n1744) );
  OAI21X1 U1660 ( .A(n1291), .B(n1316), .C(n1744), .Y(n1038) );
  NAND2X1 U1661 ( .A(\mem<7><4> ), .B(n67), .Y(n1745) );
  OAI21X1 U1662 ( .A(n1291), .B(n1318), .C(n1745), .Y(n1039) );
  NAND2X1 U1663 ( .A(\mem<7><5> ), .B(n67), .Y(n1746) );
  OAI21X1 U1664 ( .A(n1291), .B(n1320), .C(n1746), .Y(n1040) );
  NAND2X1 U1665 ( .A(\mem<7><6> ), .B(n67), .Y(n1747) );
  OAI21X1 U1666 ( .A(n1291), .B(n1322), .C(n1747), .Y(n1041) );
  NAND2X1 U1667 ( .A(\mem<7><7> ), .B(n67), .Y(n1748) );
  OAI21X1 U1668 ( .A(n1291), .B(n1241), .C(n1748), .Y(n1042) );
  NAND2X1 U1669 ( .A(\mem<7><8> ), .B(n67), .Y(n1749) );
  OAI21X1 U1670 ( .A(n1292), .B(n1324), .C(n1749), .Y(n1043) );
  NAND2X1 U1671 ( .A(\mem<7><9> ), .B(n67), .Y(n1750) );
  OAI21X1 U1672 ( .A(n1292), .B(n1326), .C(n1750), .Y(n1044) );
  NAND2X1 U1673 ( .A(\mem<7><10> ), .B(n67), .Y(n1751) );
  OAI21X1 U1674 ( .A(n1292), .B(n1328), .C(n1751), .Y(n1045) );
  NAND2X1 U1675 ( .A(\mem<7><11> ), .B(n67), .Y(n1752) );
  OAI21X1 U1676 ( .A(n1292), .B(n1330), .C(n1752), .Y(n1046) );
  NAND2X1 U1677 ( .A(\mem<7><12> ), .B(n67), .Y(n1753) );
  OAI21X1 U1678 ( .A(n1292), .B(n1332), .C(n1753), .Y(n1047) );
  NAND2X1 U1679 ( .A(\mem<7><13> ), .B(n67), .Y(n1754) );
  OAI21X1 U1680 ( .A(n1292), .B(n1334), .C(n1754), .Y(n1048) );
  NAND2X1 U1681 ( .A(\mem<7><14> ), .B(n67), .Y(n1755) );
  OAI21X1 U1682 ( .A(n1292), .B(n1227), .C(n1755), .Y(n1049) );
  NAND2X1 U1683 ( .A(\mem<7><15> ), .B(n67), .Y(n1756) );
  OAI21X1 U1684 ( .A(n1292), .B(n1337), .C(n1756), .Y(n1050) );
  NAND2X1 U1685 ( .A(\mem<6><0> ), .B(n13), .Y(n1757) );
  OAI21X1 U1686 ( .A(n1293), .B(n1311), .C(n1757), .Y(n1051) );
  NAND2X1 U1687 ( .A(\mem<6><1> ), .B(n13), .Y(n1758) );
  OAI21X1 U1688 ( .A(n1293), .B(n1312), .C(n1758), .Y(n1052) );
  NAND2X1 U1689 ( .A(\mem<6><2> ), .B(n13), .Y(n1759) );
  OAI21X1 U1690 ( .A(n1293), .B(n1314), .C(n1759), .Y(n1053) );
  NAND2X1 U1691 ( .A(\mem<6><3> ), .B(n13), .Y(n1760) );
  OAI21X1 U1692 ( .A(n1293), .B(n1316), .C(n1760), .Y(n1054) );
  NAND2X1 U1693 ( .A(\mem<6><4> ), .B(n13), .Y(n1761) );
  OAI21X1 U1694 ( .A(n1293), .B(n1318), .C(n1761), .Y(n1055) );
  NAND2X1 U1695 ( .A(\mem<6><5> ), .B(n13), .Y(n1762) );
  OAI21X1 U1696 ( .A(n1293), .B(n1320), .C(n1762), .Y(n1056) );
  NAND2X1 U1697 ( .A(\mem<6><6> ), .B(n13), .Y(n1763) );
  OAI21X1 U1698 ( .A(n1293), .B(n1322), .C(n1763), .Y(n1057) );
  NAND2X1 U1699 ( .A(\mem<6><7> ), .B(n13), .Y(n1764) );
  OAI21X1 U1700 ( .A(n1293), .B(n1242), .C(n1764), .Y(n1058) );
  NAND2X1 U1701 ( .A(\mem<6><8> ), .B(n13), .Y(n1765) );
  OAI21X1 U1702 ( .A(n1294), .B(n1324), .C(n1765), .Y(n1059) );
  NAND2X1 U1703 ( .A(\mem<6><9> ), .B(n13), .Y(n1766) );
  OAI21X1 U1704 ( .A(n1294), .B(n1326), .C(n1766), .Y(n1060) );
  NAND2X1 U1705 ( .A(\mem<6><10> ), .B(n13), .Y(n1767) );
  OAI21X1 U1706 ( .A(n1294), .B(n1328), .C(n1767), .Y(n1061) );
  NAND2X1 U1707 ( .A(\mem<6><11> ), .B(n13), .Y(n1768) );
  OAI21X1 U1708 ( .A(n1294), .B(n1330), .C(n1768), .Y(n1062) );
  NAND2X1 U1709 ( .A(\mem<6><12> ), .B(n13), .Y(n1769) );
  OAI21X1 U1710 ( .A(n1294), .B(n1332), .C(n1769), .Y(n1063) );
  NAND2X1 U1711 ( .A(\mem<6><13> ), .B(n13), .Y(n1770) );
  OAI21X1 U1712 ( .A(n1294), .B(n1334), .C(n1770), .Y(n1064) );
  NAND2X1 U1713 ( .A(\mem<6><14> ), .B(n13), .Y(n1771) );
  OAI21X1 U1714 ( .A(n1294), .B(n1233), .C(n1771), .Y(n1065) );
  NAND2X1 U1715 ( .A(\mem<6><15> ), .B(n13), .Y(n1772) );
  OAI21X1 U1716 ( .A(n1294), .B(n1337), .C(n1772), .Y(n1066) );
  NAND2X1 U1717 ( .A(\mem<5><0> ), .B(n15), .Y(n1774) );
  OAI21X1 U1718 ( .A(n1295), .B(n1311), .C(n1774), .Y(n1067) );
  NAND2X1 U1719 ( .A(\mem<5><1> ), .B(n15), .Y(n1775) );
  OAI21X1 U1720 ( .A(n1295), .B(n1312), .C(n1775), .Y(n1068) );
  NAND2X1 U1721 ( .A(\mem<5><2> ), .B(n15), .Y(n1776) );
  OAI21X1 U1722 ( .A(n1295), .B(n1314), .C(n1776), .Y(n1069) );
  NAND2X1 U1723 ( .A(\mem<5><3> ), .B(n15), .Y(n1777) );
  OAI21X1 U1724 ( .A(n1295), .B(n1316), .C(n1777), .Y(n1070) );
  NAND2X1 U1725 ( .A(\mem<5><4> ), .B(n15), .Y(n1778) );
  OAI21X1 U1726 ( .A(n1295), .B(n1318), .C(n1778), .Y(n1071) );
  NAND2X1 U1727 ( .A(\mem<5><5> ), .B(n15), .Y(n1779) );
  OAI21X1 U1728 ( .A(n1295), .B(n1320), .C(n1779), .Y(n1072) );
  NAND2X1 U1729 ( .A(\mem<5><6> ), .B(n15), .Y(n1780) );
  OAI21X1 U1730 ( .A(n1295), .B(n1322), .C(n1780), .Y(n1073) );
  NAND2X1 U1731 ( .A(\mem<5><7> ), .B(n15), .Y(n1781) );
  OAI21X1 U1732 ( .A(n1295), .B(n1242), .C(n1781), .Y(n1074) );
  NAND2X1 U1733 ( .A(\mem<5><8> ), .B(n15), .Y(n1782) );
  OAI21X1 U1734 ( .A(n1296), .B(n1324), .C(n1782), .Y(n1075) );
  NAND2X1 U1735 ( .A(\mem<5><9> ), .B(n15), .Y(n1783) );
  OAI21X1 U1736 ( .A(n1296), .B(n1326), .C(n1783), .Y(n1076) );
  NAND2X1 U1737 ( .A(\mem<5><10> ), .B(n15), .Y(n1784) );
  OAI21X1 U1738 ( .A(n1296), .B(n1328), .C(n1784), .Y(n1077) );
  NAND2X1 U1739 ( .A(\mem<5><11> ), .B(n15), .Y(n1785) );
  OAI21X1 U1740 ( .A(n1296), .B(n1330), .C(n1785), .Y(n1078) );
  NAND2X1 U1741 ( .A(\mem<5><12> ), .B(n15), .Y(n1786) );
  OAI21X1 U1742 ( .A(n1296), .B(n1332), .C(n1786), .Y(n1079) );
  NAND2X1 U1743 ( .A(\mem<5><13> ), .B(n15), .Y(n1787) );
  OAI21X1 U1744 ( .A(n1296), .B(n1334), .C(n1787), .Y(n1080) );
  NAND2X1 U1745 ( .A(\mem<5><14> ), .B(n15), .Y(n1788) );
  OAI21X1 U1746 ( .A(n1296), .B(n1234), .C(n1788), .Y(n1081) );
  NAND2X1 U1747 ( .A(\mem<5><15> ), .B(n15), .Y(n1789) );
  OAI21X1 U1748 ( .A(n1296), .B(n1337), .C(n1789), .Y(n1082) );
  NAND2X1 U1749 ( .A(\mem<4><0> ), .B(n17), .Y(n1791) );
  OAI21X1 U1750 ( .A(n1297), .B(n1311), .C(n1791), .Y(n1083) );
  NAND2X1 U1751 ( .A(\mem<4><1> ), .B(n17), .Y(n1792) );
  OAI21X1 U1752 ( .A(n1297), .B(n1312), .C(n1792), .Y(n1084) );
  NAND2X1 U1753 ( .A(\mem<4><2> ), .B(n17), .Y(n1793) );
  OAI21X1 U1754 ( .A(n1297), .B(n1314), .C(n1793), .Y(n1085) );
  NAND2X1 U1755 ( .A(\mem<4><3> ), .B(n17), .Y(n1794) );
  OAI21X1 U1756 ( .A(n1297), .B(n1316), .C(n1794), .Y(n1086) );
  NAND2X1 U1757 ( .A(\mem<4><4> ), .B(n17), .Y(n1795) );
  OAI21X1 U1758 ( .A(n1297), .B(n1318), .C(n1795), .Y(n1087) );
  NAND2X1 U1759 ( .A(\mem<4><5> ), .B(n17), .Y(n1796) );
  OAI21X1 U1760 ( .A(n1297), .B(n1320), .C(n1796), .Y(n1088) );
  NAND2X1 U1761 ( .A(\mem<4><6> ), .B(n17), .Y(n1797) );
  OAI21X1 U1762 ( .A(n1297), .B(n1322), .C(n1797), .Y(n1089) );
  NAND2X1 U1763 ( .A(\mem<4><7> ), .B(n17), .Y(n1798) );
  OAI21X1 U1764 ( .A(n1297), .B(n1243), .C(n1798), .Y(n1090) );
  NAND2X1 U1765 ( .A(\mem<4><8> ), .B(n17), .Y(n1799) );
  OAI21X1 U1766 ( .A(n1298), .B(n1324), .C(n1799), .Y(n1091) );
  NAND2X1 U1767 ( .A(\mem<4><9> ), .B(n17), .Y(n1800) );
  OAI21X1 U1768 ( .A(n1298), .B(n1326), .C(n1800), .Y(n1092) );
  NAND2X1 U1769 ( .A(\mem<4><10> ), .B(n17), .Y(n1801) );
  OAI21X1 U1770 ( .A(n1298), .B(n1328), .C(n1801), .Y(n1093) );
  NAND2X1 U1771 ( .A(\mem<4><11> ), .B(n17), .Y(n1802) );
  OAI21X1 U1772 ( .A(n1298), .B(n1330), .C(n1802), .Y(n1094) );
  NAND2X1 U1773 ( .A(\mem<4><12> ), .B(n17), .Y(n1803) );
  OAI21X1 U1774 ( .A(n1298), .B(n1332), .C(n1803), .Y(n1095) );
  NAND2X1 U1775 ( .A(\mem<4><13> ), .B(n17), .Y(n1804) );
  OAI21X1 U1776 ( .A(n1298), .B(n1334), .C(n1804), .Y(n1096) );
  NAND2X1 U1777 ( .A(\mem<4><14> ), .B(n17), .Y(n1805) );
  OAI21X1 U1778 ( .A(n1298), .B(n1235), .C(n1805), .Y(n1097) );
  NAND2X1 U1779 ( .A(\mem<4><15> ), .B(n17), .Y(n1806) );
  OAI21X1 U1780 ( .A(n1298), .B(n1337), .C(n1806), .Y(n1098) );
  NAND2X1 U1781 ( .A(\mem<3><0> ), .B(n98), .Y(n1808) );
  OAI21X1 U1782 ( .A(n1299), .B(n1311), .C(n1808), .Y(n1099) );
  NAND2X1 U1783 ( .A(\mem<3><1> ), .B(n98), .Y(n1809) );
  OAI21X1 U1784 ( .A(n1299), .B(n1312), .C(n1809), .Y(n1100) );
  NAND2X1 U1785 ( .A(\mem<3><2> ), .B(n98), .Y(n1810) );
  OAI21X1 U1786 ( .A(n1299), .B(n1314), .C(n1810), .Y(n1101) );
  NAND2X1 U1787 ( .A(\mem<3><3> ), .B(n98), .Y(n1811) );
  OAI21X1 U1788 ( .A(n1299), .B(n1316), .C(n1811), .Y(n1102) );
  NAND2X1 U1789 ( .A(\mem<3><4> ), .B(n98), .Y(n1812) );
  OAI21X1 U1790 ( .A(n1299), .B(n1318), .C(n1812), .Y(n1103) );
  NAND2X1 U1791 ( .A(\mem<3><5> ), .B(n98), .Y(n1813) );
  OAI21X1 U1792 ( .A(n1299), .B(n1320), .C(n1813), .Y(n1104) );
  NAND2X1 U1793 ( .A(\mem<3><6> ), .B(n98), .Y(n1814) );
  OAI21X1 U1794 ( .A(n1299), .B(n1322), .C(n1814), .Y(n1105) );
  NAND2X1 U1795 ( .A(\mem<3><7> ), .B(n98), .Y(n1815) );
  OAI21X1 U1796 ( .A(n1299), .B(n1244), .C(n1815), .Y(n1106) );
  NAND2X1 U1797 ( .A(\mem<3><8> ), .B(n98), .Y(n1816) );
  OAI21X1 U1798 ( .A(n1300), .B(n1324), .C(n1816), .Y(n1107) );
  NAND2X1 U1799 ( .A(\mem<3><9> ), .B(n98), .Y(n1817) );
  OAI21X1 U1800 ( .A(n1300), .B(n1326), .C(n1817), .Y(n1108) );
  NAND2X1 U1801 ( .A(\mem<3><10> ), .B(n98), .Y(n1818) );
  OAI21X1 U1802 ( .A(n1300), .B(n1328), .C(n1818), .Y(n1109) );
  NAND2X1 U1803 ( .A(\mem<3><11> ), .B(n98), .Y(n1819) );
  OAI21X1 U1804 ( .A(n1300), .B(n1330), .C(n1819), .Y(n1110) );
  NAND2X1 U1805 ( .A(\mem<3><12> ), .B(n98), .Y(n1820) );
  OAI21X1 U1806 ( .A(n1300), .B(n1332), .C(n1820), .Y(n1111) );
  NAND2X1 U1807 ( .A(\mem<3><13> ), .B(n98), .Y(n1821) );
  OAI21X1 U1808 ( .A(n1300), .B(n1334), .C(n1821), .Y(n1112) );
  NAND2X1 U1809 ( .A(\mem<3><14> ), .B(n98), .Y(n1822) );
  OAI21X1 U1810 ( .A(n1300), .B(n1224), .C(n1822), .Y(n1113) );
  NAND2X1 U1811 ( .A(\mem<3><15> ), .B(n98), .Y(n1823) );
  OAI21X1 U1812 ( .A(n1300), .B(n1337), .C(n1823), .Y(n1114) );
  NAND2X1 U1813 ( .A(\mem<2><0> ), .B(n99), .Y(n1825) );
  OAI21X1 U1814 ( .A(n1301), .B(n1311), .C(n1825), .Y(n1115) );
  NAND2X1 U1815 ( .A(\mem<2><1> ), .B(n99), .Y(n1826) );
  OAI21X1 U1816 ( .A(n1301), .B(n1312), .C(n1826), .Y(n1116) );
  NAND2X1 U1817 ( .A(\mem<2><2> ), .B(n99), .Y(n1827) );
  OAI21X1 U1818 ( .A(n1301), .B(n1314), .C(n1827), .Y(n1117) );
  NAND2X1 U1819 ( .A(\mem<2><3> ), .B(n99), .Y(n1828) );
  OAI21X1 U1820 ( .A(n1301), .B(n1316), .C(n1828), .Y(n1118) );
  NAND2X1 U1821 ( .A(\mem<2><4> ), .B(n99), .Y(n1829) );
  OAI21X1 U1822 ( .A(n1301), .B(n1318), .C(n1829), .Y(n1119) );
  NAND2X1 U1823 ( .A(\mem<2><5> ), .B(n99), .Y(n1830) );
  OAI21X1 U1824 ( .A(n1301), .B(n1320), .C(n1830), .Y(n1120) );
  NAND2X1 U1825 ( .A(\mem<2><6> ), .B(n99), .Y(n1831) );
  OAI21X1 U1826 ( .A(n1301), .B(n1322), .C(n1831), .Y(n1121) );
  NAND2X1 U1827 ( .A(\mem<2><7> ), .B(n99), .Y(n1832) );
  OAI21X1 U1828 ( .A(n1301), .B(n1241), .C(n1832), .Y(n1122) );
  NAND2X1 U1829 ( .A(\mem<2><8> ), .B(n99), .Y(n1833) );
  OAI21X1 U1830 ( .A(n1302), .B(n1324), .C(n1833), .Y(n1123) );
  NAND2X1 U1831 ( .A(\mem<2><9> ), .B(n99), .Y(n1834) );
  OAI21X1 U1832 ( .A(n1302), .B(n1326), .C(n1834), .Y(n1124) );
  NAND2X1 U1833 ( .A(\mem<2><10> ), .B(n99), .Y(n1835) );
  OAI21X1 U1834 ( .A(n1302), .B(n1328), .C(n1835), .Y(n1125) );
  NAND2X1 U1835 ( .A(\mem<2><11> ), .B(n99), .Y(n1836) );
  OAI21X1 U1836 ( .A(n1302), .B(n1330), .C(n1836), .Y(n1126) );
  NAND2X1 U1837 ( .A(\mem<2><12> ), .B(n99), .Y(n1837) );
  OAI21X1 U1838 ( .A(n1302), .B(n1332), .C(n1837), .Y(n1127) );
  NAND2X1 U1839 ( .A(\mem<2><13> ), .B(n99), .Y(n1838) );
  OAI21X1 U1840 ( .A(n1302), .B(n1334), .C(n1838), .Y(n1128) );
  NAND2X1 U1841 ( .A(\mem<2><14> ), .B(n99), .Y(n1839) );
  OAI21X1 U1842 ( .A(n1302), .B(n1221), .C(n1839), .Y(n1129) );
  NAND2X1 U1843 ( .A(\mem<2><15> ), .B(n99), .Y(n1840) );
  OAI21X1 U1844 ( .A(n1302), .B(n1337), .C(n1840), .Y(n1130) );
  NAND2X1 U1845 ( .A(\mem<1><0> ), .B(n100), .Y(n1842) );
  OAI21X1 U1846 ( .A(n1303), .B(n1311), .C(n1842), .Y(n1131) );
  NAND2X1 U1847 ( .A(\mem<1><1> ), .B(n100), .Y(n1843) );
  OAI21X1 U1848 ( .A(n1303), .B(n1312), .C(n1843), .Y(n1132) );
  NAND2X1 U1849 ( .A(\mem<1><2> ), .B(n100), .Y(n1844) );
  OAI21X1 U1850 ( .A(n1303), .B(n1314), .C(n1844), .Y(n1133) );
  NAND2X1 U1851 ( .A(\mem<1><3> ), .B(n100), .Y(n1845) );
  OAI21X1 U1852 ( .A(n1303), .B(n1316), .C(n1845), .Y(n1134) );
  NAND2X1 U1853 ( .A(\mem<1><4> ), .B(n100), .Y(n1846) );
  OAI21X1 U1854 ( .A(n1303), .B(n1318), .C(n1846), .Y(n1135) );
  NAND2X1 U1855 ( .A(\mem<1><5> ), .B(n100), .Y(n1847) );
  OAI21X1 U1856 ( .A(n1303), .B(n1320), .C(n1847), .Y(n1136) );
  NAND2X1 U1857 ( .A(\mem<1><6> ), .B(n100), .Y(n1848) );
  OAI21X1 U1858 ( .A(n1303), .B(n1322), .C(n1848), .Y(n1137) );
  NAND2X1 U1859 ( .A(\mem<1><7> ), .B(n100), .Y(n1849) );
  OAI21X1 U1860 ( .A(n1303), .B(n1240), .C(n1849), .Y(n1138) );
  NAND2X1 U1861 ( .A(\mem<1><8> ), .B(n100), .Y(n1850) );
  OAI21X1 U1862 ( .A(n1304), .B(n1324), .C(n1850), .Y(n1139) );
  NAND2X1 U1863 ( .A(\mem<1><9> ), .B(n100), .Y(n1851) );
  OAI21X1 U1864 ( .A(n1304), .B(n1326), .C(n1851), .Y(n1140) );
  NAND2X1 U1865 ( .A(\mem<1><10> ), .B(n100), .Y(n1852) );
  OAI21X1 U1866 ( .A(n1304), .B(n1328), .C(n1852), .Y(n1141) );
  NAND2X1 U1867 ( .A(\mem<1><11> ), .B(n100), .Y(n1853) );
  OAI21X1 U1868 ( .A(n1304), .B(n1330), .C(n1853), .Y(n1142) );
  NAND2X1 U1869 ( .A(\mem<1><12> ), .B(n100), .Y(n1854) );
  OAI21X1 U1870 ( .A(n1304), .B(n1332), .C(n1854), .Y(n1143) );
  NAND2X1 U1871 ( .A(\mem<1><13> ), .B(n100), .Y(n1855) );
  OAI21X1 U1872 ( .A(n1304), .B(n1334), .C(n1855), .Y(n1144) );
  NAND2X1 U1873 ( .A(\mem<1><14> ), .B(n100), .Y(n1856) );
  OAI21X1 U1874 ( .A(n1304), .B(n1222), .C(n1856), .Y(n1145) );
  NAND2X1 U1875 ( .A(\mem<1><15> ), .B(n100), .Y(n1857) );
  OAI21X1 U1876 ( .A(n1304), .B(n1337), .C(n1857), .Y(n1146) );
  NAND2X1 U1877 ( .A(\mem<0><0> ), .B(n69), .Y(n1860) );
  OAI21X1 U1878 ( .A(n1305), .B(n1311), .C(n1860), .Y(n1147) );
  NAND2X1 U1879 ( .A(\mem<0><1> ), .B(n69), .Y(n1861) );
  OAI21X1 U1880 ( .A(n1305), .B(n1312), .C(n1861), .Y(n1148) );
  NAND2X1 U1881 ( .A(\mem<0><2> ), .B(n69), .Y(n1862) );
  OAI21X1 U1882 ( .A(n1305), .B(n1314), .C(n1862), .Y(n1149) );
  NAND2X1 U1883 ( .A(\mem<0><3> ), .B(n69), .Y(n1863) );
  OAI21X1 U1884 ( .A(n1305), .B(n1316), .C(n1863), .Y(n1150) );
  NAND2X1 U1885 ( .A(\mem<0><4> ), .B(n69), .Y(n1864) );
  OAI21X1 U1886 ( .A(n1305), .B(n1318), .C(n1864), .Y(n1151) );
  NAND2X1 U1887 ( .A(\mem<0><5> ), .B(n69), .Y(n1865) );
  OAI21X1 U1888 ( .A(n1305), .B(n1320), .C(n1865), .Y(n1152) );
  NAND2X1 U1889 ( .A(\mem<0><6> ), .B(n69), .Y(n1866) );
  OAI21X1 U1890 ( .A(n1305), .B(n1322), .C(n1866), .Y(n1153) );
  NAND2X1 U1891 ( .A(\mem<0><7> ), .B(n69), .Y(n1867) );
  OAI21X1 U1892 ( .A(n1305), .B(n1238), .C(n1867), .Y(n1154) );
  NAND2X1 U1893 ( .A(\mem<0><8> ), .B(n69), .Y(n1868) );
  OAI21X1 U1894 ( .A(n1305), .B(n1324), .C(n1868), .Y(n1155) );
  NAND2X1 U1895 ( .A(\mem<0><9> ), .B(n69), .Y(n1869) );
  OAI21X1 U1896 ( .A(n1305), .B(n1326), .C(n1869), .Y(n1156) );
  NAND2X1 U1897 ( .A(\mem<0><10> ), .B(n69), .Y(n1870) );
  OAI21X1 U1898 ( .A(n1305), .B(n1328), .C(n1870), .Y(n1157) );
  NAND2X1 U1899 ( .A(\mem<0><11> ), .B(n69), .Y(n1871) );
  OAI21X1 U1900 ( .A(n1305), .B(n1330), .C(n1871), .Y(n1158) );
  NAND2X1 U1901 ( .A(\mem<0><12> ), .B(n69), .Y(n1872) );
  OAI21X1 U1902 ( .A(n1305), .B(n1332), .C(n1872), .Y(n1159) );
  NAND2X1 U1903 ( .A(\mem<0><13> ), .B(n69), .Y(n1873) );
  OAI21X1 U1904 ( .A(n1305), .B(n1334), .C(n1873), .Y(n1160) );
  NAND2X1 U1905 ( .A(\mem<0><14> ), .B(n69), .Y(n1874) );
  OAI21X1 U1906 ( .A(n1305), .B(n1227), .C(n1874), .Y(n1161) );
  NAND2X1 U1907 ( .A(\mem<0><15> ), .B(n69), .Y(n1875) );
  OAI21X1 U1908 ( .A(n1305), .B(n1337), .C(n1875), .Y(n1162) );
endmodule


module memc_Size16_6 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1853), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1854), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1855), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1856), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1857), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1858), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1859), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1860), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1861), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1862), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1863), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1864), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1865), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1866), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1867), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1868), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1869), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1870), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1871), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1872), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1873), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1874), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1875), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1876), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1877), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1878), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1879), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1880), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1881), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1882), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1883), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1884), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1885), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1886), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1887), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1888), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1889), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1890), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1891), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1892), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1893), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1894), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1895), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1896), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1897), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1898), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1899), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1900), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1901), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1902), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1903), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1904), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1905), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1906), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1907), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1908), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1909), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1910), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1911), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1912), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1913), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1914), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1915), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1916), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1917), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1918), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1919), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1920), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1921), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1922), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1923), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1924), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1925), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1926), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1927), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1928), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1929), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1930), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1931), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1932), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1933), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1934), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1935), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1936), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1937), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1938), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1939), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1940), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1941), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1942), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1943), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1944), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1945), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1946), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1947), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1948), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1949), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1950), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1951), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1952), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1953), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1954), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1955), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1956), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1957), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1958), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1959), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1960), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1961), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1962), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1963), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1964), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1965), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1966), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1967), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1968), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1969), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1970), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1971), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1972), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1973), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1974), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1975), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1976), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1977), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1978), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1979), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1980), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1981), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1982), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1983), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1984), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1985), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1986), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1987), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1988), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1989), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1990), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1991), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1992), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1993), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1994), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1995), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1996), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1997), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1998), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1999), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2000), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2001), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2002), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2003), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2004), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2005), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2006), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2007), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2008), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2009), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2010), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2011), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2012), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2013), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2014), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2015), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2016), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2017), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2018), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2019), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2020), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2021), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2022), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2023), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2024), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2025), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2026), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2027), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2028), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2029), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2030), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2031), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2032), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2033), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2034), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2035), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2036), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2037), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2038), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2039), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2040), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2041), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2042), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2043), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2044), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2045), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2046), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2047), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2048), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2049), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2050), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2051), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2052), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2053), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2054), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2055), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2056), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2057), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2058), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2059), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2060), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2061), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2062), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2063), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2064), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2065), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2066), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2067), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2068), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2069), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2070), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2071), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2072), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2073), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2074), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2075), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2076), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2077), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2078), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2079), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2080), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2081), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2082), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2083), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2084), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2085), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2086), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2087), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2088), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2089), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2090), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2091), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2092), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2093), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2094), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2095), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2096), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2097), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2098), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2099), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2100), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2101), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2102), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2103), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2104), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2105), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2106), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2107), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2108), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2109), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2110), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2111), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2112), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2113), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2114), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2115), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2116), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2117), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2118), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2119), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2120), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2121), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2122), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2123), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2124), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2125), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2126), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2127), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2128), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2129), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2130), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2131), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2132), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2133), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2134), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2135), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2136), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2137), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2138), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2139), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2140), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2141), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2142), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2143), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2144), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2145), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2146), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2147), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2148), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2149), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2150), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2151), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2152), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2153), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2154), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2155), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2156), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2157), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2158), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2159), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2160), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2161), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2162), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2163), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2164), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2165), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2166), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2167), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2168), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2169), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2170), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2171), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2172), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2173), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2174), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2175), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2176), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2177), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2178), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2179), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2180), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2181), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2182), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2183), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2184), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2185), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2186), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2187), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2188), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2189), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2190), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2191), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2192), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2193), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2194), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2195), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2196), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2197), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2198), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2199), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2200), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2201), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2202), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2203), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2204), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2205), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2206), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2207), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2208), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2209), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2210), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2211), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2212), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2213), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2214), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2215), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2216), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2217), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2218), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2219), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2220), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2221), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2222), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2223), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2224), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2225), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2226), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2227), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2228), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2229), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2230), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2231), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2232), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2233), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2234), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2235), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2236), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2237), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2238), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2239), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2240), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2241), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2242), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2243), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2244), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2245), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2246), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2247), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2248), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2249), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2250), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2251), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2252), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2253), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2254), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2255), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2256), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2257), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2258), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2259), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2260), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2261), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2262), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2263), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2264), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2265), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2266), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2267), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2268), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2269), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2270), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2271), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2272), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2273), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2274), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2275), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2276), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2277), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2278), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2279), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2280), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2281), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2282), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2283), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2284), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2285), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2286), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2287), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2288), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2289), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2290), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2291), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2292), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2293), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2294), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2295), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2296), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2297), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2298), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2299), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2300), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2301), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2302), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2303), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2304), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2305), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2306), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2307), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2308), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2309), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2310), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2311), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2312), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2313), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2314), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2315), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2316), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2317), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2318), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2319), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2320), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2321), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2322), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2323), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2324), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2325), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2326), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2327), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2328), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2329), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2330), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2331), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2332), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2333), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2334), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2335), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2336), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2337), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2338), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2339), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2340), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2341), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2342), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2343), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2344), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2345), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2346), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2347), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2348), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2349), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2350), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2351), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2352), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2353), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2354), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2355), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2356), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2357), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2358), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2359), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2360), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2361), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2362), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2363), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2364), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2365) );
  INVX4 U2 ( .A(n76), .Y(n77) );
  INVX4 U3 ( .A(n74), .Y(n75) );
  INVX4 U4 ( .A(n72), .Y(n73) );
  INVX4 U5 ( .A(n70), .Y(n71) );
  INVX4 U6 ( .A(n68), .Y(n69) );
  INVX4 U7 ( .A(n66), .Y(n67) );
  INVX4 U8 ( .A(n64), .Y(n65) );
  INVX4 U9 ( .A(n36), .Y(n37) );
  INVX4 U10 ( .A(n34), .Y(n35) );
  INVX4 U11 ( .A(n28), .Y(n29) );
  INVX4 U12 ( .A(n22), .Y(n23) );
  INVX4 U13 ( .A(n18), .Y(n19) );
  INVX4 U14 ( .A(n62), .Y(n63) );
  INVX4 U15 ( .A(n60), .Y(n61) );
  INVX4 U16 ( .A(n58), .Y(n59) );
  INVX4 U17 ( .A(n56), .Y(n57) );
  INVX4 U18 ( .A(n54), .Y(n55) );
  INVX4 U19 ( .A(n52), .Y(n53) );
  INVX4 U20 ( .A(n50), .Y(n51) );
  INVX4 U21 ( .A(n48), .Y(n49) );
  INVX4 U22 ( .A(n46), .Y(n47) );
  INVX4 U23 ( .A(n44), .Y(n45) );
  INVX4 U24 ( .A(n38), .Y(n39) );
  INVX4 U25 ( .A(n32), .Y(n33) );
  INVX4 U26 ( .A(n30), .Y(n31) );
  INVX4 U27 ( .A(n26), .Y(n27) );
  INVX4 U28 ( .A(n24), .Y(n25) );
  INVX4 U29 ( .A(n20), .Y(n21) );
  INVX4 U30 ( .A(n42), .Y(n43) );
  INVX4 U31 ( .A(n40), .Y(n41) );
  INVX2 U32 ( .A(n2), .Y(n3) );
  INVX1 U33 ( .A(n639), .Y(N32) );
  INVX1 U34 ( .A(n640), .Y(N31) );
  INVX1 U35 ( .A(n641), .Y(N30) );
  INVX1 U36 ( .A(n642), .Y(N29) );
  INVX1 U37 ( .A(n643), .Y(N28) );
  INVX1 U38 ( .A(n644), .Y(N27) );
  INVX1 U39 ( .A(n645), .Y(N26) );
  INVX1 U40 ( .A(n646), .Y(N25) );
  INVX1 U41 ( .A(n647), .Y(N24) );
  INVX1 U42 ( .A(n648), .Y(N23) );
  INVX1 U43 ( .A(n649), .Y(N22) );
  INVX1 U44 ( .A(n650), .Y(N21) );
  INVX1 U45 ( .A(n1163), .Y(N20) );
  INVX1 U46 ( .A(n1164), .Y(N19) );
  INVX1 U47 ( .A(n1165), .Y(N18) );
  INVX1 U48 ( .A(n1166), .Y(N17) );
  INVX1 U49 ( .A(n1217), .Y(n1219) );
  INVX1 U50 ( .A(n1219), .Y(n1194) );
  INVX1 U51 ( .A(n1219), .Y(n1193) );
  INVX1 U52 ( .A(n1219), .Y(n1192) );
  INVX1 U53 ( .A(n1218), .Y(n1191) );
  INVX2 U54 ( .A(n1218), .Y(n1190) );
  INVX2 U55 ( .A(n1194), .Y(n1196) );
  INVX1 U56 ( .A(n1194), .Y(n1195) );
  INVX1 U57 ( .A(n1188), .Y(n1177) );
  INVX2 U58 ( .A(n1193), .Y(n1198) );
  INVX1 U59 ( .A(n1188), .Y(n1178) );
  INVX1 U60 ( .A(n1321), .Y(n1174) );
  INVX1 U61 ( .A(n1188), .Y(n1179) );
  INVX2 U62 ( .A(n1192), .Y(n1201) );
  INVX2 U63 ( .A(n1192), .Y(n1202) );
  INVX1 U64 ( .A(n1176), .Y(n1180) );
  INVX1 U65 ( .A(n1321), .Y(n1173) );
  INVX1 U66 ( .A(n1176), .Y(n1181) );
  INVX2 U67 ( .A(n1176), .Y(n1182) );
  INVX1 U68 ( .A(n1321), .Y(n1172) );
  INVX1 U69 ( .A(n1175), .Y(n1183) );
  INVX1 U70 ( .A(n1175), .Y(n1184) );
  INVX2 U71 ( .A(n1175), .Y(n1185) );
  INVX2 U72 ( .A(n1176), .Y(n1186) );
  INVX2 U73 ( .A(n1175), .Y(n1187) );
  BUFX2 U74 ( .A(n103), .Y(n1220) );
  BUFX2 U75 ( .A(n105), .Y(n1222) );
  BUFX2 U76 ( .A(n107), .Y(n1224) );
  BUFX2 U77 ( .A(n109), .Y(n1226) );
  BUFX2 U78 ( .A(n111), .Y(n1228) );
  BUFX2 U79 ( .A(n113), .Y(n1230) );
  BUFX2 U80 ( .A(n115), .Y(n1232) );
  BUFX2 U81 ( .A(n117), .Y(n1235) );
  BUFX2 U82 ( .A(n119), .Y(n1237) );
  BUFX2 U83 ( .A(n121), .Y(n1239) );
  BUFX2 U84 ( .A(n123), .Y(n1241) );
  BUFX2 U85 ( .A(n125), .Y(n1243) );
  BUFX2 U86 ( .A(n127), .Y(n1245) );
  BUFX2 U87 ( .A(n129), .Y(n1247) );
  BUFX2 U88 ( .A(n131), .Y(n1250) );
  BUFX2 U89 ( .A(n133), .Y(n1252) );
  BUFX2 U90 ( .A(n135), .Y(n1254) );
  BUFX2 U91 ( .A(n137), .Y(n1256) );
  BUFX2 U92 ( .A(n139), .Y(n1258) );
  BUFX2 U93 ( .A(n141), .Y(n1260) );
  BUFX2 U94 ( .A(n143), .Y(n1262) );
  BUFX2 U95 ( .A(n145), .Y(n1265) );
  BUFX2 U96 ( .A(n147), .Y(n1267) );
  BUFX2 U97 ( .A(n149), .Y(n1269) );
  BUFX2 U98 ( .A(n151), .Y(n1271) );
  BUFX2 U99 ( .A(n153), .Y(n1273) );
  BUFX2 U100 ( .A(n155), .Y(n1275) );
  BUFX2 U101 ( .A(n157), .Y(n1277) );
  INVX2 U102 ( .A(n2), .Y(n1) );
  INVX1 U103 ( .A(n1217), .Y(n1218) );
  INVX1 U104 ( .A(n1318), .Y(n1188) );
  INVX1 U105 ( .A(n1323), .Y(n1169) );
  INVX1 U106 ( .A(n1323), .Y(n1168) );
  INVX1 U107 ( .A(N12), .Y(n1321) );
  INVX1 U108 ( .A(n1321), .Y(n1170) );
  INVX1 U109 ( .A(n1321), .Y(n1171) );
  INVX1 U110 ( .A(n1325), .Y(n1324) );
  INVX1 U111 ( .A(N14), .Y(n1325) );
  INVX1 U112 ( .A(n1316), .Y(n1217) );
  INVX2 U113 ( .A(n1316), .Y(n1189) );
  INVX1 U114 ( .A(n1323), .Y(n1322) );
  INVX1 U115 ( .A(N13), .Y(n1323) );
  INVX1 U116 ( .A(n1318), .Y(n1175) );
  INVX1 U117 ( .A(n1318), .Y(n1176) );
  INVX1 U118 ( .A(rst), .Y(n1315) );
  BUFX2 U119 ( .A(n107), .Y(n1225) );
  BUFX2 U120 ( .A(n109), .Y(n1227) );
  INVX1 U121 ( .A(n1325), .Y(n1167) );
  INVX1 U122 ( .A(n99), .Y(n1249) );
  INVX1 U123 ( .A(n101), .Y(n1279) );
  INVX1 U124 ( .A(n100), .Y(n1264) );
  INVX1 U125 ( .A(n98), .Y(n1234) );
  BUFX2 U126 ( .A(n103), .Y(n1221) );
  BUFX2 U127 ( .A(n105), .Y(n1223) );
  BUFX2 U128 ( .A(n119), .Y(n1238) );
  BUFX2 U129 ( .A(n121), .Y(n1240) );
  BUFX2 U130 ( .A(n123), .Y(n1242) );
  BUFX2 U131 ( .A(n111), .Y(n1229) );
  BUFX2 U132 ( .A(n113), .Y(n1231) );
  BUFX2 U133 ( .A(n115), .Y(n1233) );
  BUFX2 U134 ( .A(n117), .Y(n1236) );
  BUFX2 U135 ( .A(n131), .Y(n1251) );
  BUFX2 U136 ( .A(n145), .Y(n1266) );
  BUFX2 U137 ( .A(n157), .Y(n1278) );
  BUFX2 U138 ( .A(n125), .Y(n1244) );
  BUFX2 U139 ( .A(n127), .Y(n1246) );
  BUFX2 U140 ( .A(n129), .Y(n1248) );
  BUFX2 U141 ( .A(n133), .Y(n1253) );
  BUFX2 U142 ( .A(n135), .Y(n1255) );
  BUFX2 U143 ( .A(n137), .Y(n1257) );
  BUFX2 U144 ( .A(n139), .Y(n1259) );
  BUFX2 U145 ( .A(n141), .Y(n1261) );
  BUFX2 U146 ( .A(n143), .Y(n1263) );
  BUFX2 U147 ( .A(n147), .Y(n1268) );
  BUFX2 U148 ( .A(n149), .Y(n1270) );
  BUFX2 U149 ( .A(n151), .Y(n1272) );
  BUFX2 U150 ( .A(n153), .Y(n1274) );
  BUFX2 U151 ( .A(n155), .Y(n1276) );
  INVX4 U152 ( .A(n16), .Y(n83) );
  INVX4 U153 ( .A(n15), .Y(n82) );
  INVX4 U154 ( .A(n17), .Y(n1282) );
  OR2X2 U155 ( .A(write), .B(rst), .Y(n2) );
  AND2X2 U156 ( .A(\data_in<0> ), .B(n1281), .Y(n4) );
  AND2X2 U157 ( .A(\data_in<1> ), .B(n1280), .Y(n5) );
  AND2X2 U158 ( .A(\data_in<2> ), .B(n1280), .Y(n6) );
  AND2X2 U159 ( .A(\data_in<3> ), .B(n17), .Y(n7) );
  AND2X2 U160 ( .A(\data_in<4> ), .B(n1281), .Y(n8) );
  AND2X2 U161 ( .A(\data_in<5> ), .B(n1281), .Y(n9) );
  AND2X2 U162 ( .A(\data_in<6> ), .B(n1280), .Y(n10) );
  AND2X2 U163 ( .A(\data_in<7> ), .B(n17), .Y(n11) );
  AND2X2 U164 ( .A(\data_in<8> ), .B(n1281), .Y(n12) );
  AND2X2 U165 ( .A(\data_in<9> ), .B(n1281), .Y(n13) );
  AND2X2 U166 ( .A(\data_in<10> ), .B(n1280), .Y(n14) );
  AND2X2 U167 ( .A(n1280), .B(n99), .Y(n15) );
  AND2X2 U168 ( .A(n1280), .B(n101), .Y(n16) );
  AND2X2 U169 ( .A(write), .B(n1315), .Y(n17) );
  AND2X2 U170 ( .A(n1281), .B(n110), .Y(n18) );
  AND2X2 U171 ( .A(n1280), .B(n112), .Y(n20) );
  AND2X2 U172 ( .A(n1281), .B(n114), .Y(n22) );
  AND2X2 U173 ( .A(n1280), .B(n98), .Y(n24) );
  AND2X2 U174 ( .A(n1280), .B(n116), .Y(n26) );
  AND2X2 U175 ( .A(n1281), .B(n118), .Y(n28) );
  AND2X2 U176 ( .A(n1280), .B(n120), .Y(n30) );
  AND2X2 U177 ( .A(n1280), .B(n102), .Y(n32) );
  AND2X2 U178 ( .A(n1281), .B(n122), .Y(n34) );
  AND2X2 U179 ( .A(n1281), .B(n156), .Y(n36) );
  AND2X2 U180 ( .A(n1280), .B(n104), .Y(n38) );
  AND2X2 U181 ( .A(n17), .B(n106), .Y(n40) );
  AND2X2 U182 ( .A(n17), .B(n108), .Y(n42) );
  AND2X2 U183 ( .A(n1280), .B(n124), .Y(n44) );
  AND2X2 U184 ( .A(n1280), .B(n126), .Y(n46) );
  AND2X2 U185 ( .A(n1280), .B(n128), .Y(n48) );
  AND2X2 U186 ( .A(n1280), .B(n130), .Y(n50) );
  AND2X2 U187 ( .A(n1280), .B(n132), .Y(n52) );
  AND2X2 U188 ( .A(n1280), .B(n134), .Y(n54) );
  AND2X2 U189 ( .A(n1280), .B(n136), .Y(n56) );
  AND2X2 U190 ( .A(n1280), .B(n138), .Y(n58) );
  AND2X2 U191 ( .A(n1280), .B(n140), .Y(n60) );
  AND2X2 U192 ( .A(n1280), .B(n142), .Y(n62) );
  AND2X2 U193 ( .A(n1281), .B(n100), .Y(n64) );
  AND2X2 U194 ( .A(n1281), .B(n144), .Y(n66) );
  AND2X2 U195 ( .A(n1281), .B(n146), .Y(n68) );
  AND2X2 U196 ( .A(n1281), .B(n148), .Y(n70) );
  AND2X2 U197 ( .A(n1281), .B(n150), .Y(n72) );
  AND2X2 U198 ( .A(n1281), .B(n152), .Y(n74) );
  AND2X2 U199 ( .A(n1281), .B(n154), .Y(n76) );
  AND2X2 U200 ( .A(\data_in<12> ), .B(n1281), .Y(n78) );
  AND2X2 U201 ( .A(\data_in<13> ), .B(n1281), .Y(n79) );
  AND2X2 U202 ( .A(\data_in<14> ), .B(n1281), .Y(n80) );
  AND2X2 U203 ( .A(\data_in<15> ), .B(n1281), .Y(n81) );
  INVX1 U204 ( .A(n1321), .Y(n1320) );
  INVX1 U205 ( .A(n1317), .Y(n1316) );
  AND2X1 U206 ( .A(n1320), .B(n1318), .Y(n84) );
  INVX1 U207 ( .A(n1319), .Y(n1318) );
  AND2X1 U208 ( .A(n2365), .B(n1324), .Y(n85) );
  AND2X2 U209 ( .A(\data_in<11> ), .B(n1281), .Y(n86) );
  BUFX2 U210 ( .A(n1358), .Y(n87) );
  INVX1 U211 ( .A(n87), .Y(n1750) );
  BUFX2 U212 ( .A(n1375), .Y(n88) );
  INVX1 U213 ( .A(n88), .Y(n1767) );
  BUFX2 U214 ( .A(n1392), .Y(n89) );
  INVX1 U215 ( .A(n89), .Y(n1784) );
  BUFX2 U216 ( .A(n1409), .Y(n90) );
  INVX1 U217 ( .A(n90), .Y(n1801) );
  BUFX2 U218 ( .A(n1426), .Y(n91) );
  INVX1 U219 ( .A(n91), .Y(n1818) );
  BUFX2 U220 ( .A(n1587), .Y(n92) );
  INVX1 U221 ( .A(n92), .Y(n1700) );
  BUFX2 U222 ( .A(n1717), .Y(n93) );
  INVX1 U223 ( .A(n93), .Y(n1835) );
  AND2X1 U224 ( .A(n1316), .B(n84), .Y(n94) );
  AND2X1 U225 ( .A(n1322), .B(n85), .Y(n95) );
  AND2X1 U226 ( .A(n1317), .B(n84), .Y(n96) );
  AND2X1 U227 ( .A(n1323), .B(n85), .Y(n97) );
  AND2X1 U228 ( .A(n95), .B(n1836), .Y(n98) );
  AND2X1 U229 ( .A(n1836), .B(n97), .Y(n99) );
  AND2X1 U230 ( .A(n1836), .B(n1700), .Y(n100) );
  AND2X1 U231 ( .A(n1836), .B(n1835), .Y(n101) );
  AND2X1 U232 ( .A(n94), .B(n95), .Y(n102) );
  INVX1 U233 ( .A(n102), .Y(n103) );
  AND2X1 U234 ( .A(n95), .B(n96), .Y(n104) );
  INVX1 U235 ( .A(n104), .Y(n105) );
  AND2X1 U236 ( .A(n95), .B(n1750), .Y(n106) );
  INVX1 U237 ( .A(n106), .Y(n107) );
  AND2X1 U238 ( .A(n95), .B(n1767), .Y(n108) );
  INVX1 U239 ( .A(n108), .Y(n109) );
  AND2X1 U240 ( .A(n95), .B(n1784), .Y(n110) );
  INVX1 U241 ( .A(n110), .Y(n111) );
  AND2X1 U242 ( .A(n95), .B(n1801), .Y(n112) );
  INVX1 U243 ( .A(n112), .Y(n113) );
  AND2X1 U244 ( .A(n95), .B(n1818), .Y(n114) );
  INVX1 U245 ( .A(n114), .Y(n115) );
  AND2X1 U246 ( .A(n94), .B(n97), .Y(n116) );
  INVX1 U247 ( .A(n116), .Y(n117) );
  AND2X1 U248 ( .A(n96), .B(n97), .Y(n118) );
  INVX1 U249 ( .A(n118), .Y(n119) );
  AND2X1 U250 ( .A(n1750), .B(n97), .Y(n120) );
  INVX1 U251 ( .A(n120), .Y(n121) );
  AND2X1 U252 ( .A(n1767), .B(n97), .Y(n122) );
  INVX1 U253 ( .A(n122), .Y(n123) );
  AND2X1 U254 ( .A(n1784), .B(n97), .Y(n124) );
  INVX1 U255 ( .A(n124), .Y(n125) );
  AND2X1 U256 ( .A(n1801), .B(n97), .Y(n126) );
  INVX1 U257 ( .A(n126), .Y(n127) );
  AND2X1 U258 ( .A(n1818), .B(n97), .Y(n128) );
  INVX1 U259 ( .A(n128), .Y(n129) );
  AND2X1 U260 ( .A(n94), .B(n1700), .Y(n130) );
  INVX1 U261 ( .A(n130), .Y(n131) );
  AND2X1 U262 ( .A(n96), .B(n1700), .Y(n132) );
  INVX1 U263 ( .A(n132), .Y(n133) );
  AND2X1 U264 ( .A(n1750), .B(n1700), .Y(n134) );
  INVX1 U265 ( .A(n134), .Y(n135) );
  AND2X1 U266 ( .A(n1767), .B(n1700), .Y(n136) );
  INVX1 U267 ( .A(n136), .Y(n137) );
  AND2X1 U268 ( .A(n1784), .B(n1700), .Y(n138) );
  INVX1 U269 ( .A(n138), .Y(n139) );
  AND2X1 U270 ( .A(n1801), .B(n1700), .Y(n140) );
  INVX1 U271 ( .A(n140), .Y(n141) );
  AND2X1 U272 ( .A(n1818), .B(n1700), .Y(n142) );
  INVX1 U273 ( .A(n142), .Y(n143) );
  AND2X1 U274 ( .A(n94), .B(n1835), .Y(n144) );
  INVX1 U275 ( .A(n144), .Y(n145) );
  AND2X1 U276 ( .A(n96), .B(n1835), .Y(n146) );
  INVX1 U277 ( .A(n146), .Y(n147) );
  AND2X1 U278 ( .A(n1750), .B(n1835), .Y(n148) );
  INVX1 U279 ( .A(n148), .Y(n149) );
  AND2X1 U280 ( .A(n1767), .B(n1835), .Y(n150) );
  INVX1 U281 ( .A(n150), .Y(n151) );
  AND2X1 U282 ( .A(n1784), .B(n1835), .Y(n152) );
  INVX1 U283 ( .A(n152), .Y(n153) );
  AND2X1 U284 ( .A(n1801), .B(n1835), .Y(n154) );
  INVX1 U285 ( .A(n154), .Y(n155) );
  AND2X1 U286 ( .A(n1818), .B(n1835), .Y(n156) );
  INVX1 U287 ( .A(n156), .Y(n157) );
  MUX2X1 U288 ( .B(n159), .A(n160), .S(n1177), .Y(n158) );
  MUX2X1 U289 ( .B(n162), .A(n163), .S(n1177), .Y(n161) );
  MUX2X1 U290 ( .B(n165), .A(n166), .S(n1177), .Y(n164) );
  MUX2X1 U291 ( .B(n168), .A(n169), .S(n1177), .Y(n167) );
  MUX2X1 U292 ( .B(n171), .A(n172), .S(n1169), .Y(n170) );
  MUX2X1 U293 ( .B(n174), .A(n175), .S(n1177), .Y(n173) );
  MUX2X1 U294 ( .B(n177), .A(n178), .S(n1177), .Y(n176) );
  MUX2X1 U295 ( .B(n180), .A(n181), .S(n1177), .Y(n179) );
  MUX2X1 U296 ( .B(n183), .A(n184), .S(n1177), .Y(n182) );
  MUX2X1 U297 ( .B(n186), .A(n187), .S(n1169), .Y(n185) );
  MUX2X1 U298 ( .B(n189), .A(n190), .S(n1178), .Y(n188) );
  MUX2X1 U299 ( .B(n192), .A(n193), .S(n1178), .Y(n191) );
  MUX2X1 U300 ( .B(n195), .A(n196), .S(n1178), .Y(n194) );
  MUX2X1 U301 ( .B(n198), .A(n199), .S(n1178), .Y(n197) );
  MUX2X1 U302 ( .B(n201), .A(n202), .S(n1169), .Y(n200) );
  MUX2X1 U303 ( .B(n204), .A(n205), .S(n1178), .Y(n203) );
  MUX2X1 U304 ( .B(n207), .A(n208), .S(n1178), .Y(n206) );
  MUX2X1 U305 ( .B(n210), .A(n211), .S(n1178), .Y(n209) );
  MUX2X1 U306 ( .B(n213), .A(n215), .S(n1178), .Y(n212) );
  MUX2X1 U307 ( .B(n217), .A(n218), .S(n1169), .Y(n216) );
  MUX2X1 U308 ( .B(n220), .A(n221), .S(n1178), .Y(n219) );
  MUX2X1 U309 ( .B(n223), .A(n224), .S(n1178), .Y(n222) );
  MUX2X1 U310 ( .B(n226), .A(n227), .S(n1178), .Y(n225) );
  MUX2X1 U311 ( .B(n229), .A(n230), .S(n1178), .Y(n228) );
  MUX2X1 U312 ( .B(n232), .A(n233), .S(n1169), .Y(n231) );
  MUX2X1 U313 ( .B(n235), .A(n236), .S(n1179), .Y(n234) );
  MUX2X1 U314 ( .B(n238), .A(n239), .S(n1179), .Y(n237) );
  MUX2X1 U315 ( .B(n241), .A(n242), .S(n1179), .Y(n240) );
  MUX2X1 U316 ( .B(n244), .A(n245), .S(n1179), .Y(n243) );
  MUX2X1 U317 ( .B(n247), .A(n248), .S(n1169), .Y(n246) );
  MUX2X1 U318 ( .B(n250), .A(n251), .S(n1179), .Y(n249) );
  MUX2X1 U319 ( .B(n253), .A(n254), .S(n1179), .Y(n252) );
  MUX2X1 U320 ( .B(n256), .A(n257), .S(n1179), .Y(n255) );
  MUX2X1 U321 ( .B(n259), .A(n260), .S(n1179), .Y(n258) );
  MUX2X1 U322 ( .B(n262), .A(n263), .S(n1169), .Y(n261) );
  MUX2X1 U323 ( .B(n265), .A(n266), .S(n1179), .Y(n264) );
  MUX2X1 U324 ( .B(n268), .A(n269), .S(n1179), .Y(n267) );
  MUX2X1 U325 ( .B(n271), .A(n272), .S(n1179), .Y(n270) );
  MUX2X1 U326 ( .B(n274), .A(n275), .S(n1179), .Y(n273) );
  MUX2X1 U327 ( .B(n277), .A(n278), .S(n1169), .Y(n276) );
  MUX2X1 U328 ( .B(n280), .A(n281), .S(n1180), .Y(n279) );
  MUX2X1 U329 ( .B(n283), .A(n284), .S(n1180), .Y(n282) );
  MUX2X1 U330 ( .B(n286), .A(n287), .S(n1180), .Y(n285) );
  MUX2X1 U331 ( .B(n289), .A(n290), .S(n1180), .Y(n288) );
  MUX2X1 U332 ( .B(n292), .A(n293), .S(n1169), .Y(n291) );
  MUX2X1 U333 ( .B(n295), .A(n296), .S(n1180), .Y(n294) );
  MUX2X1 U334 ( .B(n298), .A(n299), .S(n1180), .Y(n297) );
  MUX2X1 U335 ( .B(n301), .A(n302), .S(n1180), .Y(n300) );
  MUX2X1 U336 ( .B(n304), .A(n305), .S(n1180), .Y(n303) );
  MUX2X1 U337 ( .B(n307), .A(n308), .S(n1169), .Y(n306) );
  MUX2X1 U338 ( .B(n310), .A(n311), .S(n1180), .Y(n309) );
  MUX2X1 U339 ( .B(n313), .A(n314), .S(n1180), .Y(n312) );
  MUX2X1 U340 ( .B(n316), .A(n317), .S(n1180), .Y(n315) );
  MUX2X1 U341 ( .B(n319), .A(n320), .S(n1180), .Y(n318) );
  MUX2X1 U342 ( .B(n322), .A(n323), .S(n1169), .Y(n321) );
  MUX2X1 U343 ( .B(n325), .A(n326), .S(n1181), .Y(n324) );
  MUX2X1 U344 ( .B(n328), .A(n329), .S(n1181), .Y(n327) );
  MUX2X1 U345 ( .B(n331), .A(n332), .S(n1181), .Y(n330) );
  MUX2X1 U346 ( .B(n334), .A(n335), .S(n1181), .Y(n333) );
  MUX2X1 U347 ( .B(n337), .A(n338), .S(n1169), .Y(n336) );
  MUX2X1 U348 ( .B(n340), .A(n341), .S(n1181), .Y(n339) );
  MUX2X1 U349 ( .B(n343), .A(n344), .S(n1181), .Y(n342) );
  MUX2X1 U350 ( .B(n346), .A(n347), .S(n1181), .Y(n345) );
  MUX2X1 U351 ( .B(n349), .A(n350), .S(n1181), .Y(n348) );
  MUX2X1 U352 ( .B(n352), .A(n353), .S(n1168), .Y(n351) );
  MUX2X1 U353 ( .B(n355), .A(n356), .S(n1181), .Y(n354) );
  MUX2X1 U354 ( .B(n358), .A(n359), .S(n1181), .Y(n357) );
  MUX2X1 U355 ( .B(n361), .A(n362), .S(n1181), .Y(n360) );
  MUX2X1 U356 ( .B(n364), .A(n365), .S(n1181), .Y(n363) );
  MUX2X1 U357 ( .B(n367), .A(n368), .S(n1168), .Y(n366) );
  MUX2X1 U358 ( .B(n370), .A(n371), .S(n1182), .Y(n369) );
  MUX2X1 U359 ( .B(n373), .A(n374), .S(n1182), .Y(n372) );
  MUX2X1 U360 ( .B(n376), .A(n377), .S(n1182), .Y(n375) );
  MUX2X1 U361 ( .B(n379), .A(n380), .S(n1182), .Y(n378) );
  MUX2X1 U362 ( .B(n382), .A(n383), .S(n1168), .Y(n381) );
  MUX2X1 U363 ( .B(n385), .A(n386), .S(n1182), .Y(n384) );
  MUX2X1 U364 ( .B(n388), .A(n389), .S(n1182), .Y(n387) );
  MUX2X1 U365 ( .B(n391), .A(n392), .S(n1182), .Y(n390) );
  MUX2X1 U366 ( .B(n394), .A(n395), .S(n1182), .Y(n393) );
  MUX2X1 U367 ( .B(n397), .A(n398), .S(n1168), .Y(n396) );
  MUX2X1 U368 ( .B(n400), .A(n401), .S(n1182), .Y(n399) );
  MUX2X1 U369 ( .B(n403), .A(n404), .S(n1182), .Y(n402) );
  MUX2X1 U370 ( .B(n406), .A(n407), .S(n1182), .Y(n405) );
  MUX2X1 U371 ( .B(n409), .A(n410), .S(n1182), .Y(n408) );
  MUX2X1 U372 ( .B(n412), .A(n413), .S(n1168), .Y(n411) );
  MUX2X1 U373 ( .B(n415), .A(n416), .S(n1183), .Y(n414) );
  MUX2X1 U374 ( .B(n418), .A(n419), .S(n1183), .Y(n417) );
  MUX2X1 U375 ( .B(n421), .A(n422), .S(n1183), .Y(n420) );
  MUX2X1 U376 ( .B(n424), .A(n425), .S(n1183), .Y(n423) );
  MUX2X1 U377 ( .B(n427), .A(n428), .S(n1168), .Y(n426) );
  MUX2X1 U378 ( .B(n430), .A(n431), .S(n1183), .Y(n429) );
  MUX2X1 U379 ( .B(n433), .A(n434), .S(n1183), .Y(n432) );
  MUX2X1 U380 ( .B(n436), .A(n437), .S(n1183), .Y(n435) );
  MUX2X1 U381 ( .B(n439), .A(n440), .S(n1183), .Y(n438) );
  MUX2X1 U382 ( .B(n442), .A(n443), .S(n1168), .Y(n441) );
  MUX2X1 U383 ( .B(n445), .A(n446), .S(n1183), .Y(n444) );
  MUX2X1 U384 ( .B(n448), .A(n449), .S(n1183), .Y(n447) );
  MUX2X1 U385 ( .B(n451), .A(n452), .S(n1183), .Y(n450) );
  MUX2X1 U386 ( .B(n454), .A(n455), .S(n1183), .Y(n453) );
  MUX2X1 U387 ( .B(n457), .A(n458), .S(n1168), .Y(n456) );
  MUX2X1 U388 ( .B(n460), .A(n461), .S(n1184), .Y(n459) );
  MUX2X1 U389 ( .B(n463), .A(n464), .S(n1184), .Y(n462) );
  MUX2X1 U390 ( .B(n466), .A(n467), .S(n1184), .Y(n465) );
  MUX2X1 U391 ( .B(n469), .A(n470), .S(n1184), .Y(n468) );
  MUX2X1 U392 ( .B(n472), .A(n473), .S(n1168), .Y(n471) );
  MUX2X1 U393 ( .B(n475), .A(n476), .S(n1184), .Y(n474) );
  MUX2X1 U394 ( .B(n478), .A(n479), .S(n1184), .Y(n477) );
  MUX2X1 U395 ( .B(n481), .A(n482), .S(n1184), .Y(n480) );
  MUX2X1 U396 ( .B(n484), .A(n485), .S(n1184), .Y(n483) );
  MUX2X1 U397 ( .B(n487), .A(n488), .S(n1168), .Y(n486) );
  MUX2X1 U398 ( .B(n490), .A(n491), .S(n1184), .Y(n489) );
  MUX2X1 U399 ( .B(n493), .A(n494), .S(n1184), .Y(n492) );
  MUX2X1 U400 ( .B(n496), .A(n497), .S(n1184), .Y(n495) );
  MUX2X1 U401 ( .B(n499), .A(n500), .S(n1184), .Y(n498) );
  MUX2X1 U402 ( .B(n502), .A(n503), .S(n1168), .Y(n501) );
  MUX2X1 U403 ( .B(n505), .A(n506), .S(n1185), .Y(n504) );
  MUX2X1 U404 ( .B(n508), .A(n509), .S(n1185), .Y(n507) );
  MUX2X1 U405 ( .B(n511), .A(n512), .S(n1185), .Y(n510) );
  MUX2X1 U406 ( .B(n514), .A(n515), .S(n1185), .Y(n513) );
  MUX2X1 U407 ( .B(n517), .A(n518), .S(n1168), .Y(n516) );
  MUX2X1 U408 ( .B(n520), .A(n521), .S(n1185), .Y(n519) );
  MUX2X1 U409 ( .B(n523), .A(n524), .S(n1185), .Y(n522) );
  MUX2X1 U410 ( .B(n526), .A(n527), .S(n1185), .Y(n525) );
  MUX2X1 U411 ( .B(n529), .A(n530), .S(n1185), .Y(n528) );
  MUX2X1 U412 ( .B(n532), .A(n533), .S(n1168), .Y(n531) );
  MUX2X1 U413 ( .B(n535), .A(n536), .S(n1185), .Y(n534) );
  MUX2X1 U414 ( .B(n538), .A(n539), .S(n1185), .Y(n537) );
  MUX2X1 U415 ( .B(n541), .A(n542), .S(n1185), .Y(n540) );
  MUX2X1 U416 ( .B(n544), .A(n545), .S(n1185), .Y(n543) );
  MUX2X1 U417 ( .B(n547), .A(n548), .S(n1168), .Y(n546) );
  MUX2X1 U418 ( .B(n550), .A(n551), .S(n1186), .Y(n549) );
  MUX2X1 U419 ( .B(n553), .A(n554), .S(n1186), .Y(n552) );
  MUX2X1 U420 ( .B(n556), .A(n557), .S(n1186), .Y(n555) );
  MUX2X1 U421 ( .B(n559), .A(n560), .S(n1186), .Y(n558) );
  MUX2X1 U422 ( .B(n562), .A(n563), .S(n1169), .Y(n561) );
  MUX2X1 U423 ( .B(n565), .A(n566), .S(n1186), .Y(n564) );
  MUX2X1 U424 ( .B(n568), .A(n569), .S(n1186), .Y(n567) );
  MUX2X1 U425 ( .B(n571), .A(n572), .S(n1186), .Y(n570) );
  MUX2X1 U426 ( .B(n574), .A(n575), .S(n1186), .Y(n573) );
  MUX2X1 U427 ( .B(n577), .A(n578), .S(n1169), .Y(n576) );
  MUX2X1 U428 ( .B(n580), .A(n581), .S(n1186), .Y(n579) );
  MUX2X1 U429 ( .B(n583), .A(n584), .S(n1186), .Y(n582) );
  MUX2X1 U430 ( .B(n586), .A(n587), .S(n1186), .Y(n585) );
  MUX2X1 U431 ( .B(n589), .A(n590), .S(n1186), .Y(n588) );
  MUX2X1 U432 ( .B(n592), .A(n593), .S(n1168), .Y(n591) );
  MUX2X1 U433 ( .B(n595), .A(n596), .S(n1187), .Y(n594) );
  MUX2X1 U434 ( .B(n598), .A(n599), .S(n1187), .Y(n597) );
  MUX2X1 U435 ( .B(n601), .A(n602), .S(n1187), .Y(n600) );
  MUX2X1 U436 ( .B(n604), .A(n605), .S(n1187), .Y(n603) );
  MUX2X1 U437 ( .B(n607), .A(n608), .S(n1168), .Y(n606) );
  MUX2X1 U438 ( .B(n610), .A(n611), .S(n1187), .Y(n609) );
  MUX2X1 U439 ( .B(n613), .A(n614), .S(n1187), .Y(n612) );
  MUX2X1 U440 ( .B(n616), .A(n617), .S(n1187), .Y(n615) );
  MUX2X1 U441 ( .B(n619), .A(n620), .S(n1187), .Y(n618) );
  MUX2X1 U442 ( .B(n622), .A(n623), .S(n1169), .Y(n621) );
  MUX2X1 U443 ( .B(n625), .A(n626), .S(n1187), .Y(n624) );
  MUX2X1 U444 ( .B(n628), .A(n629), .S(n1187), .Y(n627) );
  MUX2X1 U445 ( .B(n631), .A(n632), .S(n1187), .Y(n630) );
  MUX2X1 U446 ( .B(n634), .A(n635), .S(n1187), .Y(n633) );
  MUX2X1 U447 ( .B(n637), .A(n638), .S(n1169), .Y(n636) );
  MUX2X1 U448 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1195), .Y(n160) );
  MUX2X1 U449 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1195), .Y(n159) );
  MUX2X1 U450 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1195), .Y(n163) );
  MUX2X1 U451 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1195), .Y(n162) );
  MUX2X1 U452 ( .B(n161), .A(n158), .S(n1174), .Y(n172) );
  MUX2X1 U453 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1196), .Y(n166) );
  MUX2X1 U454 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1196), .Y(n165) );
  MUX2X1 U455 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1196), .Y(n169) );
  MUX2X1 U456 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1196), .Y(n168) );
  MUX2X1 U457 ( .B(n167), .A(n164), .S(n1174), .Y(n171) );
  MUX2X1 U458 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1196), .Y(n175) );
  MUX2X1 U459 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1196), .Y(n174) );
  MUX2X1 U460 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1196), .Y(n178) );
  MUX2X1 U461 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1196), .Y(n177) );
  MUX2X1 U462 ( .B(n176), .A(n173), .S(n1174), .Y(n187) );
  MUX2X1 U463 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1196), .Y(n181) );
  MUX2X1 U464 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1196), .Y(n180) );
  MUX2X1 U465 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1196), .Y(n184) );
  MUX2X1 U466 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1196), .Y(n183) );
  MUX2X1 U467 ( .B(n182), .A(n179), .S(n1174), .Y(n186) );
  MUX2X1 U468 ( .B(n185), .A(n170), .S(n1167), .Y(n639) );
  MUX2X1 U469 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1197), .Y(n190) );
  MUX2X1 U470 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1197), .Y(n189) );
  MUX2X1 U471 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1197), .Y(n193) );
  MUX2X1 U472 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1197), .Y(n192) );
  MUX2X1 U473 ( .B(n191), .A(n188), .S(n1174), .Y(n202) );
  MUX2X1 U474 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1197), .Y(n196) );
  MUX2X1 U475 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1197), .Y(n195) );
  MUX2X1 U476 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1197), .Y(n199) );
  MUX2X1 U477 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1197), .Y(n198) );
  MUX2X1 U478 ( .B(n197), .A(n194), .S(n1174), .Y(n201) );
  MUX2X1 U479 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1197), .Y(n205) );
  MUX2X1 U480 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1197), .Y(n204) );
  MUX2X1 U481 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1197), .Y(n208) );
  MUX2X1 U482 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1197), .Y(n207) );
  MUX2X1 U483 ( .B(n206), .A(n203), .S(n1174), .Y(n218) );
  MUX2X1 U484 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1198), .Y(n211) );
  MUX2X1 U485 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1198), .Y(n210) );
  MUX2X1 U486 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1198), .Y(n215) );
  MUX2X1 U487 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1198), .Y(n213) );
  MUX2X1 U488 ( .B(n212), .A(n209), .S(n1174), .Y(n217) );
  MUX2X1 U489 ( .B(n216), .A(n200), .S(n1167), .Y(n640) );
  MUX2X1 U490 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1198), .Y(n221) );
  MUX2X1 U491 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1198), .Y(n220) );
  MUX2X1 U492 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1198), .Y(n224) );
  MUX2X1 U493 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1198), .Y(n223) );
  MUX2X1 U494 ( .B(n222), .A(n219), .S(n1174), .Y(n233) );
  MUX2X1 U495 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1198), .Y(n227) );
  MUX2X1 U496 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1198), .Y(n226) );
  MUX2X1 U497 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1198), .Y(n230) );
  MUX2X1 U498 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1198), .Y(n229) );
  MUX2X1 U499 ( .B(n228), .A(n225), .S(n1174), .Y(n232) );
  MUX2X1 U500 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1199), .Y(n236) );
  MUX2X1 U501 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1199), .Y(n235) );
  MUX2X1 U502 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1199), .Y(n239) );
  MUX2X1 U503 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1199), .Y(n238) );
  MUX2X1 U504 ( .B(n237), .A(n234), .S(n1174), .Y(n248) );
  MUX2X1 U505 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1199), .Y(n242) );
  MUX2X1 U506 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1199), .Y(n241) );
  MUX2X1 U507 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1199), .Y(n245) );
  MUX2X1 U508 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1199), .Y(n244) );
  MUX2X1 U509 ( .B(n243), .A(n240), .S(n1174), .Y(n247) );
  MUX2X1 U510 ( .B(n246), .A(n231), .S(n1167), .Y(n641) );
  MUX2X1 U511 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1199), .Y(n251) );
  MUX2X1 U512 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1199), .Y(n250) );
  MUX2X1 U513 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1199), .Y(n254) );
  MUX2X1 U514 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1199), .Y(n253) );
  MUX2X1 U515 ( .B(n252), .A(n249), .S(n1173), .Y(n263) );
  MUX2X1 U516 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1200), .Y(n257) );
  MUX2X1 U517 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1200), .Y(n256) );
  MUX2X1 U518 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1200), .Y(n260) );
  MUX2X1 U519 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1200), .Y(n259) );
  MUX2X1 U520 ( .B(n258), .A(n255), .S(n1173), .Y(n262) );
  MUX2X1 U521 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1200), .Y(n266) );
  MUX2X1 U522 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1200), .Y(n265) );
  MUX2X1 U523 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1200), .Y(n269) );
  MUX2X1 U524 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1200), .Y(n268) );
  MUX2X1 U525 ( .B(n267), .A(n264), .S(n1173), .Y(n278) );
  MUX2X1 U526 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1200), .Y(n272) );
  MUX2X1 U527 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1200), .Y(n271) );
  MUX2X1 U528 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1200), .Y(n275) );
  MUX2X1 U529 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1200), .Y(n274) );
  MUX2X1 U530 ( .B(n273), .A(n270), .S(n1173), .Y(n277) );
  MUX2X1 U531 ( .B(n276), .A(n261), .S(n1167), .Y(n642) );
  MUX2X1 U532 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1201), .Y(n281) );
  MUX2X1 U533 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1201), .Y(n280) );
  MUX2X1 U534 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1201), .Y(n284) );
  MUX2X1 U535 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1201), .Y(n283) );
  MUX2X1 U536 ( .B(n282), .A(n279), .S(n1173), .Y(n293) );
  MUX2X1 U537 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1201), .Y(n287) );
  MUX2X1 U538 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1201), .Y(n286) );
  MUX2X1 U539 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1201), .Y(n290) );
  MUX2X1 U540 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1201), .Y(n289) );
  MUX2X1 U541 ( .B(n288), .A(n285), .S(n1173), .Y(n292) );
  MUX2X1 U542 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1201), .Y(n296) );
  MUX2X1 U543 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1201), .Y(n295) );
  MUX2X1 U544 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1201), .Y(n299) );
  MUX2X1 U545 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1201), .Y(n298) );
  MUX2X1 U546 ( .B(n297), .A(n294), .S(n1173), .Y(n308) );
  MUX2X1 U547 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1202), .Y(n302) );
  MUX2X1 U548 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1202), .Y(n301) );
  MUX2X1 U549 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1202), .Y(n305) );
  MUX2X1 U550 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1202), .Y(n304) );
  MUX2X1 U551 ( .B(n303), .A(n300), .S(n1173), .Y(n307) );
  MUX2X1 U552 ( .B(n306), .A(n291), .S(n1167), .Y(n643) );
  MUX2X1 U553 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1202), .Y(n311) );
  MUX2X1 U554 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1202), .Y(n310) );
  MUX2X1 U555 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1202), .Y(n314) );
  MUX2X1 U556 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1202), .Y(n313) );
  MUX2X1 U557 ( .B(n312), .A(n309), .S(n1173), .Y(n323) );
  MUX2X1 U558 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1202), .Y(n317) );
  MUX2X1 U559 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1202), .Y(n316) );
  MUX2X1 U560 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1202), .Y(n320) );
  MUX2X1 U561 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1202), .Y(n319) );
  MUX2X1 U562 ( .B(n318), .A(n315), .S(n1173), .Y(n322) );
  MUX2X1 U563 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1203), .Y(n326) );
  MUX2X1 U564 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1203), .Y(n325) );
  MUX2X1 U565 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1203), .Y(n329) );
  MUX2X1 U566 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1203), .Y(n328) );
  MUX2X1 U567 ( .B(n327), .A(n324), .S(n1173), .Y(n338) );
  MUX2X1 U568 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1203), .Y(n332) );
  MUX2X1 U569 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1203), .Y(n331) );
  MUX2X1 U570 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1203), .Y(n335) );
  MUX2X1 U571 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1203), .Y(n334) );
  MUX2X1 U572 ( .B(n333), .A(n330), .S(n1173), .Y(n337) );
  MUX2X1 U573 ( .B(n336), .A(n321), .S(n1167), .Y(n644) );
  MUX2X1 U574 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1203), .Y(n341) );
  MUX2X1 U575 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1203), .Y(n340) );
  MUX2X1 U576 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1203), .Y(n344) );
  MUX2X1 U577 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1203), .Y(n343) );
  MUX2X1 U578 ( .B(n342), .A(n339), .S(n1172), .Y(n353) );
  MUX2X1 U579 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1204), .Y(n347) );
  MUX2X1 U580 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1204), .Y(n346) );
  MUX2X1 U581 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1204), .Y(n350) );
  MUX2X1 U582 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1204), .Y(n349) );
  MUX2X1 U583 ( .B(n348), .A(n345), .S(n1172), .Y(n352) );
  MUX2X1 U584 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1204), .Y(n356) );
  MUX2X1 U585 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1204), .Y(n355) );
  MUX2X1 U586 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1204), .Y(n359) );
  MUX2X1 U587 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1204), .Y(n358) );
  MUX2X1 U588 ( .B(n357), .A(n354), .S(n1172), .Y(n368) );
  MUX2X1 U589 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1204), .Y(n362) );
  MUX2X1 U590 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1204), .Y(n361) );
  MUX2X1 U591 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1204), .Y(n365) );
  MUX2X1 U592 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1204), .Y(n364) );
  MUX2X1 U593 ( .B(n363), .A(n360), .S(n1172), .Y(n367) );
  MUX2X1 U594 ( .B(n366), .A(n351), .S(n1167), .Y(n645) );
  MUX2X1 U595 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1205), .Y(n371) );
  MUX2X1 U596 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1205), .Y(n370) );
  MUX2X1 U597 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1205), .Y(n374) );
  MUX2X1 U598 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1205), .Y(n373) );
  MUX2X1 U599 ( .B(n372), .A(n369), .S(n1172), .Y(n383) );
  MUX2X1 U600 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1205), .Y(n377) );
  MUX2X1 U601 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1205), .Y(n376) );
  MUX2X1 U602 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1205), .Y(n380) );
  MUX2X1 U603 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1205), .Y(n379) );
  MUX2X1 U604 ( .B(n378), .A(n375), .S(n1172), .Y(n382) );
  MUX2X1 U605 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1205), .Y(n386) );
  MUX2X1 U606 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1205), .Y(n385) );
  MUX2X1 U607 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1205), .Y(n389) );
  MUX2X1 U608 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1205), .Y(n388) );
  MUX2X1 U609 ( .B(n387), .A(n384), .S(n1172), .Y(n398) );
  MUX2X1 U610 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1206), .Y(n392) );
  MUX2X1 U611 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1206), .Y(n391) );
  MUX2X1 U612 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1206), .Y(n395) );
  MUX2X1 U613 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1206), .Y(n394) );
  MUX2X1 U614 ( .B(n393), .A(n390), .S(n1172), .Y(n397) );
  MUX2X1 U615 ( .B(n396), .A(n381), .S(n1167), .Y(n646) );
  MUX2X1 U616 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1206), .Y(n401) );
  MUX2X1 U617 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1206), .Y(n400) );
  MUX2X1 U618 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1206), .Y(n404) );
  MUX2X1 U619 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1206), .Y(n403) );
  MUX2X1 U620 ( .B(n402), .A(n399), .S(n1172), .Y(n413) );
  MUX2X1 U621 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1206), .Y(n407) );
  MUX2X1 U622 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1206), .Y(n406) );
  MUX2X1 U623 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1206), .Y(n410) );
  MUX2X1 U624 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1206), .Y(n409) );
  MUX2X1 U625 ( .B(n408), .A(n405), .S(n1172), .Y(n412) );
  MUX2X1 U626 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1207), .Y(n416) );
  MUX2X1 U627 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1207), .Y(n415) );
  MUX2X1 U628 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1207), .Y(n419) );
  MUX2X1 U629 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1207), .Y(n418) );
  MUX2X1 U630 ( .B(n417), .A(n414), .S(n1172), .Y(n428) );
  MUX2X1 U631 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1207), .Y(n422) );
  MUX2X1 U632 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1207), .Y(n421) );
  MUX2X1 U633 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1207), .Y(n425) );
  MUX2X1 U634 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1207), .Y(n424) );
  MUX2X1 U635 ( .B(n423), .A(n420), .S(n1172), .Y(n427) );
  MUX2X1 U636 ( .B(n426), .A(n411), .S(n1167), .Y(n647) );
  MUX2X1 U637 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1207), .Y(n431) );
  MUX2X1 U638 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1207), .Y(n430) );
  MUX2X1 U639 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1207), .Y(n434) );
  MUX2X1 U640 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1207), .Y(n433) );
  MUX2X1 U641 ( .B(n432), .A(n429), .S(n1171), .Y(n443) );
  MUX2X1 U642 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1208), .Y(n437) );
  MUX2X1 U643 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1208), .Y(n436) );
  MUX2X1 U644 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1208), .Y(n440) );
  MUX2X1 U645 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1208), .Y(n439) );
  MUX2X1 U646 ( .B(n438), .A(n435), .S(n1171), .Y(n442) );
  MUX2X1 U647 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1208), .Y(n446) );
  MUX2X1 U648 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1208), .Y(n445) );
  MUX2X1 U649 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1208), .Y(n449) );
  MUX2X1 U650 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1208), .Y(n448) );
  MUX2X1 U651 ( .B(n447), .A(n444), .S(n1171), .Y(n458) );
  MUX2X1 U652 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1208), .Y(n452) );
  MUX2X1 U653 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1208), .Y(n451) );
  MUX2X1 U654 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1208), .Y(n455) );
  MUX2X1 U655 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1208), .Y(n454) );
  MUX2X1 U656 ( .B(n453), .A(n450), .S(n1171), .Y(n457) );
  MUX2X1 U657 ( .B(n456), .A(n441), .S(n1167), .Y(n648) );
  MUX2X1 U658 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1209), .Y(n461) );
  MUX2X1 U659 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1209), .Y(n460) );
  MUX2X1 U660 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1209), .Y(n464) );
  MUX2X1 U661 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1209), .Y(n463) );
  MUX2X1 U662 ( .B(n462), .A(n459), .S(n1171), .Y(n473) );
  MUX2X1 U663 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1209), .Y(n467) );
  MUX2X1 U664 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1209), .Y(n466) );
  MUX2X1 U665 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1209), .Y(n470) );
  MUX2X1 U666 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1209), .Y(n469) );
  MUX2X1 U667 ( .B(n468), .A(n465), .S(n1171), .Y(n472) );
  MUX2X1 U668 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1209), .Y(n476) );
  MUX2X1 U669 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1209), .Y(n475) );
  MUX2X1 U670 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1209), .Y(n479) );
  MUX2X1 U671 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1209), .Y(n478) );
  MUX2X1 U672 ( .B(n477), .A(n474), .S(n1171), .Y(n488) );
  MUX2X1 U673 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1210), .Y(n482) );
  MUX2X1 U674 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1210), .Y(n481) );
  MUX2X1 U675 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1210), .Y(n485) );
  MUX2X1 U676 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1210), .Y(n484) );
  MUX2X1 U677 ( .B(n483), .A(n480), .S(n1171), .Y(n487) );
  MUX2X1 U678 ( .B(n486), .A(n471), .S(n1167), .Y(n649) );
  MUX2X1 U679 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1210), .Y(n491) );
  MUX2X1 U680 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1210), .Y(n490) );
  MUX2X1 U681 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1210), .Y(n494) );
  MUX2X1 U682 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1210), .Y(n493) );
  MUX2X1 U683 ( .B(n492), .A(n489), .S(n1171), .Y(n503) );
  MUX2X1 U684 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1210), .Y(n497) );
  MUX2X1 U685 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1210), .Y(n496) );
  MUX2X1 U686 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1210), .Y(n500) );
  MUX2X1 U687 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1210), .Y(n499) );
  MUX2X1 U688 ( .B(n498), .A(n495), .S(n1171), .Y(n502) );
  MUX2X1 U689 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1211), .Y(n506) );
  MUX2X1 U690 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1211), .Y(n505) );
  MUX2X1 U691 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1211), .Y(n509) );
  MUX2X1 U692 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1211), .Y(n508) );
  MUX2X1 U693 ( .B(n507), .A(n504), .S(n1171), .Y(n518) );
  MUX2X1 U694 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1211), .Y(n512) );
  MUX2X1 U695 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1211), .Y(n511) );
  MUX2X1 U696 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1211), .Y(n515) );
  MUX2X1 U697 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1211), .Y(n514) );
  MUX2X1 U698 ( .B(n513), .A(n510), .S(n1171), .Y(n517) );
  MUX2X1 U699 ( .B(n516), .A(n501), .S(n1167), .Y(n650) );
  MUX2X1 U700 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1211), .Y(n521) );
  MUX2X1 U701 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1211), .Y(n520) );
  MUX2X1 U702 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1211), .Y(n524) );
  MUX2X1 U703 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1211), .Y(n523) );
  MUX2X1 U704 ( .B(n522), .A(n519), .S(n1170), .Y(n533) );
  MUX2X1 U705 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1212), .Y(n527) );
  MUX2X1 U706 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1212), .Y(n526) );
  MUX2X1 U707 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1212), .Y(n530) );
  MUX2X1 U708 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1212), .Y(n529) );
  MUX2X1 U709 ( .B(n528), .A(n525), .S(n1170), .Y(n532) );
  MUX2X1 U710 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1212), .Y(n536) );
  MUX2X1 U711 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1212), .Y(n535) );
  MUX2X1 U712 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1212), .Y(n539) );
  MUX2X1 U713 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1212), .Y(n538) );
  MUX2X1 U714 ( .B(n537), .A(n534), .S(n1170), .Y(n548) );
  MUX2X1 U715 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1212), .Y(n542) );
  MUX2X1 U716 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1212), .Y(n541) );
  MUX2X1 U717 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1212), .Y(n545) );
  MUX2X1 U718 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1212), .Y(n544) );
  MUX2X1 U719 ( .B(n543), .A(n540), .S(n1170), .Y(n547) );
  MUX2X1 U720 ( .B(n546), .A(n531), .S(n1167), .Y(n1163) );
  MUX2X1 U721 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1213), .Y(n551) );
  MUX2X1 U722 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1213), .Y(n550) );
  MUX2X1 U723 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1213), .Y(n554) );
  MUX2X1 U724 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1213), .Y(n553) );
  MUX2X1 U725 ( .B(n552), .A(n549), .S(n1170), .Y(n563) );
  MUX2X1 U726 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1213), .Y(n557) );
  MUX2X1 U727 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1213), .Y(n556) );
  MUX2X1 U728 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1213), .Y(n560) );
  MUX2X1 U729 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1213), .Y(n559) );
  MUX2X1 U730 ( .B(n558), .A(n555), .S(n1170), .Y(n562) );
  MUX2X1 U731 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1213), .Y(n566) );
  MUX2X1 U732 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1213), .Y(n565) );
  MUX2X1 U733 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1213), .Y(n569) );
  MUX2X1 U734 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1213), .Y(n568) );
  MUX2X1 U735 ( .B(n567), .A(n564), .S(n1170), .Y(n578) );
  MUX2X1 U736 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1214), .Y(n572) );
  MUX2X1 U737 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1214), .Y(n571) );
  MUX2X1 U738 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1214), .Y(n575) );
  MUX2X1 U739 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1214), .Y(n574) );
  MUX2X1 U740 ( .B(n573), .A(n570), .S(n1170), .Y(n577) );
  MUX2X1 U741 ( .B(n576), .A(n561), .S(n1167), .Y(n1164) );
  MUX2X1 U742 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1214), .Y(n581) );
  MUX2X1 U743 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1214), .Y(n580) );
  MUX2X1 U744 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1214), .Y(n584) );
  MUX2X1 U745 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1214), .Y(n583) );
  MUX2X1 U746 ( .B(n582), .A(n579), .S(n1170), .Y(n593) );
  MUX2X1 U747 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1214), .Y(n587) );
  MUX2X1 U748 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1214), .Y(n586) );
  MUX2X1 U749 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1214), .Y(n590) );
  MUX2X1 U750 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1214), .Y(n589) );
  MUX2X1 U751 ( .B(n588), .A(n585), .S(n1170), .Y(n592) );
  MUX2X1 U752 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1215), .Y(n596) );
  MUX2X1 U753 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1215), .Y(n595) );
  MUX2X1 U754 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1215), .Y(n599) );
  MUX2X1 U755 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1215), .Y(n598) );
  MUX2X1 U756 ( .B(n597), .A(n594), .S(n1170), .Y(n608) );
  MUX2X1 U757 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1215), .Y(n602) );
  MUX2X1 U758 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1215), .Y(n601) );
  MUX2X1 U759 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1215), .Y(n605) );
  MUX2X1 U760 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1215), .Y(n604) );
  MUX2X1 U761 ( .B(n603), .A(n600), .S(n1170), .Y(n607) );
  MUX2X1 U762 ( .B(n606), .A(n591), .S(n1167), .Y(n1165) );
  MUX2X1 U763 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1215), .Y(n611) );
  MUX2X1 U764 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1215), .Y(n610) );
  MUX2X1 U765 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1215), .Y(n614) );
  MUX2X1 U766 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1215), .Y(n613) );
  MUX2X1 U767 ( .B(n612), .A(n609), .S(n1170), .Y(n623) );
  MUX2X1 U768 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1216), .Y(n617) );
  MUX2X1 U769 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1216), .Y(n616) );
  MUX2X1 U770 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1216), .Y(n620) );
  MUX2X1 U771 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1216), .Y(n619) );
  MUX2X1 U772 ( .B(n618), .A(n615), .S(n1171), .Y(n622) );
  MUX2X1 U773 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1216), .Y(n626) );
  MUX2X1 U774 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1216), .Y(n625) );
  MUX2X1 U775 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1216), .Y(n629) );
  MUX2X1 U776 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1216), .Y(n628) );
  MUX2X1 U777 ( .B(n627), .A(n624), .S(n1170), .Y(n638) );
  MUX2X1 U778 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1216), .Y(n632) );
  MUX2X1 U779 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1216), .Y(n631) );
  MUX2X1 U780 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1216), .Y(n635) );
  MUX2X1 U781 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1216), .Y(n634) );
  MUX2X1 U782 ( .B(n633), .A(n630), .S(n1171), .Y(n637) );
  MUX2X1 U783 ( .B(n636), .A(n621), .S(n1167), .Y(n1166) );
  INVX8 U784 ( .A(n1194), .Y(n1197) );
  INVX8 U785 ( .A(n1193), .Y(n1199) );
  INVX8 U786 ( .A(n1193), .Y(n1200) );
  INVX8 U787 ( .A(n1192), .Y(n1203) );
  INVX8 U788 ( .A(n1191), .Y(n1204) );
  INVX8 U789 ( .A(n1191), .Y(n1205) );
  INVX8 U790 ( .A(n1191), .Y(n1206) );
  INVX8 U791 ( .A(n1190), .Y(n1207) );
  INVX8 U792 ( .A(n1190), .Y(n1208) );
  INVX8 U793 ( .A(n1190), .Y(n1209) );
  INVX8 U794 ( .A(n1189), .Y(n1210) );
  INVX8 U795 ( .A(n1189), .Y(n1211) );
  INVX8 U796 ( .A(n1189), .Y(n1212) );
  INVX8 U797 ( .A(n1189), .Y(n1213) );
  INVX8 U798 ( .A(n1189), .Y(n1214) );
  INVX8 U799 ( .A(n1189), .Y(n1215) );
  INVX8 U800 ( .A(n1189), .Y(n1216) );
  INVX1 U801 ( .A(N11), .Y(n1319) );
  INVX1 U802 ( .A(N10), .Y(n1317) );
  INVX8 U803 ( .A(n1282), .Y(n1280) );
  INVX8 U804 ( .A(n1282), .Y(n1281) );
  INVX8 U805 ( .A(n4), .Y(n1283) );
  INVX8 U806 ( .A(n4), .Y(n1284) );
  INVX8 U807 ( .A(n5), .Y(n1285) );
  INVX8 U808 ( .A(n5), .Y(n1286) );
  INVX8 U809 ( .A(n6), .Y(n1287) );
  INVX8 U810 ( .A(n6), .Y(n1288) );
  INVX8 U811 ( .A(n7), .Y(n1289) );
  INVX8 U812 ( .A(n7), .Y(n1290) );
  INVX8 U813 ( .A(n8), .Y(n1291) );
  INVX8 U814 ( .A(n8), .Y(n1292) );
  INVX8 U815 ( .A(n9), .Y(n1293) );
  INVX8 U816 ( .A(n9), .Y(n1294) );
  INVX8 U817 ( .A(n10), .Y(n1295) );
  INVX8 U818 ( .A(n10), .Y(n1296) );
  INVX8 U819 ( .A(n11), .Y(n1297) );
  INVX8 U820 ( .A(n11), .Y(n1298) );
  INVX8 U821 ( .A(n12), .Y(n1299) );
  INVX8 U822 ( .A(n12), .Y(n1300) );
  INVX8 U823 ( .A(n13), .Y(n1301) );
  INVX8 U824 ( .A(n13), .Y(n1302) );
  INVX8 U825 ( .A(n14), .Y(n1303) );
  INVX8 U826 ( .A(n14), .Y(n1304) );
  INVX8 U827 ( .A(n86), .Y(n1305) );
  INVX8 U828 ( .A(n86), .Y(n1306) );
  INVX8 U829 ( .A(n78), .Y(n1307) );
  INVX8 U830 ( .A(n78), .Y(n1308) );
  INVX8 U831 ( .A(n79), .Y(n1309) );
  INVX8 U832 ( .A(n79), .Y(n1310) );
  INVX8 U833 ( .A(n80), .Y(n1311) );
  INVX8 U834 ( .A(n80), .Y(n1312) );
  INVX8 U835 ( .A(n81), .Y(n1313) );
  INVX8 U836 ( .A(n81), .Y(n1314) );
  AND2X2 U837 ( .A(N32), .B(n3), .Y(\data_out<0> ) );
  AND2X2 U838 ( .A(n3), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U839 ( .A(n1), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U840 ( .A(n1), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U841 ( .A(n1), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U842 ( .A(n1), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U843 ( .A(N26), .B(n3), .Y(\data_out<6> ) );
  AND2X2 U844 ( .A(n3), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U845 ( .A(n1), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U846 ( .A(n1), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U847 ( .A(n1), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U848 ( .A(N21), .B(n3), .Y(\data_out<11> ) );
  AND2X2 U849 ( .A(N20), .B(n3), .Y(\data_out<12> ) );
  AND2X2 U850 ( .A(n1), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U851 ( .A(n1), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U852 ( .A(n1), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U853 ( .A(\mem<31><0> ), .B(n33), .Y(n1326) );
  OAI21X1 U854 ( .A(n1221), .B(n1283), .C(n1326), .Y(n2364) );
  NAND2X1 U855 ( .A(\mem<31><1> ), .B(n33), .Y(n1327) );
  OAI21X1 U856 ( .A(n1286), .B(n1220), .C(n1327), .Y(n2363) );
  NAND2X1 U857 ( .A(\mem<31><2> ), .B(n33), .Y(n1328) );
  OAI21X1 U858 ( .A(n1288), .B(n1220), .C(n1328), .Y(n2362) );
  NAND2X1 U859 ( .A(\mem<31><3> ), .B(n33), .Y(n1329) );
  OAI21X1 U860 ( .A(n1290), .B(n1220), .C(n1329), .Y(n2361) );
  NAND2X1 U861 ( .A(\mem<31><4> ), .B(n33), .Y(n1330) );
  OAI21X1 U862 ( .A(n1292), .B(n1220), .C(n1330), .Y(n2360) );
  NAND2X1 U863 ( .A(\mem<31><5> ), .B(n33), .Y(n1331) );
  OAI21X1 U864 ( .A(n1294), .B(n1220), .C(n1331), .Y(n2359) );
  NAND2X1 U865 ( .A(\mem<31><6> ), .B(n33), .Y(n1332) );
  OAI21X1 U866 ( .A(n1296), .B(n1220), .C(n1332), .Y(n2358) );
  NAND2X1 U867 ( .A(\mem<31><7> ), .B(n33), .Y(n1333) );
  OAI21X1 U868 ( .A(n1298), .B(n1220), .C(n1333), .Y(n2357) );
  NAND2X1 U869 ( .A(\mem<31><8> ), .B(n33), .Y(n1334) );
  OAI21X1 U870 ( .A(n1300), .B(n1220), .C(n1334), .Y(n2356) );
  NAND2X1 U871 ( .A(\mem<31><9> ), .B(n33), .Y(n1335) );
  OAI21X1 U872 ( .A(n1302), .B(n1221), .C(n1335), .Y(n2355) );
  NAND2X1 U873 ( .A(\mem<31><10> ), .B(n33), .Y(n1336) );
  OAI21X1 U874 ( .A(n1304), .B(n1221), .C(n1336), .Y(n2354) );
  NAND2X1 U875 ( .A(\mem<31><11> ), .B(n33), .Y(n1337) );
  OAI21X1 U876 ( .A(n1306), .B(n1221), .C(n1337), .Y(n2353) );
  NAND2X1 U877 ( .A(\mem<31><12> ), .B(n33), .Y(n1338) );
  OAI21X1 U878 ( .A(n1308), .B(n1221), .C(n1338), .Y(n2352) );
  NAND2X1 U879 ( .A(\mem<31><13> ), .B(n33), .Y(n1339) );
  OAI21X1 U880 ( .A(n1310), .B(n1221), .C(n1339), .Y(n2351) );
  NAND2X1 U881 ( .A(\mem<31><14> ), .B(n33), .Y(n1340) );
  OAI21X1 U882 ( .A(n1312), .B(n1221), .C(n1340), .Y(n2350) );
  NAND2X1 U883 ( .A(\mem<31><15> ), .B(n33), .Y(n1341) );
  OAI21X1 U884 ( .A(n1314), .B(n1221), .C(n1341), .Y(n2349) );
  NAND2X1 U885 ( .A(\mem<30><0> ), .B(n39), .Y(n1342) );
  OAI21X1 U886 ( .A(n1222), .B(n1283), .C(n1342), .Y(n2348) );
  NAND2X1 U887 ( .A(\mem<30><1> ), .B(n39), .Y(n1343) );
  OAI21X1 U888 ( .A(n1222), .B(n1286), .C(n1343), .Y(n2347) );
  NAND2X1 U889 ( .A(\mem<30><2> ), .B(n39), .Y(n1344) );
  OAI21X1 U890 ( .A(n1222), .B(n1288), .C(n1344), .Y(n2346) );
  NAND2X1 U891 ( .A(\mem<30><3> ), .B(n39), .Y(n1345) );
  OAI21X1 U892 ( .A(n1222), .B(n1290), .C(n1345), .Y(n2345) );
  NAND2X1 U893 ( .A(\mem<30><4> ), .B(n39), .Y(n1346) );
  OAI21X1 U894 ( .A(n1222), .B(n1292), .C(n1346), .Y(n2344) );
  NAND2X1 U895 ( .A(\mem<30><5> ), .B(n39), .Y(n1347) );
  OAI21X1 U896 ( .A(n1222), .B(n1294), .C(n1347), .Y(n2343) );
  NAND2X1 U897 ( .A(\mem<30><6> ), .B(n39), .Y(n1348) );
  OAI21X1 U898 ( .A(n1222), .B(n1296), .C(n1348), .Y(n2342) );
  NAND2X1 U899 ( .A(\mem<30><7> ), .B(n39), .Y(n1349) );
  OAI21X1 U900 ( .A(n1222), .B(n1298), .C(n1349), .Y(n2341) );
  NAND2X1 U901 ( .A(\mem<30><8> ), .B(n39), .Y(n1350) );
  OAI21X1 U902 ( .A(n1223), .B(n1299), .C(n1350), .Y(n2340) );
  NAND2X1 U903 ( .A(\mem<30><9> ), .B(n39), .Y(n1351) );
  OAI21X1 U904 ( .A(n1223), .B(n1301), .C(n1351), .Y(n2339) );
  NAND2X1 U905 ( .A(\mem<30><10> ), .B(n39), .Y(n1352) );
  OAI21X1 U906 ( .A(n1223), .B(n1303), .C(n1352), .Y(n2338) );
  NAND2X1 U907 ( .A(\mem<30><11> ), .B(n39), .Y(n1353) );
  OAI21X1 U908 ( .A(n1223), .B(n1305), .C(n1353), .Y(n2337) );
  NAND2X1 U909 ( .A(\mem<30><12> ), .B(n39), .Y(n1354) );
  OAI21X1 U910 ( .A(n1223), .B(n1307), .C(n1354), .Y(n2336) );
  NAND2X1 U911 ( .A(\mem<30><13> ), .B(n39), .Y(n1355) );
  OAI21X1 U912 ( .A(n1223), .B(n1309), .C(n1355), .Y(n2335) );
  NAND2X1 U913 ( .A(\mem<30><14> ), .B(n39), .Y(n1356) );
  OAI21X1 U914 ( .A(n1223), .B(n1311), .C(n1356), .Y(n2334) );
  NAND2X1 U915 ( .A(\mem<30><15> ), .B(n39), .Y(n1357) );
  OAI21X1 U916 ( .A(n1223), .B(n1313), .C(n1357), .Y(n2333) );
  NAND3X1 U917 ( .A(n1316), .B(n1320), .C(n1319), .Y(n1358) );
  NAND2X1 U918 ( .A(\mem<29><0> ), .B(n41), .Y(n1359) );
  OAI21X1 U919 ( .A(n1224), .B(n1283), .C(n1359), .Y(n2332) );
  NAND2X1 U920 ( .A(\mem<29><1> ), .B(n41), .Y(n1360) );
  OAI21X1 U921 ( .A(n1224), .B(n1285), .C(n1360), .Y(n2331) );
  NAND2X1 U922 ( .A(\mem<29><2> ), .B(n41), .Y(n1361) );
  OAI21X1 U923 ( .A(n1224), .B(n1287), .C(n1361), .Y(n2330) );
  NAND2X1 U924 ( .A(\mem<29><3> ), .B(n41), .Y(n1362) );
  OAI21X1 U925 ( .A(n1224), .B(n1289), .C(n1362), .Y(n2329) );
  NAND2X1 U926 ( .A(\mem<29><4> ), .B(n41), .Y(n1363) );
  OAI21X1 U927 ( .A(n1224), .B(n1291), .C(n1363), .Y(n2328) );
  NAND2X1 U928 ( .A(\mem<29><5> ), .B(n41), .Y(n1364) );
  OAI21X1 U929 ( .A(n1224), .B(n1293), .C(n1364), .Y(n2327) );
  NAND2X1 U930 ( .A(\mem<29><6> ), .B(n41), .Y(n1365) );
  OAI21X1 U931 ( .A(n1224), .B(n1295), .C(n1365), .Y(n2326) );
  NAND2X1 U932 ( .A(\mem<29><7> ), .B(n41), .Y(n1366) );
  OAI21X1 U933 ( .A(n1224), .B(n1297), .C(n1366), .Y(n2325) );
  NAND2X1 U934 ( .A(\mem<29><8> ), .B(n41), .Y(n1367) );
  OAI21X1 U935 ( .A(n1225), .B(n1300), .C(n1367), .Y(n2324) );
  NAND2X1 U936 ( .A(\mem<29><9> ), .B(n41), .Y(n1368) );
  OAI21X1 U937 ( .A(n1225), .B(n1302), .C(n1368), .Y(n2323) );
  NAND2X1 U938 ( .A(\mem<29><10> ), .B(n41), .Y(n1369) );
  OAI21X1 U939 ( .A(n1225), .B(n1304), .C(n1369), .Y(n2322) );
  NAND2X1 U940 ( .A(\mem<29><11> ), .B(n41), .Y(n1370) );
  OAI21X1 U941 ( .A(n1225), .B(n1306), .C(n1370), .Y(n2321) );
  NAND2X1 U942 ( .A(\mem<29><12> ), .B(n41), .Y(n1371) );
  OAI21X1 U943 ( .A(n1225), .B(n1308), .C(n1371), .Y(n2320) );
  NAND2X1 U944 ( .A(\mem<29><13> ), .B(n41), .Y(n1372) );
  OAI21X1 U945 ( .A(n1225), .B(n1310), .C(n1372), .Y(n2319) );
  NAND2X1 U946 ( .A(\mem<29><14> ), .B(n41), .Y(n1373) );
  OAI21X1 U947 ( .A(n1225), .B(n1312), .C(n1373), .Y(n2318) );
  NAND2X1 U948 ( .A(\mem<29><15> ), .B(n41), .Y(n1374) );
  OAI21X1 U949 ( .A(n1225), .B(n1314), .C(n1374), .Y(n2317) );
  NAND3X1 U950 ( .A(n1320), .B(n1319), .C(n1317), .Y(n1375) );
  NAND2X1 U951 ( .A(\mem<28><0> ), .B(n43), .Y(n1376) );
  OAI21X1 U952 ( .A(n1226), .B(n1283), .C(n1376), .Y(n2316) );
  NAND2X1 U953 ( .A(\mem<28><1> ), .B(n43), .Y(n1377) );
  OAI21X1 U954 ( .A(n1226), .B(n1286), .C(n1377), .Y(n2315) );
  NAND2X1 U955 ( .A(\mem<28><2> ), .B(n43), .Y(n1378) );
  OAI21X1 U956 ( .A(n1226), .B(n1288), .C(n1378), .Y(n2314) );
  NAND2X1 U957 ( .A(\mem<28><3> ), .B(n43), .Y(n1379) );
  OAI21X1 U958 ( .A(n1226), .B(n1290), .C(n1379), .Y(n2313) );
  NAND2X1 U959 ( .A(\mem<28><4> ), .B(n43), .Y(n1380) );
  OAI21X1 U960 ( .A(n1226), .B(n1292), .C(n1380), .Y(n2312) );
  NAND2X1 U961 ( .A(\mem<28><5> ), .B(n43), .Y(n1381) );
  OAI21X1 U962 ( .A(n1226), .B(n1294), .C(n1381), .Y(n2311) );
  NAND2X1 U963 ( .A(\mem<28><6> ), .B(n43), .Y(n1382) );
  OAI21X1 U964 ( .A(n1226), .B(n1296), .C(n1382), .Y(n2310) );
  NAND2X1 U965 ( .A(\mem<28><7> ), .B(n43), .Y(n1383) );
  OAI21X1 U966 ( .A(n1226), .B(n1298), .C(n1383), .Y(n2309) );
  NAND2X1 U967 ( .A(\mem<28><8> ), .B(n43), .Y(n1384) );
  OAI21X1 U968 ( .A(n1227), .B(n1299), .C(n1384), .Y(n2308) );
  NAND2X1 U969 ( .A(\mem<28><9> ), .B(n43), .Y(n1385) );
  OAI21X1 U970 ( .A(n1227), .B(n1301), .C(n1385), .Y(n2307) );
  NAND2X1 U971 ( .A(\mem<28><10> ), .B(n43), .Y(n1386) );
  OAI21X1 U972 ( .A(n1227), .B(n1303), .C(n1386), .Y(n2306) );
  NAND2X1 U973 ( .A(\mem<28><11> ), .B(n43), .Y(n1387) );
  OAI21X1 U974 ( .A(n1227), .B(n1305), .C(n1387), .Y(n2305) );
  NAND2X1 U975 ( .A(\mem<28><12> ), .B(n43), .Y(n1388) );
  OAI21X1 U976 ( .A(n1227), .B(n1307), .C(n1388), .Y(n2304) );
  NAND2X1 U977 ( .A(\mem<28><13> ), .B(n43), .Y(n1389) );
  OAI21X1 U978 ( .A(n1227), .B(n1309), .C(n1389), .Y(n2303) );
  NAND2X1 U979 ( .A(\mem<28><14> ), .B(n43), .Y(n1390) );
  OAI21X1 U980 ( .A(n1227), .B(n1311), .C(n1390), .Y(n2302) );
  NAND2X1 U981 ( .A(\mem<28><15> ), .B(n43), .Y(n1391) );
  OAI21X1 U982 ( .A(n1227), .B(n1313), .C(n1391), .Y(n2301) );
  NAND3X1 U983 ( .A(n1316), .B(n1318), .C(n1321), .Y(n1392) );
  NAND2X1 U984 ( .A(\mem<27><0> ), .B(n19), .Y(n1393) );
  OAI21X1 U985 ( .A(n1228), .B(n1283), .C(n1393), .Y(n2300) );
  NAND2X1 U986 ( .A(\mem<27><1> ), .B(n19), .Y(n1394) );
  OAI21X1 U987 ( .A(n1228), .B(n1285), .C(n1394), .Y(n2299) );
  NAND2X1 U988 ( .A(\mem<27><2> ), .B(n19), .Y(n1395) );
  OAI21X1 U989 ( .A(n1228), .B(n1287), .C(n1395), .Y(n2298) );
  NAND2X1 U990 ( .A(\mem<27><3> ), .B(n19), .Y(n1396) );
  OAI21X1 U991 ( .A(n1228), .B(n1289), .C(n1396), .Y(n2297) );
  NAND2X1 U992 ( .A(\mem<27><4> ), .B(n19), .Y(n1397) );
  OAI21X1 U993 ( .A(n1228), .B(n1291), .C(n1397), .Y(n2296) );
  NAND2X1 U994 ( .A(\mem<27><5> ), .B(n19), .Y(n1398) );
  OAI21X1 U995 ( .A(n1228), .B(n1293), .C(n1398), .Y(n2295) );
  NAND2X1 U996 ( .A(\mem<27><6> ), .B(n19), .Y(n1399) );
  OAI21X1 U997 ( .A(n1228), .B(n1295), .C(n1399), .Y(n2294) );
  NAND2X1 U998 ( .A(\mem<27><7> ), .B(n19), .Y(n1400) );
  OAI21X1 U999 ( .A(n1228), .B(n1297), .C(n1400), .Y(n2293) );
  NAND2X1 U1000 ( .A(\mem<27><8> ), .B(n19), .Y(n1401) );
  OAI21X1 U1001 ( .A(n1229), .B(n1300), .C(n1401), .Y(n2292) );
  NAND2X1 U1002 ( .A(\mem<27><9> ), .B(n19), .Y(n1402) );
  OAI21X1 U1003 ( .A(n1229), .B(n1302), .C(n1402), .Y(n2291) );
  NAND2X1 U1004 ( .A(\mem<27><10> ), .B(n19), .Y(n1403) );
  OAI21X1 U1005 ( .A(n1229), .B(n1304), .C(n1403), .Y(n2290) );
  NAND2X1 U1006 ( .A(\mem<27><11> ), .B(n19), .Y(n1404) );
  OAI21X1 U1007 ( .A(n1229), .B(n1306), .C(n1404), .Y(n2289) );
  NAND2X1 U1008 ( .A(\mem<27><12> ), .B(n19), .Y(n1405) );
  OAI21X1 U1009 ( .A(n1229), .B(n1308), .C(n1405), .Y(n2288) );
  NAND2X1 U1010 ( .A(\mem<27><13> ), .B(n19), .Y(n1406) );
  OAI21X1 U1011 ( .A(n1229), .B(n1310), .C(n1406), .Y(n2287) );
  NAND2X1 U1012 ( .A(\mem<27><14> ), .B(n19), .Y(n1407) );
  OAI21X1 U1013 ( .A(n1229), .B(n1312), .C(n1407), .Y(n2286) );
  NAND2X1 U1014 ( .A(\mem<27><15> ), .B(n19), .Y(n1408) );
  OAI21X1 U1015 ( .A(n1229), .B(n1314), .C(n1408), .Y(n2285) );
  NAND3X1 U1016 ( .A(n1321), .B(n1318), .C(n1317), .Y(n1409) );
  NAND2X1 U1017 ( .A(\mem<26><0> ), .B(n21), .Y(n1410) );
  OAI21X1 U1018 ( .A(n1230), .B(n1283), .C(n1410), .Y(n2284) );
  NAND2X1 U1019 ( .A(\mem<26><1> ), .B(n21), .Y(n1411) );
  OAI21X1 U1020 ( .A(n1230), .B(n1286), .C(n1411), .Y(n2283) );
  NAND2X1 U1021 ( .A(\mem<26><2> ), .B(n21), .Y(n1412) );
  OAI21X1 U1022 ( .A(n1230), .B(n1288), .C(n1412), .Y(n2282) );
  NAND2X1 U1023 ( .A(\mem<26><3> ), .B(n21), .Y(n1413) );
  OAI21X1 U1024 ( .A(n1230), .B(n1290), .C(n1413), .Y(n2281) );
  NAND2X1 U1025 ( .A(\mem<26><4> ), .B(n21), .Y(n1414) );
  OAI21X1 U1026 ( .A(n1230), .B(n1292), .C(n1414), .Y(n2280) );
  NAND2X1 U1027 ( .A(\mem<26><5> ), .B(n21), .Y(n1415) );
  OAI21X1 U1028 ( .A(n1230), .B(n1294), .C(n1415), .Y(n2279) );
  NAND2X1 U1029 ( .A(\mem<26><6> ), .B(n21), .Y(n1416) );
  OAI21X1 U1030 ( .A(n1230), .B(n1296), .C(n1416), .Y(n2278) );
  NAND2X1 U1031 ( .A(\mem<26><7> ), .B(n21), .Y(n1417) );
  OAI21X1 U1032 ( .A(n1230), .B(n1298), .C(n1417), .Y(n2277) );
  NAND2X1 U1033 ( .A(\mem<26><8> ), .B(n21), .Y(n1418) );
  OAI21X1 U1034 ( .A(n1231), .B(n1299), .C(n1418), .Y(n2276) );
  NAND2X1 U1035 ( .A(\mem<26><9> ), .B(n21), .Y(n1419) );
  OAI21X1 U1036 ( .A(n1231), .B(n1301), .C(n1419), .Y(n2275) );
  NAND2X1 U1037 ( .A(\mem<26><10> ), .B(n21), .Y(n1420) );
  OAI21X1 U1038 ( .A(n1231), .B(n1303), .C(n1420), .Y(n2274) );
  NAND2X1 U1039 ( .A(\mem<26><11> ), .B(n21), .Y(n1421) );
  OAI21X1 U1040 ( .A(n1231), .B(n1305), .C(n1421), .Y(n2273) );
  NAND2X1 U1041 ( .A(\mem<26><12> ), .B(n21), .Y(n1422) );
  OAI21X1 U1042 ( .A(n1231), .B(n1307), .C(n1422), .Y(n2272) );
  NAND2X1 U1043 ( .A(\mem<26><13> ), .B(n21), .Y(n1423) );
  OAI21X1 U1044 ( .A(n1231), .B(n1309), .C(n1423), .Y(n2271) );
  NAND2X1 U1045 ( .A(\mem<26><14> ), .B(n21), .Y(n1424) );
  OAI21X1 U1046 ( .A(n1231), .B(n1311), .C(n1424), .Y(n2270) );
  NAND2X1 U1047 ( .A(\mem<26><15> ), .B(n21), .Y(n1425) );
  OAI21X1 U1048 ( .A(n1231), .B(n1313), .C(n1425), .Y(n2269) );
  NAND3X1 U1049 ( .A(n1316), .B(n1321), .C(n1319), .Y(n1426) );
  NAND2X1 U1050 ( .A(\mem<25><0> ), .B(n23), .Y(n1427) );
  OAI21X1 U1051 ( .A(n1232), .B(n1283), .C(n1427), .Y(n2268) );
  NAND2X1 U1052 ( .A(\mem<25><1> ), .B(n23), .Y(n1428) );
  OAI21X1 U1053 ( .A(n1232), .B(n1285), .C(n1428), .Y(n2267) );
  NAND2X1 U1054 ( .A(\mem<25><2> ), .B(n23), .Y(n1429) );
  OAI21X1 U1055 ( .A(n1232), .B(n1287), .C(n1429), .Y(n2266) );
  NAND2X1 U1056 ( .A(\mem<25><3> ), .B(n23), .Y(n1430) );
  OAI21X1 U1057 ( .A(n1232), .B(n1289), .C(n1430), .Y(n2265) );
  NAND2X1 U1058 ( .A(\mem<25><4> ), .B(n23), .Y(n1431) );
  OAI21X1 U1059 ( .A(n1232), .B(n1291), .C(n1431), .Y(n2264) );
  NAND2X1 U1060 ( .A(\mem<25><5> ), .B(n23), .Y(n1432) );
  OAI21X1 U1061 ( .A(n1232), .B(n1293), .C(n1432), .Y(n2263) );
  NAND2X1 U1062 ( .A(\mem<25><6> ), .B(n23), .Y(n1433) );
  OAI21X1 U1063 ( .A(n1232), .B(n1295), .C(n1433), .Y(n2262) );
  NAND2X1 U1064 ( .A(\mem<25><7> ), .B(n23), .Y(n1434) );
  OAI21X1 U1065 ( .A(n1232), .B(n1297), .C(n1434), .Y(n2261) );
  NAND2X1 U1066 ( .A(\mem<25><8> ), .B(n23), .Y(n1435) );
  OAI21X1 U1067 ( .A(n1233), .B(n1300), .C(n1435), .Y(n2260) );
  NAND2X1 U1068 ( .A(\mem<25><9> ), .B(n23), .Y(n1436) );
  OAI21X1 U1069 ( .A(n1233), .B(n1302), .C(n1436), .Y(n2259) );
  NAND2X1 U1070 ( .A(\mem<25><10> ), .B(n23), .Y(n1437) );
  OAI21X1 U1071 ( .A(n1233), .B(n1304), .C(n1437), .Y(n2258) );
  NAND2X1 U1072 ( .A(\mem<25><11> ), .B(n23), .Y(n1438) );
  OAI21X1 U1073 ( .A(n1233), .B(n1306), .C(n1438), .Y(n2257) );
  NAND2X1 U1074 ( .A(\mem<25><12> ), .B(n23), .Y(n1439) );
  OAI21X1 U1075 ( .A(n1233), .B(n1308), .C(n1439), .Y(n2256) );
  NAND2X1 U1076 ( .A(\mem<25><13> ), .B(n23), .Y(n1440) );
  OAI21X1 U1077 ( .A(n1233), .B(n1310), .C(n1440), .Y(n2255) );
  NAND2X1 U1078 ( .A(\mem<25><14> ), .B(n23), .Y(n1441) );
  OAI21X1 U1079 ( .A(n1233), .B(n1312), .C(n1441), .Y(n2254) );
  NAND2X1 U1080 ( .A(\mem<25><15> ), .B(n23), .Y(n1442) );
  OAI21X1 U1081 ( .A(n1233), .B(n1314), .C(n1442), .Y(n2253) );
  NOR3X1 U1082 ( .A(n1316), .B(n1318), .C(n1320), .Y(n1836) );
  NAND2X1 U1083 ( .A(\mem<24><0> ), .B(n25), .Y(n1443) );
  OAI21X1 U1084 ( .A(n1234), .B(n1283), .C(n1443), .Y(n2252) );
  NAND2X1 U1085 ( .A(\mem<24><1> ), .B(n25), .Y(n1444) );
  OAI21X1 U1086 ( .A(n1234), .B(n1285), .C(n1444), .Y(n2251) );
  NAND2X1 U1087 ( .A(\mem<24><2> ), .B(n25), .Y(n1445) );
  OAI21X1 U1088 ( .A(n1234), .B(n1287), .C(n1445), .Y(n2250) );
  NAND2X1 U1089 ( .A(\mem<24><3> ), .B(n25), .Y(n1446) );
  OAI21X1 U1090 ( .A(n1234), .B(n1289), .C(n1446), .Y(n2249) );
  NAND2X1 U1091 ( .A(\mem<24><4> ), .B(n25), .Y(n1447) );
  OAI21X1 U1092 ( .A(n1234), .B(n1291), .C(n1447), .Y(n2248) );
  NAND2X1 U1093 ( .A(\mem<24><5> ), .B(n25), .Y(n1448) );
  OAI21X1 U1094 ( .A(n1234), .B(n1293), .C(n1448), .Y(n2247) );
  NAND2X1 U1095 ( .A(\mem<24><6> ), .B(n25), .Y(n1449) );
  OAI21X1 U1096 ( .A(n1234), .B(n1295), .C(n1449), .Y(n2246) );
  NAND2X1 U1097 ( .A(\mem<24><7> ), .B(n25), .Y(n1450) );
  OAI21X1 U1098 ( .A(n1234), .B(n1297), .C(n1450), .Y(n2245) );
  NAND2X1 U1099 ( .A(\mem<24><8> ), .B(n25), .Y(n1451) );
  OAI21X1 U1100 ( .A(n1234), .B(n1299), .C(n1451), .Y(n2244) );
  NAND2X1 U1101 ( .A(\mem<24><9> ), .B(n25), .Y(n1452) );
  OAI21X1 U1102 ( .A(n1234), .B(n1301), .C(n1452), .Y(n2243) );
  NAND2X1 U1103 ( .A(\mem<24><10> ), .B(n25), .Y(n1453) );
  OAI21X1 U1104 ( .A(n1234), .B(n1303), .C(n1453), .Y(n2242) );
  NAND2X1 U1105 ( .A(\mem<24><11> ), .B(n25), .Y(n1454) );
  OAI21X1 U1106 ( .A(n1234), .B(n1305), .C(n1454), .Y(n2241) );
  NAND2X1 U1107 ( .A(\mem<24><12> ), .B(n25), .Y(n1455) );
  OAI21X1 U1108 ( .A(n1234), .B(n1307), .C(n1455), .Y(n2240) );
  NAND2X1 U1109 ( .A(\mem<24><13> ), .B(n25), .Y(n1456) );
  OAI21X1 U1110 ( .A(n1234), .B(n1309), .C(n1456), .Y(n2239) );
  NAND2X1 U1111 ( .A(\mem<24><14> ), .B(n25), .Y(n1457) );
  OAI21X1 U1112 ( .A(n1234), .B(n1311), .C(n1457), .Y(n2238) );
  NAND2X1 U1113 ( .A(\mem<24><15> ), .B(n25), .Y(n1458) );
  OAI21X1 U1114 ( .A(n1234), .B(n1313), .C(n1458), .Y(n2237) );
  NAND2X1 U1115 ( .A(\mem<23><0> ), .B(n27), .Y(n1459) );
  OAI21X1 U1116 ( .A(n1235), .B(n1283), .C(n1459), .Y(n2236) );
  NAND2X1 U1117 ( .A(\mem<23><1> ), .B(n27), .Y(n1460) );
  OAI21X1 U1118 ( .A(n1235), .B(n1286), .C(n1460), .Y(n2235) );
  NAND2X1 U1119 ( .A(\mem<23><2> ), .B(n27), .Y(n1461) );
  OAI21X1 U1120 ( .A(n1235), .B(n1288), .C(n1461), .Y(n2234) );
  NAND2X1 U1121 ( .A(\mem<23><3> ), .B(n27), .Y(n1462) );
  OAI21X1 U1122 ( .A(n1235), .B(n1290), .C(n1462), .Y(n2233) );
  NAND2X1 U1123 ( .A(\mem<23><4> ), .B(n27), .Y(n1463) );
  OAI21X1 U1124 ( .A(n1235), .B(n1292), .C(n1463), .Y(n2232) );
  NAND2X1 U1125 ( .A(\mem<23><5> ), .B(n27), .Y(n1464) );
  OAI21X1 U1126 ( .A(n1235), .B(n1294), .C(n1464), .Y(n2231) );
  NAND2X1 U1127 ( .A(\mem<23><6> ), .B(n27), .Y(n1465) );
  OAI21X1 U1128 ( .A(n1235), .B(n1296), .C(n1465), .Y(n2230) );
  NAND2X1 U1129 ( .A(\mem<23><7> ), .B(n27), .Y(n1466) );
  OAI21X1 U1130 ( .A(n1235), .B(n1298), .C(n1466), .Y(n2229) );
  NAND2X1 U1131 ( .A(\mem<23><8> ), .B(n27), .Y(n1467) );
  OAI21X1 U1132 ( .A(n1236), .B(n1300), .C(n1467), .Y(n2228) );
  NAND2X1 U1133 ( .A(\mem<23><9> ), .B(n27), .Y(n1468) );
  OAI21X1 U1134 ( .A(n1236), .B(n1302), .C(n1468), .Y(n2227) );
  NAND2X1 U1135 ( .A(\mem<23><10> ), .B(n27), .Y(n1469) );
  OAI21X1 U1136 ( .A(n1236), .B(n1304), .C(n1469), .Y(n2226) );
  NAND2X1 U1137 ( .A(\mem<23><11> ), .B(n27), .Y(n1470) );
  OAI21X1 U1138 ( .A(n1236), .B(n1306), .C(n1470), .Y(n2225) );
  NAND2X1 U1139 ( .A(\mem<23><12> ), .B(n27), .Y(n1471) );
  OAI21X1 U1140 ( .A(n1236), .B(n1308), .C(n1471), .Y(n2224) );
  NAND2X1 U1141 ( .A(\mem<23><13> ), .B(n27), .Y(n1472) );
  OAI21X1 U1142 ( .A(n1236), .B(n1310), .C(n1472), .Y(n2223) );
  NAND2X1 U1143 ( .A(\mem<23><14> ), .B(n27), .Y(n1473) );
  OAI21X1 U1144 ( .A(n1236), .B(n1312), .C(n1473), .Y(n2222) );
  NAND2X1 U1145 ( .A(\mem<23><15> ), .B(n27), .Y(n1474) );
  OAI21X1 U1146 ( .A(n1236), .B(n1314), .C(n1474), .Y(n2221) );
  NAND2X1 U1147 ( .A(\mem<22><0> ), .B(n29), .Y(n1475) );
  OAI21X1 U1148 ( .A(n1237), .B(n1283), .C(n1475), .Y(n2220) );
  NAND2X1 U1149 ( .A(\mem<22><1> ), .B(n29), .Y(n1476) );
  OAI21X1 U1150 ( .A(n1237), .B(n1286), .C(n1476), .Y(n2219) );
  NAND2X1 U1151 ( .A(\mem<22><2> ), .B(n29), .Y(n1477) );
  OAI21X1 U1152 ( .A(n1237), .B(n1288), .C(n1477), .Y(n2218) );
  NAND2X1 U1153 ( .A(\mem<22><3> ), .B(n29), .Y(n1478) );
  OAI21X1 U1154 ( .A(n1237), .B(n1290), .C(n1478), .Y(n2217) );
  NAND2X1 U1155 ( .A(\mem<22><4> ), .B(n29), .Y(n1479) );
  OAI21X1 U1156 ( .A(n1237), .B(n1292), .C(n1479), .Y(n2216) );
  NAND2X1 U1157 ( .A(\mem<22><5> ), .B(n29), .Y(n1480) );
  OAI21X1 U1158 ( .A(n1237), .B(n1294), .C(n1480), .Y(n2215) );
  NAND2X1 U1159 ( .A(\mem<22><6> ), .B(n29), .Y(n1481) );
  OAI21X1 U1160 ( .A(n1237), .B(n1296), .C(n1481), .Y(n2214) );
  NAND2X1 U1161 ( .A(\mem<22><7> ), .B(n29), .Y(n1482) );
  OAI21X1 U1162 ( .A(n1237), .B(n1298), .C(n1482), .Y(n2213) );
  NAND2X1 U1163 ( .A(\mem<22><8> ), .B(n29), .Y(n1483) );
  OAI21X1 U1164 ( .A(n1238), .B(n1300), .C(n1483), .Y(n2212) );
  NAND2X1 U1165 ( .A(\mem<22><9> ), .B(n29), .Y(n1484) );
  OAI21X1 U1166 ( .A(n1238), .B(n1302), .C(n1484), .Y(n2211) );
  NAND2X1 U1167 ( .A(\mem<22><10> ), .B(n29), .Y(n1485) );
  OAI21X1 U1168 ( .A(n1238), .B(n1304), .C(n1485), .Y(n2210) );
  NAND2X1 U1169 ( .A(\mem<22><11> ), .B(n29), .Y(n1486) );
  OAI21X1 U1170 ( .A(n1238), .B(n1306), .C(n1486), .Y(n2209) );
  NAND2X1 U1171 ( .A(\mem<22><12> ), .B(n29), .Y(n1487) );
  OAI21X1 U1172 ( .A(n1238), .B(n1308), .C(n1487), .Y(n2208) );
  NAND2X1 U1173 ( .A(\mem<22><13> ), .B(n29), .Y(n1488) );
  OAI21X1 U1174 ( .A(n1238), .B(n1310), .C(n1488), .Y(n2207) );
  NAND2X1 U1175 ( .A(\mem<22><14> ), .B(n29), .Y(n1489) );
  OAI21X1 U1177 ( .A(n1238), .B(n1312), .C(n1489), .Y(n2206) );
  NAND2X1 U1178 ( .A(\mem<22><15> ), .B(n29), .Y(n1490) );
  OAI21X1 U1179 ( .A(n1238), .B(n1314), .C(n1490), .Y(n2205) );
  NAND2X1 U1180 ( .A(\mem<21><0> ), .B(n31), .Y(n1491) );
  OAI21X1 U1181 ( .A(n1239), .B(n1283), .C(n1491), .Y(n2204) );
  NAND2X1 U1182 ( .A(\mem<21><1> ), .B(n31), .Y(n1492) );
  OAI21X1 U1183 ( .A(n1239), .B(n1286), .C(n1492), .Y(n2203) );
  NAND2X1 U1184 ( .A(\mem<21><2> ), .B(n31), .Y(n1493) );
  OAI21X1 U1185 ( .A(n1239), .B(n1288), .C(n1493), .Y(n2202) );
  NAND2X1 U1186 ( .A(\mem<21><3> ), .B(n31), .Y(n1494) );
  OAI21X1 U1187 ( .A(n1239), .B(n1290), .C(n1494), .Y(n2201) );
  NAND2X1 U1188 ( .A(\mem<21><4> ), .B(n31), .Y(n1495) );
  OAI21X1 U1189 ( .A(n1239), .B(n1292), .C(n1495), .Y(n2200) );
  NAND2X1 U1190 ( .A(\mem<21><5> ), .B(n31), .Y(n1496) );
  OAI21X1 U1191 ( .A(n1239), .B(n1294), .C(n1496), .Y(n2199) );
  NAND2X1 U1192 ( .A(\mem<21><6> ), .B(n31), .Y(n1497) );
  OAI21X1 U1193 ( .A(n1239), .B(n1296), .C(n1497), .Y(n2198) );
  NAND2X1 U1194 ( .A(\mem<21><7> ), .B(n31), .Y(n1498) );
  OAI21X1 U1195 ( .A(n1239), .B(n1298), .C(n1498), .Y(n2197) );
  NAND2X1 U1196 ( .A(\mem<21><8> ), .B(n31), .Y(n1499) );
  OAI21X1 U1197 ( .A(n1240), .B(n1300), .C(n1499), .Y(n2196) );
  NAND2X1 U1198 ( .A(\mem<21><9> ), .B(n31), .Y(n1500) );
  OAI21X1 U1199 ( .A(n1240), .B(n1302), .C(n1500), .Y(n2195) );
  NAND2X1 U1200 ( .A(\mem<21><10> ), .B(n31), .Y(n1501) );
  OAI21X1 U1201 ( .A(n1240), .B(n1304), .C(n1501), .Y(n2194) );
  NAND2X1 U1202 ( .A(\mem<21><11> ), .B(n31), .Y(n1502) );
  OAI21X1 U1203 ( .A(n1240), .B(n1306), .C(n1502), .Y(n2193) );
  NAND2X1 U1204 ( .A(\mem<21><12> ), .B(n31), .Y(n1503) );
  OAI21X1 U1205 ( .A(n1240), .B(n1308), .C(n1503), .Y(n2192) );
  NAND2X1 U1206 ( .A(\mem<21><13> ), .B(n31), .Y(n1504) );
  OAI21X1 U1207 ( .A(n1240), .B(n1310), .C(n1504), .Y(n2191) );
  NAND2X1 U1208 ( .A(\mem<21><14> ), .B(n31), .Y(n1505) );
  OAI21X1 U1209 ( .A(n1240), .B(n1312), .C(n1505), .Y(n2190) );
  NAND2X1 U1210 ( .A(\mem<21><15> ), .B(n31), .Y(n1506) );
  OAI21X1 U1211 ( .A(n1240), .B(n1314), .C(n1506), .Y(n2189) );
  NAND2X1 U1212 ( .A(\mem<20><0> ), .B(n35), .Y(n1507) );
  OAI21X1 U1213 ( .A(n1241), .B(n1283), .C(n1507), .Y(n2188) );
  NAND2X1 U1214 ( .A(\mem<20><1> ), .B(n35), .Y(n1508) );
  OAI21X1 U1215 ( .A(n1241), .B(n1286), .C(n1508), .Y(n2187) );
  NAND2X1 U1216 ( .A(\mem<20><2> ), .B(n35), .Y(n1509) );
  OAI21X1 U1217 ( .A(n1241), .B(n1288), .C(n1509), .Y(n2186) );
  NAND2X1 U1218 ( .A(\mem<20><3> ), .B(n35), .Y(n1510) );
  OAI21X1 U1219 ( .A(n1241), .B(n1290), .C(n1510), .Y(n2185) );
  NAND2X1 U1220 ( .A(\mem<20><4> ), .B(n35), .Y(n1511) );
  OAI21X1 U1221 ( .A(n1241), .B(n1292), .C(n1511), .Y(n2184) );
  NAND2X1 U1222 ( .A(\mem<20><5> ), .B(n35), .Y(n1512) );
  OAI21X1 U1223 ( .A(n1241), .B(n1294), .C(n1512), .Y(n2183) );
  NAND2X1 U1224 ( .A(\mem<20><6> ), .B(n35), .Y(n1513) );
  OAI21X1 U1225 ( .A(n1241), .B(n1296), .C(n1513), .Y(n2182) );
  NAND2X1 U1226 ( .A(\mem<20><7> ), .B(n35), .Y(n1514) );
  OAI21X1 U1227 ( .A(n1241), .B(n1298), .C(n1514), .Y(n2181) );
  NAND2X1 U1228 ( .A(\mem<20><8> ), .B(n35), .Y(n1515) );
  OAI21X1 U1229 ( .A(n1242), .B(n1300), .C(n1515), .Y(n2180) );
  NAND2X1 U1230 ( .A(\mem<20><9> ), .B(n35), .Y(n1516) );
  OAI21X1 U1231 ( .A(n1242), .B(n1302), .C(n1516), .Y(n2179) );
  NAND2X1 U1232 ( .A(\mem<20><10> ), .B(n35), .Y(n1517) );
  OAI21X1 U1233 ( .A(n1242), .B(n1304), .C(n1517), .Y(n2178) );
  NAND2X1 U1234 ( .A(\mem<20><11> ), .B(n35), .Y(n1518) );
  OAI21X1 U1235 ( .A(n1242), .B(n1306), .C(n1518), .Y(n2177) );
  NAND2X1 U1236 ( .A(\mem<20><12> ), .B(n35), .Y(n1519) );
  OAI21X1 U1237 ( .A(n1242), .B(n1308), .C(n1519), .Y(n2176) );
  NAND2X1 U1238 ( .A(\mem<20><13> ), .B(n35), .Y(n1520) );
  OAI21X1 U1239 ( .A(n1242), .B(n1310), .C(n1520), .Y(n2175) );
  NAND2X1 U1240 ( .A(\mem<20><14> ), .B(n35), .Y(n1521) );
  OAI21X1 U1241 ( .A(n1242), .B(n1312), .C(n1521), .Y(n2174) );
  NAND2X1 U1242 ( .A(\mem<20><15> ), .B(n35), .Y(n1522) );
  OAI21X1 U1243 ( .A(n1242), .B(n1314), .C(n1522), .Y(n2173) );
  NAND2X1 U1244 ( .A(\mem<19><0> ), .B(n45), .Y(n1523) );
  OAI21X1 U1245 ( .A(n1243), .B(n1284), .C(n1523), .Y(n2172) );
  NAND2X1 U1246 ( .A(\mem<19><1> ), .B(n45), .Y(n1524) );
  OAI21X1 U1247 ( .A(n1243), .B(n1286), .C(n1524), .Y(n2171) );
  NAND2X1 U1248 ( .A(\mem<19><2> ), .B(n45), .Y(n1525) );
  OAI21X1 U1249 ( .A(n1243), .B(n1288), .C(n1525), .Y(n2170) );
  NAND2X1 U1250 ( .A(\mem<19><3> ), .B(n45), .Y(n1526) );
  OAI21X1 U1251 ( .A(n1243), .B(n1290), .C(n1526), .Y(n2169) );
  NAND2X1 U1252 ( .A(\mem<19><4> ), .B(n45), .Y(n1527) );
  OAI21X1 U1253 ( .A(n1243), .B(n1292), .C(n1527), .Y(n2168) );
  NAND2X1 U1254 ( .A(\mem<19><5> ), .B(n45), .Y(n1528) );
  OAI21X1 U1255 ( .A(n1243), .B(n1294), .C(n1528), .Y(n2167) );
  NAND2X1 U1256 ( .A(\mem<19><6> ), .B(n45), .Y(n1529) );
  OAI21X1 U1257 ( .A(n1243), .B(n1296), .C(n1529), .Y(n2166) );
  NAND2X1 U1258 ( .A(\mem<19><7> ), .B(n45), .Y(n1530) );
  OAI21X1 U1259 ( .A(n1243), .B(n1298), .C(n1530), .Y(n2165) );
  NAND2X1 U1260 ( .A(\mem<19><8> ), .B(n45), .Y(n1531) );
  OAI21X1 U1261 ( .A(n1244), .B(n1300), .C(n1531), .Y(n2164) );
  NAND2X1 U1262 ( .A(\mem<19><9> ), .B(n45), .Y(n1532) );
  OAI21X1 U1263 ( .A(n1244), .B(n1302), .C(n1532), .Y(n2163) );
  NAND2X1 U1264 ( .A(\mem<19><10> ), .B(n45), .Y(n1533) );
  OAI21X1 U1265 ( .A(n1244), .B(n1304), .C(n1533), .Y(n2162) );
  NAND2X1 U1266 ( .A(\mem<19><11> ), .B(n45), .Y(n1534) );
  OAI21X1 U1267 ( .A(n1244), .B(n1306), .C(n1534), .Y(n2161) );
  NAND2X1 U1268 ( .A(\mem<19><12> ), .B(n45), .Y(n1535) );
  OAI21X1 U1269 ( .A(n1244), .B(n1308), .C(n1535), .Y(n2160) );
  NAND2X1 U1270 ( .A(\mem<19><13> ), .B(n45), .Y(n1536) );
  OAI21X1 U1271 ( .A(n1244), .B(n1310), .C(n1536), .Y(n2159) );
  NAND2X1 U1272 ( .A(\mem<19><14> ), .B(n45), .Y(n1537) );
  OAI21X1 U1273 ( .A(n1244), .B(n1312), .C(n1537), .Y(n2158) );
  NAND2X1 U1274 ( .A(\mem<19><15> ), .B(n45), .Y(n1538) );
  OAI21X1 U1275 ( .A(n1244), .B(n1314), .C(n1538), .Y(n2157) );
  NAND2X1 U1276 ( .A(\mem<18><0> ), .B(n47), .Y(n1539) );
  OAI21X1 U1277 ( .A(n1245), .B(n1284), .C(n1539), .Y(n2156) );
  NAND2X1 U1278 ( .A(\mem<18><1> ), .B(n47), .Y(n1540) );
  OAI21X1 U1279 ( .A(n1245), .B(n1286), .C(n1540), .Y(n2155) );
  NAND2X1 U1280 ( .A(\mem<18><2> ), .B(n47), .Y(n1541) );
  OAI21X1 U1281 ( .A(n1245), .B(n1288), .C(n1541), .Y(n2154) );
  NAND2X1 U1282 ( .A(\mem<18><3> ), .B(n47), .Y(n1542) );
  OAI21X1 U1283 ( .A(n1245), .B(n1290), .C(n1542), .Y(n2153) );
  NAND2X1 U1284 ( .A(\mem<18><4> ), .B(n47), .Y(n1543) );
  OAI21X1 U1285 ( .A(n1245), .B(n1292), .C(n1543), .Y(n2152) );
  NAND2X1 U1286 ( .A(\mem<18><5> ), .B(n47), .Y(n1544) );
  OAI21X1 U1287 ( .A(n1245), .B(n1294), .C(n1544), .Y(n2151) );
  NAND2X1 U1288 ( .A(\mem<18><6> ), .B(n47), .Y(n1545) );
  OAI21X1 U1289 ( .A(n1245), .B(n1296), .C(n1545), .Y(n2150) );
  NAND2X1 U1290 ( .A(\mem<18><7> ), .B(n47), .Y(n1546) );
  OAI21X1 U1291 ( .A(n1245), .B(n1298), .C(n1546), .Y(n2149) );
  NAND2X1 U1292 ( .A(\mem<18><8> ), .B(n47), .Y(n1547) );
  OAI21X1 U1293 ( .A(n1246), .B(n1300), .C(n1547), .Y(n2148) );
  NAND2X1 U1294 ( .A(\mem<18><9> ), .B(n47), .Y(n1548) );
  OAI21X1 U1295 ( .A(n1246), .B(n1302), .C(n1548), .Y(n2147) );
  NAND2X1 U1296 ( .A(\mem<18><10> ), .B(n47), .Y(n1549) );
  OAI21X1 U1297 ( .A(n1246), .B(n1304), .C(n1549), .Y(n2146) );
  NAND2X1 U1298 ( .A(\mem<18><11> ), .B(n47), .Y(n1550) );
  OAI21X1 U1299 ( .A(n1246), .B(n1306), .C(n1550), .Y(n2145) );
  NAND2X1 U1300 ( .A(\mem<18><12> ), .B(n47), .Y(n1551) );
  OAI21X1 U1301 ( .A(n1246), .B(n1308), .C(n1551), .Y(n2144) );
  NAND2X1 U1302 ( .A(\mem<18><13> ), .B(n47), .Y(n1552) );
  OAI21X1 U1303 ( .A(n1246), .B(n1310), .C(n1552), .Y(n2143) );
  NAND2X1 U1304 ( .A(\mem<18><14> ), .B(n47), .Y(n1553) );
  OAI21X1 U1305 ( .A(n1246), .B(n1312), .C(n1553), .Y(n2142) );
  NAND2X1 U1306 ( .A(\mem<18><15> ), .B(n47), .Y(n1554) );
  OAI21X1 U1307 ( .A(n1246), .B(n1314), .C(n1554), .Y(n2141) );
  NAND2X1 U1308 ( .A(\mem<17><0> ), .B(n49), .Y(n1555) );
  OAI21X1 U1309 ( .A(n1247), .B(n1284), .C(n1555), .Y(n2140) );
  NAND2X1 U1310 ( .A(\mem<17><1> ), .B(n49), .Y(n1556) );
  OAI21X1 U1311 ( .A(n1247), .B(n1286), .C(n1556), .Y(n2139) );
  NAND2X1 U1312 ( .A(\mem<17><2> ), .B(n49), .Y(n1557) );
  OAI21X1 U1313 ( .A(n1247), .B(n1288), .C(n1557), .Y(n2138) );
  NAND2X1 U1314 ( .A(\mem<17><3> ), .B(n49), .Y(n1558) );
  OAI21X1 U1315 ( .A(n1247), .B(n1290), .C(n1558), .Y(n2137) );
  NAND2X1 U1316 ( .A(\mem<17><4> ), .B(n49), .Y(n1559) );
  OAI21X1 U1317 ( .A(n1247), .B(n1292), .C(n1559), .Y(n2136) );
  NAND2X1 U1318 ( .A(\mem<17><5> ), .B(n49), .Y(n1560) );
  OAI21X1 U1319 ( .A(n1247), .B(n1294), .C(n1560), .Y(n2135) );
  NAND2X1 U1320 ( .A(\mem<17><6> ), .B(n49), .Y(n1561) );
  OAI21X1 U1321 ( .A(n1247), .B(n1296), .C(n1561), .Y(n2134) );
  NAND2X1 U1322 ( .A(\mem<17><7> ), .B(n49), .Y(n1562) );
  OAI21X1 U1323 ( .A(n1247), .B(n1298), .C(n1562), .Y(n2133) );
  NAND2X1 U1324 ( .A(\mem<17><8> ), .B(n49), .Y(n1563) );
  OAI21X1 U1325 ( .A(n1248), .B(n1300), .C(n1563), .Y(n2132) );
  NAND2X1 U1326 ( .A(\mem<17><9> ), .B(n49), .Y(n1564) );
  OAI21X1 U1327 ( .A(n1248), .B(n1302), .C(n1564), .Y(n2131) );
  NAND2X1 U1328 ( .A(\mem<17><10> ), .B(n49), .Y(n1565) );
  OAI21X1 U1329 ( .A(n1248), .B(n1304), .C(n1565), .Y(n2130) );
  NAND2X1 U1330 ( .A(\mem<17><11> ), .B(n49), .Y(n1566) );
  OAI21X1 U1331 ( .A(n1248), .B(n1306), .C(n1566), .Y(n2129) );
  NAND2X1 U1332 ( .A(\mem<17><12> ), .B(n49), .Y(n1567) );
  OAI21X1 U1333 ( .A(n1248), .B(n1308), .C(n1567), .Y(n2128) );
  NAND2X1 U1334 ( .A(\mem<17><13> ), .B(n49), .Y(n1568) );
  OAI21X1 U1335 ( .A(n1248), .B(n1310), .C(n1568), .Y(n2127) );
  NAND2X1 U1336 ( .A(\mem<17><14> ), .B(n49), .Y(n1569) );
  OAI21X1 U1337 ( .A(n1248), .B(n1312), .C(n1569), .Y(n2126) );
  NAND2X1 U1338 ( .A(\mem<17><15> ), .B(n49), .Y(n1570) );
  OAI21X1 U1339 ( .A(n1248), .B(n1314), .C(n1570), .Y(n2125) );
  NAND2X1 U1340 ( .A(\mem<16><0> ), .B(n82), .Y(n1571) );
  OAI21X1 U1341 ( .A(n1249), .B(n1284), .C(n1571), .Y(n2124) );
  NAND2X1 U1342 ( .A(\mem<16><1> ), .B(n82), .Y(n1572) );
  OAI21X1 U1343 ( .A(n1249), .B(n1286), .C(n1572), .Y(n2123) );
  NAND2X1 U1344 ( .A(\mem<16><2> ), .B(n82), .Y(n1573) );
  OAI21X1 U1345 ( .A(n1249), .B(n1288), .C(n1573), .Y(n2122) );
  NAND2X1 U1346 ( .A(\mem<16><3> ), .B(n82), .Y(n1574) );
  OAI21X1 U1347 ( .A(n1249), .B(n1290), .C(n1574), .Y(n2121) );
  NAND2X1 U1348 ( .A(\mem<16><4> ), .B(n82), .Y(n1575) );
  OAI21X1 U1349 ( .A(n1249), .B(n1292), .C(n1575), .Y(n2120) );
  NAND2X1 U1350 ( .A(\mem<16><5> ), .B(n82), .Y(n1576) );
  OAI21X1 U1351 ( .A(n1249), .B(n1294), .C(n1576), .Y(n2119) );
  NAND2X1 U1352 ( .A(\mem<16><6> ), .B(n82), .Y(n1577) );
  OAI21X1 U1353 ( .A(n1249), .B(n1296), .C(n1577), .Y(n2118) );
  NAND2X1 U1354 ( .A(\mem<16><7> ), .B(n82), .Y(n1578) );
  OAI21X1 U1355 ( .A(n1249), .B(n1298), .C(n1578), .Y(n2117) );
  NAND2X1 U1356 ( .A(\mem<16><8> ), .B(n82), .Y(n1579) );
  OAI21X1 U1357 ( .A(n1249), .B(n1300), .C(n1579), .Y(n2116) );
  NAND2X1 U1358 ( .A(\mem<16><9> ), .B(n82), .Y(n1580) );
  OAI21X1 U1359 ( .A(n1249), .B(n1302), .C(n1580), .Y(n2115) );
  NAND2X1 U1360 ( .A(\mem<16><10> ), .B(n82), .Y(n1581) );
  OAI21X1 U1361 ( .A(n1249), .B(n1304), .C(n1581), .Y(n2114) );
  NAND2X1 U1362 ( .A(\mem<16><11> ), .B(n82), .Y(n1582) );
  OAI21X1 U1363 ( .A(n1249), .B(n1306), .C(n1582), .Y(n2113) );
  NAND2X1 U1364 ( .A(\mem<16><12> ), .B(n82), .Y(n1583) );
  OAI21X1 U1365 ( .A(n1249), .B(n1308), .C(n1583), .Y(n2112) );
  NAND2X1 U1366 ( .A(\mem<16><13> ), .B(n82), .Y(n1584) );
  OAI21X1 U1367 ( .A(n1249), .B(n1310), .C(n1584), .Y(n2111) );
  NAND2X1 U1368 ( .A(\mem<16><14> ), .B(n82), .Y(n1585) );
  OAI21X1 U1369 ( .A(n1249), .B(n1312), .C(n1585), .Y(n2110) );
  NAND2X1 U1370 ( .A(\mem<16><15> ), .B(n82), .Y(n1586) );
  OAI21X1 U1371 ( .A(n1249), .B(n1314), .C(n1586), .Y(n2109) );
  NAND3X1 U1372 ( .A(n1322), .B(n2365), .C(n1325), .Y(n1587) );
  NAND2X1 U1373 ( .A(\mem<15><0> ), .B(n51), .Y(n1588) );
  OAI21X1 U1374 ( .A(n1250), .B(n1284), .C(n1588), .Y(n2108) );
  NAND2X1 U1375 ( .A(\mem<15><1> ), .B(n51), .Y(n1589) );
  OAI21X1 U1376 ( .A(n1250), .B(n1286), .C(n1589), .Y(n2107) );
  NAND2X1 U1377 ( .A(\mem<15><2> ), .B(n51), .Y(n1590) );
  OAI21X1 U1378 ( .A(n1250), .B(n1288), .C(n1590), .Y(n2106) );
  NAND2X1 U1379 ( .A(\mem<15><3> ), .B(n51), .Y(n1591) );
  OAI21X1 U1380 ( .A(n1250), .B(n1290), .C(n1591), .Y(n2105) );
  NAND2X1 U1381 ( .A(\mem<15><4> ), .B(n51), .Y(n1592) );
  OAI21X1 U1382 ( .A(n1250), .B(n1292), .C(n1592), .Y(n2104) );
  NAND2X1 U1383 ( .A(\mem<15><5> ), .B(n51), .Y(n1593) );
  OAI21X1 U1384 ( .A(n1250), .B(n1294), .C(n1593), .Y(n2103) );
  NAND2X1 U1385 ( .A(\mem<15><6> ), .B(n51), .Y(n1594) );
  OAI21X1 U1386 ( .A(n1250), .B(n1296), .C(n1594), .Y(n2102) );
  NAND2X1 U1387 ( .A(\mem<15><7> ), .B(n51), .Y(n1595) );
  OAI21X1 U1388 ( .A(n1250), .B(n1298), .C(n1595), .Y(n2101) );
  NAND2X1 U1389 ( .A(\mem<15><8> ), .B(n51), .Y(n1596) );
  OAI21X1 U1390 ( .A(n1251), .B(n1300), .C(n1596), .Y(n2100) );
  NAND2X1 U1391 ( .A(\mem<15><9> ), .B(n51), .Y(n1597) );
  OAI21X1 U1392 ( .A(n1251), .B(n1302), .C(n1597), .Y(n2099) );
  NAND2X1 U1393 ( .A(\mem<15><10> ), .B(n51), .Y(n1598) );
  OAI21X1 U1394 ( .A(n1251), .B(n1304), .C(n1598), .Y(n2098) );
  NAND2X1 U1395 ( .A(\mem<15><11> ), .B(n51), .Y(n1599) );
  OAI21X1 U1396 ( .A(n1251), .B(n1306), .C(n1599), .Y(n2097) );
  NAND2X1 U1397 ( .A(\mem<15><12> ), .B(n51), .Y(n1600) );
  OAI21X1 U1398 ( .A(n1251), .B(n1308), .C(n1600), .Y(n2096) );
  NAND2X1 U1399 ( .A(\mem<15><13> ), .B(n51), .Y(n1601) );
  OAI21X1 U1400 ( .A(n1251), .B(n1310), .C(n1601), .Y(n2095) );
  NAND2X1 U1401 ( .A(\mem<15><14> ), .B(n51), .Y(n1602) );
  OAI21X1 U1402 ( .A(n1251), .B(n1312), .C(n1602), .Y(n2094) );
  NAND2X1 U1403 ( .A(\mem<15><15> ), .B(n51), .Y(n1603) );
  OAI21X1 U1404 ( .A(n1251), .B(n1314), .C(n1603), .Y(n2093) );
  NAND2X1 U1405 ( .A(\mem<14><0> ), .B(n53), .Y(n1604) );
  OAI21X1 U1406 ( .A(n1252), .B(n1284), .C(n1604), .Y(n2092) );
  NAND2X1 U1407 ( .A(\mem<14><1> ), .B(n53), .Y(n1605) );
  OAI21X1 U1408 ( .A(n1252), .B(n1286), .C(n1605), .Y(n2091) );
  NAND2X1 U1409 ( .A(\mem<14><2> ), .B(n53), .Y(n1606) );
  OAI21X1 U1410 ( .A(n1252), .B(n1288), .C(n1606), .Y(n2090) );
  NAND2X1 U1411 ( .A(\mem<14><3> ), .B(n53), .Y(n1607) );
  OAI21X1 U1412 ( .A(n1252), .B(n1290), .C(n1607), .Y(n2089) );
  NAND2X1 U1413 ( .A(\mem<14><4> ), .B(n53), .Y(n1608) );
  OAI21X1 U1414 ( .A(n1252), .B(n1292), .C(n1608), .Y(n2088) );
  NAND2X1 U1415 ( .A(\mem<14><5> ), .B(n53), .Y(n1609) );
  OAI21X1 U1416 ( .A(n1252), .B(n1294), .C(n1609), .Y(n2087) );
  NAND2X1 U1417 ( .A(\mem<14><6> ), .B(n53), .Y(n1610) );
  OAI21X1 U1418 ( .A(n1252), .B(n1296), .C(n1610), .Y(n2086) );
  NAND2X1 U1419 ( .A(\mem<14><7> ), .B(n53), .Y(n1611) );
  OAI21X1 U1420 ( .A(n1252), .B(n1298), .C(n1611), .Y(n2085) );
  NAND2X1 U1421 ( .A(\mem<14><8> ), .B(n53), .Y(n1612) );
  OAI21X1 U1422 ( .A(n1253), .B(n1300), .C(n1612), .Y(n2084) );
  NAND2X1 U1423 ( .A(\mem<14><9> ), .B(n53), .Y(n1613) );
  OAI21X1 U1424 ( .A(n1253), .B(n1302), .C(n1613), .Y(n2083) );
  NAND2X1 U1425 ( .A(\mem<14><10> ), .B(n53), .Y(n1614) );
  OAI21X1 U1426 ( .A(n1253), .B(n1304), .C(n1614), .Y(n2082) );
  NAND2X1 U1427 ( .A(\mem<14><11> ), .B(n53), .Y(n1615) );
  OAI21X1 U1428 ( .A(n1253), .B(n1306), .C(n1615), .Y(n2081) );
  NAND2X1 U1429 ( .A(\mem<14><12> ), .B(n53), .Y(n1616) );
  OAI21X1 U1430 ( .A(n1253), .B(n1308), .C(n1616), .Y(n2080) );
  NAND2X1 U1431 ( .A(\mem<14><13> ), .B(n53), .Y(n1617) );
  OAI21X1 U1432 ( .A(n1253), .B(n1310), .C(n1617), .Y(n2079) );
  NAND2X1 U1433 ( .A(\mem<14><14> ), .B(n53), .Y(n1618) );
  OAI21X1 U1434 ( .A(n1253), .B(n1312), .C(n1618), .Y(n2078) );
  NAND2X1 U1435 ( .A(\mem<14><15> ), .B(n53), .Y(n1619) );
  OAI21X1 U1436 ( .A(n1253), .B(n1314), .C(n1619), .Y(n2077) );
  NAND2X1 U1437 ( .A(\mem<13><0> ), .B(n55), .Y(n1620) );
  OAI21X1 U1438 ( .A(n1254), .B(n1284), .C(n1620), .Y(n2076) );
  NAND2X1 U1439 ( .A(\mem<13><1> ), .B(n55), .Y(n1621) );
  OAI21X1 U1440 ( .A(n1254), .B(n1286), .C(n1621), .Y(n2075) );
  NAND2X1 U1441 ( .A(\mem<13><2> ), .B(n55), .Y(n1622) );
  OAI21X1 U1442 ( .A(n1254), .B(n1288), .C(n1622), .Y(n2074) );
  NAND2X1 U1443 ( .A(\mem<13><3> ), .B(n55), .Y(n1623) );
  OAI21X1 U1444 ( .A(n1254), .B(n1290), .C(n1623), .Y(n2073) );
  NAND2X1 U1445 ( .A(\mem<13><4> ), .B(n55), .Y(n1624) );
  OAI21X1 U1446 ( .A(n1254), .B(n1292), .C(n1624), .Y(n2072) );
  NAND2X1 U1447 ( .A(\mem<13><5> ), .B(n55), .Y(n1625) );
  OAI21X1 U1448 ( .A(n1254), .B(n1294), .C(n1625), .Y(n2071) );
  NAND2X1 U1449 ( .A(\mem<13><6> ), .B(n55), .Y(n1626) );
  OAI21X1 U1450 ( .A(n1254), .B(n1296), .C(n1626), .Y(n2070) );
  NAND2X1 U1451 ( .A(\mem<13><7> ), .B(n55), .Y(n1627) );
  OAI21X1 U1452 ( .A(n1254), .B(n1298), .C(n1627), .Y(n2069) );
  NAND2X1 U1453 ( .A(\mem<13><8> ), .B(n55), .Y(n1628) );
  OAI21X1 U1454 ( .A(n1255), .B(n1300), .C(n1628), .Y(n2068) );
  NAND2X1 U1455 ( .A(\mem<13><9> ), .B(n55), .Y(n1629) );
  OAI21X1 U1456 ( .A(n1255), .B(n1302), .C(n1629), .Y(n2067) );
  NAND2X1 U1457 ( .A(\mem<13><10> ), .B(n55), .Y(n1630) );
  OAI21X1 U1458 ( .A(n1255), .B(n1304), .C(n1630), .Y(n2066) );
  NAND2X1 U1459 ( .A(\mem<13><11> ), .B(n55), .Y(n1631) );
  OAI21X1 U1460 ( .A(n1255), .B(n1306), .C(n1631), .Y(n2065) );
  NAND2X1 U1461 ( .A(\mem<13><12> ), .B(n55), .Y(n1632) );
  OAI21X1 U1462 ( .A(n1255), .B(n1308), .C(n1632), .Y(n2064) );
  NAND2X1 U1463 ( .A(\mem<13><13> ), .B(n55), .Y(n1633) );
  OAI21X1 U1464 ( .A(n1255), .B(n1310), .C(n1633), .Y(n2063) );
  NAND2X1 U1465 ( .A(\mem<13><14> ), .B(n55), .Y(n1634) );
  OAI21X1 U1466 ( .A(n1255), .B(n1312), .C(n1634), .Y(n2062) );
  NAND2X1 U1467 ( .A(\mem<13><15> ), .B(n55), .Y(n1635) );
  OAI21X1 U1468 ( .A(n1255), .B(n1314), .C(n1635), .Y(n2061) );
  NAND2X1 U1469 ( .A(\mem<12><0> ), .B(n57), .Y(n1636) );
  OAI21X1 U1470 ( .A(n1256), .B(n1284), .C(n1636), .Y(n2060) );
  NAND2X1 U1471 ( .A(\mem<12><1> ), .B(n57), .Y(n1637) );
  OAI21X1 U1472 ( .A(n1256), .B(n1286), .C(n1637), .Y(n2059) );
  NAND2X1 U1473 ( .A(\mem<12><2> ), .B(n57), .Y(n1638) );
  OAI21X1 U1474 ( .A(n1256), .B(n1288), .C(n1638), .Y(n2058) );
  NAND2X1 U1475 ( .A(\mem<12><3> ), .B(n57), .Y(n1639) );
  OAI21X1 U1476 ( .A(n1256), .B(n1290), .C(n1639), .Y(n2057) );
  NAND2X1 U1477 ( .A(\mem<12><4> ), .B(n57), .Y(n1640) );
  OAI21X1 U1478 ( .A(n1256), .B(n1292), .C(n1640), .Y(n2056) );
  NAND2X1 U1479 ( .A(\mem<12><5> ), .B(n57), .Y(n1641) );
  OAI21X1 U1480 ( .A(n1256), .B(n1294), .C(n1641), .Y(n2055) );
  NAND2X1 U1481 ( .A(\mem<12><6> ), .B(n57), .Y(n1642) );
  OAI21X1 U1482 ( .A(n1256), .B(n1296), .C(n1642), .Y(n2054) );
  NAND2X1 U1483 ( .A(\mem<12><7> ), .B(n57), .Y(n1643) );
  OAI21X1 U1484 ( .A(n1256), .B(n1298), .C(n1643), .Y(n2053) );
  NAND2X1 U1485 ( .A(\mem<12><8> ), .B(n57), .Y(n1644) );
  OAI21X1 U1486 ( .A(n1257), .B(n1300), .C(n1644), .Y(n2052) );
  NAND2X1 U1487 ( .A(\mem<12><9> ), .B(n57), .Y(n1645) );
  OAI21X1 U1488 ( .A(n1257), .B(n1302), .C(n1645), .Y(n2051) );
  NAND2X1 U1489 ( .A(\mem<12><10> ), .B(n57), .Y(n1646) );
  OAI21X1 U1490 ( .A(n1257), .B(n1304), .C(n1646), .Y(n2050) );
  NAND2X1 U1491 ( .A(\mem<12><11> ), .B(n57), .Y(n1647) );
  OAI21X1 U1492 ( .A(n1257), .B(n1306), .C(n1647), .Y(n2049) );
  NAND2X1 U1493 ( .A(\mem<12><12> ), .B(n57), .Y(n1648) );
  OAI21X1 U1494 ( .A(n1257), .B(n1308), .C(n1648), .Y(n2048) );
  NAND2X1 U1495 ( .A(\mem<12><13> ), .B(n57), .Y(n1649) );
  OAI21X1 U1496 ( .A(n1257), .B(n1310), .C(n1649), .Y(n2047) );
  NAND2X1 U1497 ( .A(\mem<12><14> ), .B(n57), .Y(n1650) );
  OAI21X1 U1498 ( .A(n1257), .B(n1312), .C(n1650), .Y(n2046) );
  NAND2X1 U1499 ( .A(\mem<12><15> ), .B(n57), .Y(n1651) );
  OAI21X1 U1500 ( .A(n1257), .B(n1314), .C(n1651), .Y(n2045) );
  NAND2X1 U1501 ( .A(\mem<11><0> ), .B(n59), .Y(n1652) );
  OAI21X1 U1502 ( .A(n1258), .B(n1284), .C(n1652), .Y(n2044) );
  NAND2X1 U1503 ( .A(\mem<11><1> ), .B(n59), .Y(n1653) );
  OAI21X1 U1504 ( .A(n1258), .B(n1285), .C(n1653), .Y(n2043) );
  NAND2X1 U1505 ( .A(\mem<11><2> ), .B(n59), .Y(n1654) );
  OAI21X1 U1506 ( .A(n1258), .B(n1287), .C(n1654), .Y(n2042) );
  NAND2X1 U1507 ( .A(\mem<11><3> ), .B(n59), .Y(n1655) );
  OAI21X1 U1508 ( .A(n1258), .B(n1289), .C(n1655), .Y(n2041) );
  NAND2X1 U1509 ( .A(\mem<11><4> ), .B(n59), .Y(n1656) );
  OAI21X1 U1510 ( .A(n1258), .B(n1291), .C(n1656), .Y(n2040) );
  NAND2X1 U1511 ( .A(\mem<11><5> ), .B(n59), .Y(n1657) );
  OAI21X1 U1512 ( .A(n1258), .B(n1293), .C(n1657), .Y(n2039) );
  NAND2X1 U1513 ( .A(\mem<11><6> ), .B(n59), .Y(n1658) );
  OAI21X1 U1514 ( .A(n1258), .B(n1295), .C(n1658), .Y(n2038) );
  NAND2X1 U1515 ( .A(\mem<11><7> ), .B(n59), .Y(n1659) );
  OAI21X1 U1516 ( .A(n1258), .B(n1297), .C(n1659), .Y(n2037) );
  NAND2X1 U1517 ( .A(\mem<11><8> ), .B(n59), .Y(n1660) );
  OAI21X1 U1518 ( .A(n1259), .B(n1299), .C(n1660), .Y(n2036) );
  NAND2X1 U1519 ( .A(\mem<11><9> ), .B(n59), .Y(n1661) );
  OAI21X1 U1520 ( .A(n1259), .B(n1301), .C(n1661), .Y(n2035) );
  NAND2X1 U1521 ( .A(\mem<11><10> ), .B(n59), .Y(n1662) );
  OAI21X1 U1522 ( .A(n1259), .B(n1303), .C(n1662), .Y(n2034) );
  NAND2X1 U1523 ( .A(\mem<11><11> ), .B(n59), .Y(n1663) );
  OAI21X1 U1524 ( .A(n1259), .B(n1305), .C(n1663), .Y(n2033) );
  NAND2X1 U1525 ( .A(\mem<11><12> ), .B(n59), .Y(n1664) );
  OAI21X1 U1526 ( .A(n1259), .B(n1307), .C(n1664), .Y(n2032) );
  NAND2X1 U1527 ( .A(\mem<11><13> ), .B(n59), .Y(n1665) );
  OAI21X1 U1528 ( .A(n1259), .B(n1309), .C(n1665), .Y(n2031) );
  NAND2X1 U1529 ( .A(\mem<11><14> ), .B(n59), .Y(n1666) );
  OAI21X1 U1530 ( .A(n1259), .B(n1311), .C(n1666), .Y(n2030) );
  NAND2X1 U1531 ( .A(\mem<11><15> ), .B(n59), .Y(n1667) );
  OAI21X1 U1532 ( .A(n1259), .B(n1313), .C(n1667), .Y(n2029) );
  NAND2X1 U1533 ( .A(\mem<10><0> ), .B(n61), .Y(n1668) );
  OAI21X1 U1534 ( .A(n1260), .B(n1284), .C(n1668), .Y(n2028) );
  NAND2X1 U1535 ( .A(\mem<10><1> ), .B(n61), .Y(n1669) );
  OAI21X1 U1536 ( .A(n1260), .B(n1285), .C(n1669), .Y(n2027) );
  NAND2X1 U1537 ( .A(\mem<10><2> ), .B(n61), .Y(n1670) );
  OAI21X1 U1538 ( .A(n1260), .B(n1287), .C(n1670), .Y(n2026) );
  NAND2X1 U1539 ( .A(\mem<10><3> ), .B(n61), .Y(n1671) );
  OAI21X1 U1540 ( .A(n1260), .B(n1289), .C(n1671), .Y(n2025) );
  NAND2X1 U1541 ( .A(\mem<10><4> ), .B(n61), .Y(n1672) );
  OAI21X1 U1542 ( .A(n1260), .B(n1291), .C(n1672), .Y(n2024) );
  NAND2X1 U1543 ( .A(\mem<10><5> ), .B(n61), .Y(n1673) );
  OAI21X1 U1544 ( .A(n1260), .B(n1293), .C(n1673), .Y(n2023) );
  NAND2X1 U1545 ( .A(\mem<10><6> ), .B(n61), .Y(n1674) );
  OAI21X1 U1546 ( .A(n1260), .B(n1295), .C(n1674), .Y(n2022) );
  NAND2X1 U1547 ( .A(\mem<10><7> ), .B(n61), .Y(n1675) );
  OAI21X1 U1548 ( .A(n1260), .B(n1297), .C(n1675), .Y(n2021) );
  NAND2X1 U1549 ( .A(\mem<10><8> ), .B(n61), .Y(n1676) );
  OAI21X1 U1550 ( .A(n1261), .B(n1299), .C(n1676), .Y(n2020) );
  NAND2X1 U1551 ( .A(\mem<10><9> ), .B(n61), .Y(n1677) );
  OAI21X1 U1552 ( .A(n1261), .B(n1301), .C(n1677), .Y(n2019) );
  NAND2X1 U1553 ( .A(\mem<10><10> ), .B(n61), .Y(n1678) );
  OAI21X1 U1554 ( .A(n1261), .B(n1303), .C(n1678), .Y(n2018) );
  NAND2X1 U1555 ( .A(\mem<10><11> ), .B(n61), .Y(n1679) );
  OAI21X1 U1556 ( .A(n1261), .B(n1305), .C(n1679), .Y(n2017) );
  NAND2X1 U1557 ( .A(\mem<10><12> ), .B(n61), .Y(n1680) );
  OAI21X1 U1558 ( .A(n1261), .B(n1307), .C(n1680), .Y(n2016) );
  NAND2X1 U1559 ( .A(\mem<10><13> ), .B(n61), .Y(n1681) );
  OAI21X1 U1560 ( .A(n1261), .B(n1309), .C(n1681), .Y(n2015) );
  NAND2X1 U1561 ( .A(\mem<10><14> ), .B(n61), .Y(n1682) );
  OAI21X1 U1562 ( .A(n1261), .B(n1311), .C(n1682), .Y(n2014) );
  NAND2X1 U1563 ( .A(\mem<10><15> ), .B(n61), .Y(n1683) );
  OAI21X1 U1564 ( .A(n1261), .B(n1313), .C(n1683), .Y(n2013) );
  NAND2X1 U1565 ( .A(\mem<9><0> ), .B(n63), .Y(n1684) );
  OAI21X1 U1566 ( .A(n1262), .B(n1284), .C(n1684), .Y(n2012) );
  NAND2X1 U1567 ( .A(\mem<9><1> ), .B(n63), .Y(n1685) );
  OAI21X1 U1568 ( .A(n1262), .B(n1285), .C(n1685), .Y(n2011) );
  NAND2X1 U1569 ( .A(\mem<9><2> ), .B(n63), .Y(n1686) );
  OAI21X1 U1570 ( .A(n1262), .B(n1287), .C(n1686), .Y(n2010) );
  NAND2X1 U1571 ( .A(\mem<9><3> ), .B(n63), .Y(n1687) );
  OAI21X1 U1572 ( .A(n1262), .B(n1289), .C(n1687), .Y(n2009) );
  NAND2X1 U1573 ( .A(\mem<9><4> ), .B(n63), .Y(n1688) );
  OAI21X1 U1574 ( .A(n1262), .B(n1291), .C(n1688), .Y(n2008) );
  NAND2X1 U1575 ( .A(\mem<9><5> ), .B(n63), .Y(n1689) );
  OAI21X1 U1576 ( .A(n1262), .B(n1293), .C(n1689), .Y(n2007) );
  NAND2X1 U1577 ( .A(\mem<9><6> ), .B(n63), .Y(n1690) );
  OAI21X1 U1578 ( .A(n1262), .B(n1295), .C(n1690), .Y(n2006) );
  NAND2X1 U1579 ( .A(\mem<9><7> ), .B(n63), .Y(n1691) );
  OAI21X1 U1580 ( .A(n1262), .B(n1297), .C(n1691), .Y(n2005) );
  NAND2X1 U1581 ( .A(\mem<9><8> ), .B(n63), .Y(n1692) );
  OAI21X1 U1582 ( .A(n1263), .B(n1299), .C(n1692), .Y(n2004) );
  NAND2X1 U1583 ( .A(\mem<9><9> ), .B(n63), .Y(n1693) );
  OAI21X1 U1584 ( .A(n1263), .B(n1301), .C(n1693), .Y(n2003) );
  NAND2X1 U1585 ( .A(\mem<9><10> ), .B(n63), .Y(n1694) );
  OAI21X1 U1586 ( .A(n1263), .B(n1303), .C(n1694), .Y(n2002) );
  NAND2X1 U1587 ( .A(\mem<9><11> ), .B(n63), .Y(n1695) );
  OAI21X1 U1588 ( .A(n1263), .B(n1305), .C(n1695), .Y(n2001) );
  NAND2X1 U1589 ( .A(\mem<9><12> ), .B(n63), .Y(n1696) );
  OAI21X1 U1590 ( .A(n1263), .B(n1307), .C(n1696), .Y(n2000) );
  NAND2X1 U1591 ( .A(\mem<9><13> ), .B(n63), .Y(n1697) );
  OAI21X1 U1592 ( .A(n1263), .B(n1309), .C(n1697), .Y(n1999) );
  NAND2X1 U1593 ( .A(\mem<9><14> ), .B(n63), .Y(n1698) );
  OAI21X1 U1594 ( .A(n1263), .B(n1311), .C(n1698), .Y(n1998) );
  NAND2X1 U1595 ( .A(\mem<9><15> ), .B(n63), .Y(n1699) );
  OAI21X1 U1596 ( .A(n1263), .B(n1313), .C(n1699), .Y(n1997) );
  NAND2X1 U1597 ( .A(\mem<8><0> ), .B(n65), .Y(n1701) );
  OAI21X1 U1598 ( .A(n1264), .B(n1284), .C(n1701), .Y(n1996) );
  NAND2X1 U1599 ( .A(\mem<8><1> ), .B(n65), .Y(n1702) );
  OAI21X1 U1600 ( .A(n1264), .B(n1285), .C(n1702), .Y(n1995) );
  NAND2X1 U1601 ( .A(\mem<8><2> ), .B(n65), .Y(n1703) );
  OAI21X1 U1602 ( .A(n1264), .B(n1287), .C(n1703), .Y(n1994) );
  NAND2X1 U1603 ( .A(\mem<8><3> ), .B(n65), .Y(n1704) );
  OAI21X1 U1604 ( .A(n1264), .B(n1289), .C(n1704), .Y(n1993) );
  NAND2X1 U1605 ( .A(\mem<8><4> ), .B(n65), .Y(n1705) );
  OAI21X1 U1606 ( .A(n1264), .B(n1291), .C(n1705), .Y(n1992) );
  NAND2X1 U1607 ( .A(\mem<8><5> ), .B(n65), .Y(n1706) );
  OAI21X1 U1608 ( .A(n1264), .B(n1293), .C(n1706), .Y(n1991) );
  NAND2X1 U1609 ( .A(\mem<8><6> ), .B(n65), .Y(n1707) );
  OAI21X1 U1610 ( .A(n1264), .B(n1295), .C(n1707), .Y(n1990) );
  NAND2X1 U1611 ( .A(\mem<8><7> ), .B(n65), .Y(n1708) );
  OAI21X1 U1612 ( .A(n1264), .B(n1297), .C(n1708), .Y(n1989) );
  NAND2X1 U1613 ( .A(\mem<8><8> ), .B(n65), .Y(n1709) );
  OAI21X1 U1614 ( .A(n1264), .B(n1299), .C(n1709), .Y(n1988) );
  NAND2X1 U1615 ( .A(\mem<8><9> ), .B(n65), .Y(n1710) );
  OAI21X1 U1616 ( .A(n1264), .B(n1301), .C(n1710), .Y(n1987) );
  NAND2X1 U1617 ( .A(\mem<8><10> ), .B(n65), .Y(n1711) );
  OAI21X1 U1618 ( .A(n1264), .B(n1303), .C(n1711), .Y(n1986) );
  NAND2X1 U1619 ( .A(\mem<8><11> ), .B(n65), .Y(n1712) );
  OAI21X1 U1620 ( .A(n1264), .B(n1305), .C(n1712), .Y(n1985) );
  NAND2X1 U1621 ( .A(\mem<8><12> ), .B(n65), .Y(n1713) );
  OAI21X1 U1622 ( .A(n1264), .B(n1307), .C(n1713), .Y(n1984) );
  NAND2X1 U1623 ( .A(\mem<8><13> ), .B(n65), .Y(n1714) );
  OAI21X1 U1624 ( .A(n1264), .B(n1309), .C(n1714), .Y(n1983) );
  NAND2X1 U1625 ( .A(\mem<8><14> ), .B(n65), .Y(n1715) );
  OAI21X1 U1626 ( .A(n1264), .B(n1311), .C(n1715), .Y(n1982) );
  NAND2X1 U1627 ( .A(\mem<8><15> ), .B(n65), .Y(n1716) );
  OAI21X1 U1628 ( .A(n1264), .B(n1313), .C(n1716), .Y(n1981) );
  NAND3X1 U1629 ( .A(n1323), .B(n2365), .C(n1325), .Y(n1717) );
  NAND2X1 U1630 ( .A(\mem<7><0> ), .B(n67), .Y(n1718) );
  OAI21X1 U1631 ( .A(n1265), .B(n1283), .C(n1718), .Y(n1980) );
  NAND2X1 U1632 ( .A(\mem<7><1> ), .B(n67), .Y(n1719) );
  OAI21X1 U1633 ( .A(n1265), .B(n1285), .C(n1719), .Y(n1979) );
  NAND2X1 U1634 ( .A(\mem<7><2> ), .B(n67), .Y(n1720) );
  OAI21X1 U1635 ( .A(n1265), .B(n1287), .C(n1720), .Y(n1978) );
  NAND2X1 U1636 ( .A(\mem<7><3> ), .B(n67), .Y(n1721) );
  OAI21X1 U1637 ( .A(n1265), .B(n1289), .C(n1721), .Y(n1977) );
  NAND2X1 U1638 ( .A(\mem<7><4> ), .B(n67), .Y(n1722) );
  OAI21X1 U1639 ( .A(n1265), .B(n1291), .C(n1722), .Y(n1976) );
  NAND2X1 U1640 ( .A(\mem<7><5> ), .B(n67), .Y(n1723) );
  OAI21X1 U1641 ( .A(n1265), .B(n1293), .C(n1723), .Y(n1975) );
  NAND2X1 U1642 ( .A(\mem<7><6> ), .B(n67), .Y(n1724) );
  OAI21X1 U1643 ( .A(n1265), .B(n1295), .C(n1724), .Y(n1974) );
  NAND2X1 U1644 ( .A(\mem<7><7> ), .B(n67), .Y(n1725) );
  OAI21X1 U1645 ( .A(n1265), .B(n1297), .C(n1725), .Y(n1973) );
  NAND2X1 U1646 ( .A(\mem<7><8> ), .B(n67), .Y(n1726) );
  OAI21X1 U1647 ( .A(n1266), .B(n1299), .C(n1726), .Y(n1972) );
  NAND2X1 U1648 ( .A(\mem<7><9> ), .B(n67), .Y(n1727) );
  OAI21X1 U1649 ( .A(n1266), .B(n1301), .C(n1727), .Y(n1971) );
  NAND2X1 U1650 ( .A(\mem<7><10> ), .B(n67), .Y(n1728) );
  OAI21X1 U1651 ( .A(n1266), .B(n1303), .C(n1728), .Y(n1970) );
  NAND2X1 U1652 ( .A(\mem<7><11> ), .B(n67), .Y(n1729) );
  OAI21X1 U1653 ( .A(n1266), .B(n1305), .C(n1729), .Y(n1969) );
  NAND2X1 U1654 ( .A(\mem<7><12> ), .B(n67), .Y(n1730) );
  OAI21X1 U1655 ( .A(n1266), .B(n1307), .C(n1730), .Y(n1968) );
  NAND2X1 U1656 ( .A(\mem<7><13> ), .B(n67), .Y(n1731) );
  OAI21X1 U1657 ( .A(n1266), .B(n1309), .C(n1731), .Y(n1967) );
  NAND2X1 U1658 ( .A(\mem<7><14> ), .B(n67), .Y(n1732) );
  OAI21X1 U1659 ( .A(n1266), .B(n1311), .C(n1732), .Y(n1966) );
  NAND2X1 U1660 ( .A(\mem<7><15> ), .B(n67), .Y(n1733) );
  OAI21X1 U1661 ( .A(n1266), .B(n1313), .C(n1733), .Y(n1965) );
  NAND2X1 U1662 ( .A(\mem<6><0> ), .B(n69), .Y(n1734) );
  OAI21X1 U1663 ( .A(n1267), .B(n1284), .C(n1734), .Y(n1964) );
  NAND2X1 U1664 ( .A(\mem<6><1> ), .B(n69), .Y(n1735) );
  OAI21X1 U1665 ( .A(n1267), .B(n1285), .C(n1735), .Y(n1963) );
  NAND2X1 U1666 ( .A(\mem<6><2> ), .B(n69), .Y(n1736) );
  OAI21X1 U1667 ( .A(n1267), .B(n1287), .C(n1736), .Y(n1962) );
  NAND2X1 U1668 ( .A(\mem<6><3> ), .B(n69), .Y(n1737) );
  OAI21X1 U1669 ( .A(n1267), .B(n1289), .C(n1737), .Y(n1961) );
  NAND2X1 U1670 ( .A(\mem<6><4> ), .B(n69), .Y(n1738) );
  OAI21X1 U1671 ( .A(n1267), .B(n1291), .C(n1738), .Y(n1960) );
  NAND2X1 U1672 ( .A(\mem<6><5> ), .B(n69), .Y(n1739) );
  OAI21X1 U1673 ( .A(n1267), .B(n1293), .C(n1739), .Y(n1959) );
  NAND2X1 U1674 ( .A(\mem<6><6> ), .B(n69), .Y(n1740) );
  OAI21X1 U1675 ( .A(n1267), .B(n1295), .C(n1740), .Y(n1958) );
  NAND2X1 U1676 ( .A(\mem<6><7> ), .B(n69), .Y(n1741) );
  OAI21X1 U1677 ( .A(n1267), .B(n1297), .C(n1741), .Y(n1957) );
  NAND2X1 U1678 ( .A(\mem<6><8> ), .B(n69), .Y(n1742) );
  OAI21X1 U1679 ( .A(n1268), .B(n1299), .C(n1742), .Y(n1956) );
  NAND2X1 U1680 ( .A(\mem<6><9> ), .B(n69), .Y(n1743) );
  OAI21X1 U1681 ( .A(n1268), .B(n1301), .C(n1743), .Y(n1955) );
  NAND2X1 U1682 ( .A(\mem<6><10> ), .B(n69), .Y(n1744) );
  OAI21X1 U1683 ( .A(n1268), .B(n1303), .C(n1744), .Y(n1954) );
  NAND2X1 U1684 ( .A(\mem<6><11> ), .B(n69), .Y(n1745) );
  OAI21X1 U1685 ( .A(n1268), .B(n1305), .C(n1745), .Y(n1953) );
  NAND2X1 U1686 ( .A(\mem<6><12> ), .B(n69), .Y(n1746) );
  OAI21X1 U1687 ( .A(n1268), .B(n1307), .C(n1746), .Y(n1952) );
  NAND2X1 U1688 ( .A(\mem<6><13> ), .B(n69), .Y(n1747) );
  OAI21X1 U1689 ( .A(n1268), .B(n1309), .C(n1747), .Y(n1951) );
  NAND2X1 U1690 ( .A(\mem<6><14> ), .B(n69), .Y(n1748) );
  OAI21X1 U1691 ( .A(n1268), .B(n1311), .C(n1748), .Y(n1950) );
  NAND2X1 U1692 ( .A(\mem<6><15> ), .B(n69), .Y(n1749) );
  OAI21X1 U1693 ( .A(n1268), .B(n1313), .C(n1749), .Y(n1949) );
  NAND2X1 U1694 ( .A(\mem<5><0> ), .B(n71), .Y(n1751) );
  OAI21X1 U1695 ( .A(n1269), .B(n1283), .C(n1751), .Y(n1948) );
  NAND2X1 U1696 ( .A(\mem<5><1> ), .B(n71), .Y(n1752) );
  OAI21X1 U1697 ( .A(n1269), .B(n1285), .C(n1752), .Y(n1947) );
  NAND2X1 U1698 ( .A(\mem<5><2> ), .B(n71), .Y(n1753) );
  OAI21X1 U1699 ( .A(n1269), .B(n1287), .C(n1753), .Y(n1946) );
  NAND2X1 U1700 ( .A(\mem<5><3> ), .B(n71), .Y(n1754) );
  OAI21X1 U1701 ( .A(n1269), .B(n1289), .C(n1754), .Y(n1945) );
  NAND2X1 U1702 ( .A(\mem<5><4> ), .B(n71), .Y(n1755) );
  OAI21X1 U1703 ( .A(n1269), .B(n1291), .C(n1755), .Y(n1944) );
  NAND2X1 U1704 ( .A(\mem<5><5> ), .B(n71), .Y(n1756) );
  OAI21X1 U1705 ( .A(n1269), .B(n1293), .C(n1756), .Y(n1943) );
  NAND2X1 U1706 ( .A(\mem<5><6> ), .B(n71), .Y(n1757) );
  OAI21X1 U1707 ( .A(n1269), .B(n1295), .C(n1757), .Y(n1942) );
  NAND2X1 U1708 ( .A(\mem<5><7> ), .B(n71), .Y(n1758) );
  OAI21X1 U1709 ( .A(n1269), .B(n1297), .C(n1758), .Y(n1941) );
  NAND2X1 U1710 ( .A(\mem<5><8> ), .B(n71), .Y(n1759) );
  OAI21X1 U1711 ( .A(n1270), .B(n1299), .C(n1759), .Y(n1940) );
  NAND2X1 U1712 ( .A(\mem<5><9> ), .B(n71), .Y(n1760) );
  OAI21X1 U1713 ( .A(n1270), .B(n1301), .C(n1760), .Y(n1939) );
  NAND2X1 U1714 ( .A(\mem<5><10> ), .B(n71), .Y(n1761) );
  OAI21X1 U1715 ( .A(n1270), .B(n1303), .C(n1761), .Y(n1938) );
  NAND2X1 U1716 ( .A(\mem<5><11> ), .B(n71), .Y(n1762) );
  OAI21X1 U1717 ( .A(n1270), .B(n1305), .C(n1762), .Y(n1937) );
  NAND2X1 U1718 ( .A(\mem<5><12> ), .B(n71), .Y(n1763) );
  OAI21X1 U1719 ( .A(n1270), .B(n1307), .C(n1763), .Y(n1936) );
  NAND2X1 U1720 ( .A(\mem<5><13> ), .B(n71), .Y(n1764) );
  OAI21X1 U1721 ( .A(n1270), .B(n1309), .C(n1764), .Y(n1935) );
  NAND2X1 U1722 ( .A(\mem<5><14> ), .B(n71), .Y(n1765) );
  OAI21X1 U1723 ( .A(n1270), .B(n1311), .C(n1765), .Y(n1934) );
  NAND2X1 U1724 ( .A(\mem<5><15> ), .B(n71), .Y(n1766) );
  OAI21X1 U1725 ( .A(n1270), .B(n1313), .C(n1766), .Y(n1933) );
  NAND2X1 U1726 ( .A(\mem<4><0> ), .B(n73), .Y(n1768) );
  OAI21X1 U1727 ( .A(n1271), .B(n1284), .C(n1768), .Y(n1932) );
  NAND2X1 U1728 ( .A(\mem<4><1> ), .B(n73), .Y(n1769) );
  OAI21X1 U1729 ( .A(n1271), .B(n1285), .C(n1769), .Y(n1931) );
  NAND2X1 U1730 ( .A(\mem<4><2> ), .B(n73), .Y(n1770) );
  OAI21X1 U1731 ( .A(n1271), .B(n1287), .C(n1770), .Y(n1930) );
  NAND2X1 U1732 ( .A(\mem<4><3> ), .B(n73), .Y(n1771) );
  OAI21X1 U1733 ( .A(n1271), .B(n1289), .C(n1771), .Y(n1929) );
  NAND2X1 U1734 ( .A(\mem<4><4> ), .B(n73), .Y(n1772) );
  OAI21X1 U1735 ( .A(n1271), .B(n1291), .C(n1772), .Y(n1928) );
  NAND2X1 U1736 ( .A(\mem<4><5> ), .B(n73), .Y(n1773) );
  OAI21X1 U1737 ( .A(n1271), .B(n1293), .C(n1773), .Y(n1927) );
  NAND2X1 U1738 ( .A(\mem<4><6> ), .B(n73), .Y(n1774) );
  OAI21X1 U1739 ( .A(n1271), .B(n1295), .C(n1774), .Y(n1926) );
  NAND2X1 U1740 ( .A(\mem<4><7> ), .B(n73), .Y(n1775) );
  OAI21X1 U1741 ( .A(n1271), .B(n1297), .C(n1775), .Y(n1925) );
  NAND2X1 U1742 ( .A(\mem<4><8> ), .B(n73), .Y(n1776) );
  OAI21X1 U1743 ( .A(n1272), .B(n1299), .C(n1776), .Y(n1924) );
  NAND2X1 U1744 ( .A(\mem<4><9> ), .B(n73), .Y(n1777) );
  OAI21X1 U1745 ( .A(n1272), .B(n1301), .C(n1777), .Y(n1923) );
  NAND2X1 U1746 ( .A(\mem<4><10> ), .B(n73), .Y(n1778) );
  OAI21X1 U1747 ( .A(n1272), .B(n1303), .C(n1778), .Y(n1922) );
  NAND2X1 U1748 ( .A(\mem<4><11> ), .B(n73), .Y(n1779) );
  OAI21X1 U1749 ( .A(n1272), .B(n1305), .C(n1779), .Y(n1921) );
  NAND2X1 U1750 ( .A(\mem<4><12> ), .B(n73), .Y(n1780) );
  OAI21X1 U1751 ( .A(n1272), .B(n1307), .C(n1780), .Y(n1920) );
  NAND2X1 U1752 ( .A(\mem<4><13> ), .B(n73), .Y(n1781) );
  OAI21X1 U1753 ( .A(n1272), .B(n1309), .C(n1781), .Y(n1919) );
  NAND2X1 U1754 ( .A(\mem<4><14> ), .B(n73), .Y(n1782) );
  OAI21X1 U1755 ( .A(n1272), .B(n1311), .C(n1782), .Y(n1918) );
  NAND2X1 U1756 ( .A(\mem<4><15> ), .B(n73), .Y(n1783) );
  OAI21X1 U1757 ( .A(n1272), .B(n1313), .C(n1783), .Y(n1917) );
  NAND2X1 U1758 ( .A(\mem<3><0> ), .B(n75), .Y(n1785) );
  OAI21X1 U1759 ( .A(n1273), .B(n1283), .C(n1785), .Y(n1916) );
  NAND2X1 U1760 ( .A(\mem<3><1> ), .B(n75), .Y(n1786) );
  OAI21X1 U1761 ( .A(n1273), .B(n1285), .C(n1786), .Y(n1915) );
  NAND2X1 U1762 ( .A(\mem<3><2> ), .B(n75), .Y(n1787) );
  OAI21X1 U1763 ( .A(n1273), .B(n1287), .C(n1787), .Y(n1914) );
  NAND2X1 U1764 ( .A(\mem<3><3> ), .B(n75), .Y(n1788) );
  OAI21X1 U1765 ( .A(n1273), .B(n1289), .C(n1788), .Y(n1913) );
  NAND2X1 U1766 ( .A(\mem<3><4> ), .B(n75), .Y(n1789) );
  OAI21X1 U1767 ( .A(n1273), .B(n1291), .C(n1789), .Y(n1912) );
  NAND2X1 U1768 ( .A(\mem<3><5> ), .B(n75), .Y(n1790) );
  OAI21X1 U1769 ( .A(n1273), .B(n1293), .C(n1790), .Y(n1911) );
  NAND2X1 U1770 ( .A(\mem<3><6> ), .B(n75), .Y(n1791) );
  OAI21X1 U1771 ( .A(n1273), .B(n1295), .C(n1791), .Y(n1910) );
  NAND2X1 U1772 ( .A(\mem<3><7> ), .B(n75), .Y(n1792) );
  OAI21X1 U1773 ( .A(n1273), .B(n1297), .C(n1792), .Y(n1909) );
  NAND2X1 U1774 ( .A(\mem<3><8> ), .B(n75), .Y(n1793) );
  OAI21X1 U1775 ( .A(n1274), .B(n1299), .C(n1793), .Y(n1908) );
  NAND2X1 U1776 ( .A(\mem<3><9> ), .B(n75), .Y(n1794) );
  OAI21X1 U1777 ( .A(n1274), .B(n1301), .C(n1794), .Y(n1907) );
  NAND2X1 U1778 ( .A(\mem<3><10> ), .B(n75), .Y(n1795) );
  OAI21X1 U1779 ( .A(n1274), .B(n1303), .C(n1795), .Y(n1906) );
  NAND2X1 U1780 ( .A(\mem<3><11> ), .B(n75), .Y(n1796) );
  OAI21X1 U1781 ( .A(n1274), .B(n1305), .C(n1796), .Y(n1905) );
  NAND2X1 U1782 ( .A(\mem<3><12> ), .B(n75), .Y(n1797) );
  OAI21X1 U1783 ( .A(n1274), .B(n1307), .C(n1797), .Y(n1904) );
  NAND2X1 U1784 ( .A(\mem<3><13> ), .B(n75), .Y(n1798) );
  OAI21X1 U1785 ( .A(n1274), .B(n1309), .C(n1798), .Y(n1903) );
  NAND2X1 U1786 ( .A(\mem<3><14> ), .B(n75), .Y(n1799) );
  OAI21X1 U1787 ( .A(n1274), .B(n1311), .C(n1799), .Y(n1902) );
  NAND2X1 U1788 ( .A(\mem<3><15> ), .B(n75), .Y(n1800) );
  OAI21X1 U1789 ( .A(n1274), .B(n1313), .C(n1800), .Y(n1901) );
  NAND2X1 U1790 ( .A(\mem<2><0> ), .B(n77), .Y(n1802) );
  OAI21X1 U1791 ( .A(n1275), .B(n1284), .C(n1802), .Y(n1900) );
  NAND2X1 U1792 ( .A(\mem<2><1> ), .B(n77), .Y(n1803) );
  OAI21X1 U1793 ( .A(n1275), .B(n1285), .C(n1803), .Y(n1899) );
  NAND2X1 U1794 ( .A(\mem<2><2> ), .B(n77), .Y(n1804) );
  OAI21X1 U1795 ( .A(n1275), .B(n1287), .C(n1804), .Y(n1898) );
  NAND2X1 U1796 ( .A(\mem<2><3> ), .B(n77), .Y(n1805) );
  OAI21X1 U1797 ( .A(n1275), .B(n1289), .C(n1805), .Y(n1897) );
  NAND2X1 U1798 ( .A(\mem<2><4> ), .B(n77), .Y(n1806) );
  OAI21X1 U1799 ( .A(n1275), .B(n1291), .C(n1806), .Y(n1896) );
  NAND2X1 U1800 ( .A(\mem<2><5> ), .B(n77), .Y(n1807) );
  OAI21X1 U1801 ( .A(n1275), .B(n1293), .C(n1807), .Y(n1895) );
  NAND2X1 U1802 ( .A(\mem<2><6> ), .B(n77), .Y(n1808) );
  OAI21X1 U1803 ( .A(n1275), .B(n1295), .C(n1808), .Y(n1894) );
  NAND2X1 U1804 ( .A(\mem<2><7> ), .B(n77), .Y(n1809) );
  OAI21X1 U1805 ( .A(n1275), .B(n1297), .C(n1809), .Y(n1893) );
  NAND2X1 U1806 ( .A(\mem<2><8> ), .B(n77), .Y(n1810) );
  OAI21X1 U1807 ( .A(n1276), .B(n1299), .C(n1810), .Y(n1892) );
  NAND2X1 U1808 ( .A(\mem<2><9> ), .B(n77), .Y(n1811) );
  OAI21X1 U1809 ( .A(n1276), .B(n1301), .C(n1811), .Y(n1891) );
  NAND2X1 U1810 ( .A(\mem<2><10> ), .B(n77), .Y(n1812) );
  OAI21X1 U1811 ( .A(n1276), .B(n1303), .C(n1812), .Y(n1890) );
  NAND2X1 U1812 ( .A(\mem<2><11> ), .B(n77), .Y(n1813) );
  OAI21X1 U1813 ( .A(n1276), .B(n1305), .C(n1813), .Y(n1889) );
  NAND2X1 U1814 ( .A(\mem<2><12> ), .B(n77), .Y(n1814) );
  OAI21X1 U1815 ( .A(n1276), .B(n1307), .C(n1814), .Y(n1888) );
  NAND2X1 U1816 ( .A(\mem<2><13> ), .B(n77), .Y(n1815) );
  OAI21X1 U1817 ( .A(n1276), .B(n1309), .C(n1815), .Y(n1887) );
  NAND2X1 U1818 ( .A(\mem<2><14> ), .B(n77), .Y(n1816) );
  OAI21X1 U1819 ( .A(n1276), .B(n1311), .C(n1816), .Y(n1886) );
  NAND2X1 U1820 ( .A(\mem<2><15> ), .B(n77), .Y(n1817) );
  OAI21X1 U1821 ( .A(n1276), .B(n1313), .C(n1817), .Y(n1885) );
  NAND2X1 U1822 ( .A(\mem<1><0> ), .B(n37), .Y(n1819) );
  OAI21X1 U1823 ( .A(n1277), .B(n1283), .C(n1819), .Y(n1884) );
  NAND2X1 U1824 ( .A(\mem<1><1> ), .B(n37), .Y(n1820) );
  OAI21X1 U1825 ( .A(n1277), .B(n1285), .C(n1820), .Y(n1883) );
  NAND2X1 U1826 ( .A(\mem<1><2> ), .B(n37), .Y(n1821) );
  OAI21X1 U1827 ( .A(n1277), .B(n1287), .C(n1821), .Y(n1882) );
  NAND2X1 U1828 ( .A(\mem<1><3> ), .B(n37), .Y(n1822) );
  OAI21X1 U1829 ( .A(n1277), .B(n1289), .C(n1822), .Y(n1881) );
  NAND2X1 U1830 ( .A(\mem<1><4> ), .B(n37), .Y(n1823) );
  OAI21X1 U1831 ( .A(n1277), .B(n1291), .C(n1823), .Y(n1880) );
  NAND2X1 U1832 ( .A(\mem<1><5> ), .B(n37), .Y(n1824) );
  OAI21X1 U1833 ( .A(n1277), .B(n1293), .C(n1824), .Y(n1879) );
  NAND2X1 U1834 ( .A(\mem<1><6> ), .B(n37), .Y(n1825) );
  OAI21X1 U1835 ( .A(n1277), .B(n1295), .C(n1825), .Y(n1878) );
  NAND2X1 U1836 ( .A(\mem<1><7> ), .B(n37), .Y(n1826) );
  OAI21X1 U1837 ( .A(n1277), .B(n1297), .C(n1826), .Y(n1877) );
  NAND2X1 U1838 ( .A(\mem<1><8> ), .B(n37), .Y(n1827) );
  OAI21X1 U1839 ( .A(n1278), .B(n1299), .C(n1827), .Y(n1876) );
  NAND2X1 U1840 ( .A(\mem<1><9> ), .B(n37), .Y(n1828) );
  OAI21X1 U1841 ( .A(n1278), .B(n1301), .C(n1828), .Y(n1875) );
  NAND2X1 U1842 ( .A(\mem<1><10> ), .B(n37), .Y(n1829) );
  OAI21X1 U1843 ( .A(n1278), .B(n1303), .C(n1829), .Y(n1874) );
  NAND2X1 U1844 ( .A(\mem<1><11> ), .B(n37), .Y(n1830) );
  OAI21X1 U1845 ( .A(n1278), .B(n1305), .C(n1830), .Y(n1873) );
  NAND2X1 U1846 ( .A(\mem<1><12> ), .B(n37), .Y(n1831) );
  OAI21X1 U1847 ( .A(n1278), .B(n1307), .C(n1831), .Y(n1872) );
  NAND2X1 U1848 ( .A(\mem<1><13> ), .B(n37), .Y(n1832) );
  OAI21X1 U1849 ( .A(n1278), .B(n1309), .C(n1832), .Y(n1871) );
  NAND2X1 U1850 ( .A(\mem<1><14> ), .B(n37), .Y(n1833) );
  OAI21X1 U1851 ( .A(n1278), .B(n1311), .C(n1833), .Y(n1870) );
  NAND2X1 U1852 ( .A(\mem<1><15> ), .B(n37), .Y(n1834) );
  OAI21X1 U1853 ( .A(n1278), .B(n1313), .C(n1834), .Y(n1869) );
  NAND2X1 U1854 ( .A(\mem<0><0> ), .B(n83), .Y(n1837) );
  OAI21X1 U1855 ( .A(n1279), .B(n1284), .C(n1837), .Y(n1868) );
  NAND2X1 U1856 ( .A(\mem<0><1> ), .B(n83), .Y(n1838) );
  OAI21X1 U1857 ( .A(n1279), .B(n1285), .C(n1838), .Y(n1867) );
  NAND2X1 U1858 ( .A(\mem<0><2> ), .B(n83), .Y(n1839) );
  OAI21X1 U1859 ( .A(n1279), .B(n1287), .C(n1839), .Y(n1866) );
  NAND2X1 U1860 ( .A(\mem<0><3> ), .B(n83), .Y(n1840) );
  OAI21X1 U1861 ( .A(n1279), .B(n1289), .C(n1840), .Y(n1865) );
  NAND2X1 U1862 ( .A(\mem<0><4> ), .B(n83), .Y(n1841) );
  OAI21X1 U1863 ( .A(n1279), .B(n1291), .C(n1841), .Y(n1864) );
  NAND2X1 U1864 ( .A(\mem<0><5> ), .B(n83), .Y(n1842) );
  OAI21X1 U1865 ( .A(n1279), .B(n1293), .C(n1842), .Y(n1863) );
  NAND2X1 U1866 ( .A(\mem<0><6> ), .B(n83), .Y(n1843) );
  OAI21X1 U1867 ( .A(n1279), .B(n1295), .C(n1843), .Y(n1862) );
  NAND2X1 U1868 ( .A(\mem<0><7> ), .B(n83), .Y(n1844) );
  OAI21X1 U1869 ( .A(n1279), .B(n1297), .C(n1844), .Y(n1861) );
  NAND2X1 U1870 ( .A(\mem<0><8> ), .B(n83), .Y(n1845) );
  OAI21X1 U1871 ( .A(n1279), .B(n1299), .C(n1845), .Y(n1860) );
  NAND2X1 U1872 ( .A(\mem<0><9> ), .B(n83), .Y(n1846) );
  OAI21X1 U1873 ( .A(n1279), .B(n1301), .C(n1846), .Y(n1859) );
  NAND2X1 U1874 ( .A(\mem<0><10> ), .B(n83), .Y(n1847) );
  OAI21X1 U1875 ( .A(n1279), .B(n1303), .C(n1847), .Y(n1858) );
  NAND2X1 U1876 ( .A(\mem<0><11> ), .B(n83), .Y(n1848) );
  OAI21X1 U1877 ( .A(n1279), .B(n1305), .C(n1848), .Y(n1857) );
  NAND2X1 U1878 ( .A(\mem<0><12> ), .B(n83), .Y(n1849) );
  OAI21X1 U1879 ( .A(n1279), .B(n1307), .C(n1849), .Y(n1856) );
  NAND2X1 U1880 ( .A(\mem<0><13> ), .B(n83), .Y(n1850) );
  OAI21X1 U1881 ( .A(n1279), .B(n1309), .C(n1850), .Y(n1855) );
  NAND2X1 U1882 ( .A(\mem<0><14> ), .B(n83), .Y(n1851) );
  OAI21X1 U1883 ( .A(n1279), .B(n1311), .C(n1851), .Y(n1854) );
  NAND2X1 U1884 ( .A(\mem<0><15> ), .B(n83), .Y(n1852) );
  OAI21X1 U1885 ( .A(n1279), .B(n1313), .C(n1852), .Y(n1853) );
endmodule


module memc_Size16_5 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1850), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1851), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1852), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1853), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1854), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1855), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1856), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1857), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1858), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1859), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1860), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1861), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1862), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1863), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1864), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1865), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1866), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1867), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1868), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1869), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1870), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1871), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1872), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1873), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1874), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1875), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1876), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1877), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1878), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1879), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1880), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1881), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1882), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1883), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1884), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1885), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1886), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1887), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1888), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1889), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1890), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1891), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1892), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1893), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1894), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1895), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1896), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1897), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1898), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1899), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1900), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1901), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1902), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1903), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1904), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1905), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1906), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1907), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1908), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1909), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1910), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1911), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1912), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1913), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1914), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1915), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1916), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1917), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1918), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1919), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1920), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1921), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1922), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1923), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1924), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1925), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1926), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1927), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1928), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1929), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1930), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1931), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1932), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1933), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1934), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1935), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1936), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1937), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1938), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1939), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1940), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1941), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1942), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1943), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1944), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1945), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1946), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1947), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1948), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1949), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1950), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1951), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1952), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1953), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1954), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1955), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1956), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1957), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1958), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1959), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1960), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1961), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1962), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1963), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1964), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1965), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1966), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1967), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1968), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1969), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1970), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1971), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1972), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1973), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1974), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1975), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1976), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1977), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1978), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1979), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1980), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1981), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1982), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1983), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1984), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1985), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1986), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1987), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1988), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1989), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1990), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1991), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1992), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1993), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1994), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1995), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1996), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1997), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1998), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1999), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2000), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2001), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2002), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2003), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2004), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2005), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2006), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2007), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2008), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2009), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2010), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2011), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2012), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2013), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2014), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2015), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2016), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2017), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2018), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2019), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2020), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2021), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2022), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2023), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2024), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2025), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2026), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2027), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2028), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2029), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2030), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2031), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2032), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2033), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2034), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2035), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2036), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2037), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2038), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2039), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2040), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2041), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2042), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2043), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2044), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2045), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2046), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2047), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2048), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2049), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2050), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2051), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2052), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2053), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2054), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2055), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2056), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2057), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2058), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2059), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2060), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2061), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2062), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2063), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2064), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2065), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2066), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2067), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2068), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2069), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2070), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2071), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2072), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2073), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2074), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2075), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2076), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2077), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2078), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2079), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2080), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2081), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2082), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2083), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2084), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2085), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2086), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2087), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2088), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2089), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2090), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2091), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2092), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2093), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2094), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2095), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2096), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2097), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2098), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2099), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2100), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2101), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2102), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2103), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2104), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2105), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2106), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2107), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2108), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2109), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2110), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2111), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2112), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2113), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2114), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2115), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2116), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2117), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2118), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2119), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2120), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2121), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2122), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2123), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2124), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2125), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2126), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2127), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2128), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2129), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2130), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2131), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2132), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2133), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2134), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2135), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2136), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2137), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2138), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2139), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2140), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2141), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2142), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2143), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2144), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2145), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2146), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2147), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2148), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2149), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2150), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2151), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2152), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2153), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2154), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2155), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2156), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2157), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2158), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2159), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2160), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2161), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2162), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2163), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2164), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2165), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2166), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2167), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2168), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2169), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2170), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2171), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2172), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2173), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2174), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2175), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2176), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2177), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2178), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2179), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2180), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2181), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2182), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2183), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2184), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2185), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2186), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2187), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2188), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2189), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2190), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2191), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2192), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2193), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2194), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2195), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2196), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2197), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2198), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2199), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2200), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2201), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2202), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2203), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2204), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2205), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2206), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2207), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2208), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2209), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2210), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2211), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2212), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2213), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2214), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2215), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2216), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2217), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2218), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2219), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2220), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2221), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2222), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2223), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2224), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2225), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2226), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2227), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2228), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2229), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2230), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2231), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2232), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2233), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2234), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2235), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2236), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2237), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2238), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2239), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2240), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2241), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2242), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2243), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2244), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2245), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2246), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2247), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2248), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2249), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2250), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2251), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2252), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2253), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2254), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2255), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2256), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2257), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2258), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2259), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2260), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2261), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2262), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2263), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2264), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2265), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2266), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2267), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2268), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2269), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2270), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2271), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2272), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2273), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2274), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2275), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2276), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2277), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2278), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2279), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2280), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2281), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2282), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2283), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2284), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2285), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2286), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2287), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2288), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2289), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2290), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2291), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2292), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2293), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2294), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2295), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2296), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2297), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2298), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2299), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2300), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2301), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2302), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2303), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2304), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2305), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2306), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2307), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2308), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2309), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2310), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2311), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2312), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2313), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2314), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2315), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2316), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2317), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2318), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2319), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2320), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2321), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2322), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2323), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2324), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2325), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2326), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2327), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2328), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2329), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2330), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2331), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2332), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2333), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2334), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2335), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2336), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2337), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2338), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2339), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2340), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2341), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2342), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2343), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2344), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2345), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2346), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2347), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2348), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2349), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2350), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2351), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2352), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2353), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2354), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2355), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2356), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2357), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2358), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2359), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2360), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2361), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2362) );
  INVX4 U2 ( .A(n73), .Y(n1280) );
  INVX1 U3 ( .A(n640), .Y(N32) );
  INVX1 U4 ( .A(n641), .Y(N31) );
  INVX1 U5 ( .A(n642), .Y(N30) );
  INVX1 U6 ( .A(n643), .Y(N29) );
  INVX1 U7 ( .A(n644), .Y(N28) );
  INVX1 U8 ( .A(n645), .Y(N27) );
  INVX1 U9 ( .A(n646), .Y(N26) );
  INVX1 U10 ( .A(n647), .Y(N25) );
  INVX1 U11 ( .A(n648), .Y(N24) );
  INVX1 U12 ( .A(n649), .Y(N23) );
  INVX1 U13 ( .A(n650), .Y(N22) );
  INVX1 U14 ( .A(n1163), .Y(N21) );
  INVX1 U15 ( .A(n1164), .Y(N20) );
  INVX1 U16 ( .A(n1165), .Y(N19) );
  INVX1 U17 ( .A(n1166), .Y(N18) );
  INVX1 U18 ( .A(n1167), .Y(N17) );
  INVX1 U19 ( .A(n1176), .Y(n1177) );
  INVX1 U20 ( .A(n1176), .Y(n1178) );
  INVX1 U21 ( .A(n1318), .Y(n1174) );
  INVX2 U22 ( .A(n1176), .Y(n1179) );
  INVX1 U23 ( .A(n1188), .Y(n1180) );
  INVX1 U24 ( .A(n1318), .Y(n1173) );
  INVX1 U25 ( .A(n1188), .Y(n1181) );
  INVX2 U26 ( .A(n1188), .Y(n1182) );
  INVX1 U27 ( .A(n1318), .Y(n1172) );
  INVX1 U28 ( .A(n1175), .Y(n1183) );
  INVX1 U29 ( .A(n1175), .Y(n1184) );
  INVX2 U30 ( .A(n1175), .Y(n1185) );
  INVX2 U31 ( .A(n1176), .Y(n1186) );
  INVX2 U32 ( .A(n1214), .Y(n1212) );
  INVX2 U33 ( .A(n1175), .Y(n1187) );
  BUFX2 U34 ( .A(n104), .Y(n1218) );
  BUFX2 U35 ( .A(n106), .Y(n1220) );
  BUFX2 U36 ( .A(n108), .Y(n1222) );
  BUFX2 U37 ( .A(n110), .Y(n1224) );
  BUFX2 U38 ( .A(n112), .Y(n1226) );
  BUFX2 U39 ( .A(n114), .Y(n1228) );
  BUFX2 U40 ( .A(n116), .Y(n1230) );
  BUFX2 U41 ( .A(n118), .Y(n1233) );
  BUFX2 U42 ( .A(n120), .Y(n1235) );
  BUFX2 U43 ( .A(n122), .Y(n1237) );
  BUFX2 U44 ( .A(n124), .Y(n1239) );
  BUFX2 U45 ( .A(n126), .Y(n1241) );
  BUFX2 U46 ( .A(n128), .Y(n1243) );
  BUFX2 U47 ( .A(n130), .Y(n1245) );
  BUFX2 U48 ( .A(n132), .Y(n1248) );
  BUFX2 U49 ( .A(n134), .Y(n1250) );
  BUFX2 U50 ( .A(n136), .Y(n1252) );
  BUFX2 U51 ( .A(n138), .Y(n1254) );
  BUFX2 U52 ( .A(n140), .Y(n1256) );
  BUFX2 U53 ( .A(n142), .Y(n1258) );
  BUFX2 U54 ( .A(n144), .Y(n1260) );
  BUFX2 U55 ( .A(n146), .Y(n1263) );
  BUFX2 U56 ( .A(n148), .Y(n1265) );
  BUFX2 U57 ( .A(n150), .Y(n1267) );
  BUFX2 U58 ( .A(n152), .Y(n1269) );
  BUFX2 U59 ( .A(n154), .Y(n1271) );
  BUFX2 U60 ( .A(n156), .Y(n1273) );
  BUFX2 U61 ( .A(n158), .Y(n1275) );
  INVX2 U62 ( .A(n74), .Y(n1) );
  INVX2 U63 ( .A(n74), .Y(n75) );
  BUFX2 U64 ( .A(write), .Y(n2) );
  INVX1 U65 ( .A(n1214), .Y(n1215) );
  INVX1 U66 ( .A(n1313), .Y(n1214) );
  INVX1 U67 ( .A(n1315), .Y(n1188) );
  INVX1 U68 ( .A(n1322), .Y(n1168) );
  INVX1 U69 ( .A(n1214), .Y(n1217) );
  INVX2 U70 ( .A(n1217), .Y(n1191) );
  INVX2 U71 ( .A(n1217), .Y(n1192) );
  INVX1 U72 ( .A(n1320), .Y(n1169) );
  INVX1 U73 ( .A(n1214), .Y(n1216) );
  INVX2 U74 ( .A(n1216), .Y(n1189) );
  INVX2 U75 ( .A(n1216), .Y(n1190) );
  INVX1 U76 ( .A(N12), .Y(n1318) );
  INVX1 U77 ( .A(n1318), .Y(n1170) );
  INVX1 U78 ( .A(n1318), .Y(n1171) );
  INVX1 U79 ( .A(n1320), .Y(n1319) );
  INVX1 U80 ( .A(N13), .Y(n1320) );
  INVX1 U81 ( .A(n1322), .Y(n1321) );
  INVX1 U82 ( .A(N14), .Y(n1322) );
  INVX1 U83 ( .A(n1315), .Y(n1175) );
  INVX1 U84 ( .A(n1315), .Y(n1176) );
  INVX1 U85 ( .A(rst), .Y(n1312) );
  INVX1 U86 ( .A(n100), .Y(n1247) );
  INVX1 U87 ( .A(n101), .Y(n1262) );
  INVX1 U88 ( .A(n102), .Y(n1277) );
  BUFX2 U89 ( .A(n104), .Y(n1219) );
  BUFX2 U90 ( .A(n118), .Y(n1234) );
  BUFX2 U91 ( .A(n132), .Y(n1249) );
  BUFX2 U92 ( .A(n146), .Y(n1264) );
  BUFX2 U93 ( .A(n106), .Y(n1221) );
  BUFX2 U94 ( .A(n108), .Y(n1223) );
  BUFX2 U95 ( .A(n110), .Y(n1225) );
  BUFX2 U96 ( .A(n112), .Y(n1227) );
  BUFX2 U97 ( .A(n114), .Y(n1229) );
  BUFX2 U98 ( .A(n116), .Y(n1231) );
  BUFX2 U99 ( .A(n120), .Y(n1236) );
  BUFX2 U100 ( .A(n122), .Y(n1238) );
  BUFX2 U101 ( .A(n124), .Y(n1240) );
  BUFX2 U102 ( .A(n126), .Y(n1242) );
  BUFX2 U103 ( .A(n128), .Y(n1244) );
  BUFX2 U104 ( .A(n130), .Y(n1246) );
  BUFX2 U105 ( .A(n134), .Y(n1251) );
  BUFX2 U106 ( .A(n136), .Y(n1253) );
  BUFX2 U107 ( .A(n138), .Y(n1255) );
  BUFX2 U108 ( .A(n140), .Y(n1257) );
  BUFX2 U109 ( .A(n142), .Y(n1259) );
  BUFX2 U110 ( .A(n144), .Y(n1261) );
  BUFX2 U111 ( .A(n148), .Y(n1266) );
  BUFX2 U112 ( .A(n150), .Y(n1268) );
  BUFX2 U113 ( .A(n152), .Y(n1270) );
  BUFX2 U114 ( .A(n154), .Y(n1272) );
  BUFX2 U115 ( .A(n156), .Y(n1274) );
  BUFX2 U116 ( .A(n158), .Y(n1276) );
  INVX1 U117 ( .A(n99), .Y(n1232) );
  INVX4 U118 ( .A(n53), .Y(n54) );
  INVX4 U119 ( .A(n51), .Y(n52) );
  INVX4 U120 ( .A(n49), .Y(n50) );
  INVX4 U121 ( .A(n47), .Y(n48) );
  INVX4 U122 ( .A(n45), .Y(n46) );
  INVX4 U123 ( .A(n43), .Y(n44) );
  INVX4 U124 ( .A(n41), .Y(n42) );
  INVX4 U125 ( .A(n37), .Y(n38) );
  INVX4 U126 ( .A(n35), .Y(n36) );
  INVX4 U127 ( .A(n33), .Y(n34) );
  INVX4 U128 ( .A(n31), .Y(n32) );
  INVX4 U129 ( .A(n29), .Y(n30) );
  INVX4 U130 ( .A(n27), .Y(n28) );
  INVX4 U131 ( .A(n25), .Y(n26) );
  INVX4 U132 ( .A(n21), .Y(n22) );
  INVX4 U133 ( .A(n19), .Y(n20) );
  INVX4 U134 ( .A(n17), .Y(n18) );
  INVX4 U135 ( .A(n15), .Y(n16) );
  INVX4 U136 ( .A(n13), .Y(n14) );
  INVX4 U137 ( .A(n11), .Y(n12) );
  INVX4 U138 ( .A(n3), .Y(n4) );
  INVX4 U139 ( .A(n71), .Y(n72) );
  INVX4 U140 ( .A(n39), .Y(n40) );
  INVX4 U141 ( .A(n23), .Y(n24) );
  INVX4 U142 ( .A(n69), .Y(n70) );
  INVX4 U143 ( .A(n67), .Y(n68) );
  INVX4 U144 ( .A(n65), .Y(n66) );
  INVX4 U145 ( .A(n63), .Y(n64) );
  INVX4 U146 ( .A(n61), .Y(n62) );
  INVX4 U147 ( .A(n59), .Y(n60) );
  INVX4 U148 ( .A(n57), .Y(n58) );
  INVX4 U149 ( .A(n55), .Y(n56) );
  AND2X2 U150 ( .A(n1278), .B(n103), .Y(n3) );
  AND2X2 U151 ( .A(\data_in<7> ), .B(n1279), .Y(n5) );
  AND2X2 U152 ( .A(\data_in<11> ), .B(n1279), .Y(n6) );
  AND2X2 U153 ( .A(\data_in<12> ), .B(n1279), .Y(n7) );
  AND2X2 U154 ( .A(\data_in<13> ), .B(n1279), .Y(n8) );
  AND2X2 U155 ( .A(\data_in<14> ), .B(n1279), .Y(n9) );
  AND2X2 U156 ( .A(\data_in<15> ), .B(n1279), .Y(n10) );
  AND2X2 U157 ( .A(n1279), .B(n105), .Y(n11) );
  AND2X2 U158 ( .A(n1279), .B(n107), .Y(n13) );
  AND2X2 U159 ( .A(n1279), .B(n109), .Y(n15) );
  AND2X2 U160 ( .A(n1279), .B(n111), .Y(n17) );
  AND2X2 U161 ( .A(n1279), .B(n113), .Y(n19) );
  AND2X2 U162 ( .A(n1278), .B(n115), .Y(n21) );
  AND2X2 U163 ( .A(n1279), .B(n99), .Y(n23) );
  AND2X2 U164 ( .A(n1279), .B(n117), .Y(n25) );
  AND2X2 U165 ( .A(n1278), .B(n119), .Y(n27) );
  AND2X2 U166 ( .A(n1279), .B(n121), .Y(n29) );
  AND2X2 U167 ( .A(n1278), .B(n123), .Y(n31) );
  AND2X2 U168 ( .A(n1278), .B(n125), .Y(n33) );
  AND2X2 U169 ( .A(n1278), .B(n127), .Y(n35) );
  AND2X2 U170 ( .A(n1278), .B(n129), .Y(n37) );
  AND2X2 U171 ( .A(n1278), .B(n100), .Y(n39) );
  AND2X2 U172 ( .A(n1278), .B(n131), .Y(n41) );
  AND2X2 U173 ( .A(n1278), .B(n133), .Y(n43) );
  AND2X2 U174 ( .A(n1278), .B(n135), .Y(n45) );
  AND2X2 U175 ( .A(n1278), .B(n137), .Y(n47) );
  AND2X2 U176 ( .A(n1278), .B(n139), .Y(n49) );
  AND2X2 U177 ( .A(n1278), .B(n141), .Y(n51) );
  AND2X2 U178 ( .A(n1278), .B(n143), .Y(n53) );
  AND2X2 U179 ( .A(n1279), .B(n101), .Y(n55) );
  AND2X2 U180 ( .A(n1279), .B(n145), .Y(n57) );
  AND2X2 U181 ( .A(n1279), .B(n147), .Y(n59) );
  AND2X2 U182 ( .A(n1279), .B(n149), .Y(n61) );
  AND2X2 U183 ( .A(n1279), .B(n151), .Y(n63) );
  AND2X2 U184 ( .A(n1279), .B(n153), .Y(n65) );
  AND2X2 U185 ( .A(n1279), .B(n155), .Y(n67) );
  AND2X2 U186 ( .A(n1279), .B(n157), .Y(n69) );
  AND2X2 U187 ( .A(n1278), .B(n102), .Y(n71) );
  AND2X2 U188 ( .A(n2), .B(n1312), .Y(n73) );
  OR2X2 U189 ( .A(write), .B(rst), .Y(n74) );
  INVX1 U190 ( .A(n1318), .Y(n1317) );
  INVX1 U191 ( .A(n1314), .Y(n1313) );
  AND2X1 U192 ( .A(n1317), .B(n1315), .Y(n76) );
  INVX1 U193 ( .A(n1316), .Y(n1315) );
  AND2X1 U194 ( .A(n2362), .B(n1321), .Y(n77) );
  BUFX2 U195 ( .A(n1355), .Y(n78) );
  INVX1 U196 ( .A(n78), .Y(n1747) );
  BUFX2 U197 ( .A(n1372), .Y(n79) );
  INVX1 U198 ( .A(n79), .Y(n1764) );
  BUFX2 U199 ( .A(n1389), .Y(n80) );
  INVX1 U200 ( .A(n80), .Y(n1781) );
  BUFX2 U201 ( .A(n1406), .Y(n81) );
  INVX1 U202 ( .A(n81), .Y(n1798) );
  BUFX2 U203 ( .A(n1423), .Y(n82) );
  INVX1 U204 ( .A(n82), .Y(n1815) );
  BUFX2 U205 ( .A(n1584), .Y(n83) );
  INVX1 U206 ( .A(n83), .Y(n1697) );
  BUFX2 U207 ( .A(n1714), .Y(n84) );
  INVX1 U208 ( .A(n84), .Y(n1832) );
  AND2X1 U209 ( .A(n1313), .B(n76), .Y(n85) );
  AND2X1 U210 ( .A(n1319), .B(n77), .Y(n86) );
  AND2X1 U211 ( .A(n1314), .B(n76), .Y(n87) );
  AND2X1 U212 ( .A(n1320), .B(n77), .Y(n88) );
  AND2X2 U213 ( .A(\data_in<0> ), .B(n1278), .Y(n89) );
  AND2X2 U214 ( .A(\data_in<1> ), .B(n1278), .Y(n90) );
  AND2X2 U215 ( .A(\data_in<2> ), .B(n1278), .Y(n91) );
  AND2X2 U216 ( .A(\data_in<3> ), .B(n1279), .Y(n92) );
  AND2X2 U217 ( .A(\data_in<4> ), .B(n1279), .Y(n93) );
  AND2X2 U218 ( .A(\data_in<5> ), .B(n1278), .Y(n94) );
  AND2X2 U219 ( .A(\data_in<6> ), .B(n1278), .Y(n95) );
  AND2X2 U220 ( .A(\data_in<8> ), .B(n1278), .Y(n96) );
  AND2X2 U221 ( .A(\data_in<9> ), .B(n1278), .Y(n97) );
  AND2X2 U222 ( .A(\data_in<10> ), .B(n1278), .Y(n98) );
  AND2X1 U223 ( .A(n86), .B(n1833), .Y(n99) );
  AND2X1 U224 ( .A(n1833), .B(n88), .Y(n100) );
  AND2X1 U225 ( .A(n1833), .B(n1697), .Y(n101) );
  AND2X1 U226 ( .A(n1833), .B(n1832), .Y(n102) );
  AND2X1 U227 ( .A(n85), .B(n86), .Y(n103) );
  INVX1 U228 ( .A(n103), .Y(n104) );
  AND2X1 U229 ( .A(n86), .B(n87), .Y(n105) );
  INVX1 U230 ( .A(n105), .Y(n106) );
  AND2X1 U231 ( .A(n86), .B(n1747), .Y(n107) );
  INVX1 U232 ( .A(n107), .Y(n108) );
  AND2X1 U233 ( .A(n86), .B(n1764), .Y(n109) );
  INVX1 U234 ( .A(n109), .Y(n110) );
  AND2X1 U235 ( .A(n86), .B(n1781), .Y(n111) );
  INVX1 U236 ( .A(n111), .Y(n112) );
  AND2X1 U237 ( .A(n86), .B(n1798), .Y(n113) );
  INVX1 U238 ( .A(n113), .Y(n114) );
  AND2X1 U239 ( .A(n86), .B(n1815), .Y(n115) );
  INVX1 U240 ( .A(n115), .Y(n116) );
  AND2X1 U241 ( .A(n85), .B(n88), .Y(n117) );
  INVX1 U242 ( .A(n117), .Y(n118) );
  AND2X1 U243 ( .A(n87), .B(n88), .Y(n119) );
  INVX1 U244 ( .A(n119), .Y(n120) );
  AND2X1 U245 ( .A(n1747), .B(n88), .Y(n121) );
  INVX1 U246 ( .A(n121), .Y(n122) );
  AND2X1 U247 ( .A(n1764), .B(n88), .Y(n123) );
  INVX1 U248 ( .A(n123), .Y(n124) );
  AND2X1 U249 ( .A(n1781), .B(n88), .Y(n125) );
  INVX1 U250 ( .A(n125), .Y(n126) );
  AND2X1 U251 ( .A(n1798), .B(n88), .Y(n127) );
  INVX1 U252 ( .A(n127), .Y(n128) );
  AND2X1 U253 ( .A(n1815), .B(n88), .Y(n129) );
  INVX1 U254 ( .A(n129), .Y(n130) );
  AND2X1 U255 ( .A(n85), .B(n1697), .Y(n131) );
  INVX1 U256 ( .A(n131), .Y(n132) );
  AND2X1 U257 ( .A(n87), .B(n1697), .Y(n133) );
  INVX1 U258 ( .A(n133), .Y(n134) );
  AND2X1 U259 ( .A(n1747), .B(n1697), .Y(n135) );
  INVX1 U260 ( .A(n135), .Y(n136) );
  AND2X1 U261 ( .A(n1764), .B(n1697), .Y(n137) );
  INVX1 U262 ( .A(n137), .Y(n138) );
  AND2X1 U263 ( .A(n1781), .B(n1697), .Y(n139) );
  INVX1 U264 ( .A(n139), .Y(n140) );
  AND2X1 U265 ( .A(n1798), .B(n1697), .Y(n141) );
  INVX1 U266 ( .A(n141), .Y(n142) );
  AND2X1 U267 ( .A(n1815), .B(n1697), .Y(n143) );
  INVX1 U268 ( .A(n143), .Y(n144) );
  AND2X1 U269 ( .A(n85), .B(n1832), .Y(n145) );
  INVX1 U270 ( .A(n145), .Y(n146) );
  AND2X1 U271 ( .A(n87), .B(n1832), .Y(n147) );
  INVX1 U272 ( .A(n147), .Y(n148) );
  AND2X1 U273 ( .A(n1747), .B(n1832), .Y(n149) );
  INVX1 U274 ( .A(n149), .Y(n150) );
  AND2X1 U275 ( .A(n1764), .B(n1832), .Y(n151) );
  INVX1 U276 ( .A(n151), .Y(n152) );
  AND2X1 U277 ( .A(n1781), .B(n1832), .Y(n153) );
  INVX1 U278 ( .A(n153), .Y(n154) );
  AND2X1 U279 ( .A(n1798), .B(n1832), .Y(n155) );
  INVX1 U280 ( .A(n155), .Y(n156) );
  AND2X1 U281 ( .A(n1815), .B(n1832), .Y(n157) );
  INVX1 U282 ( .A(n157), .Y(n158) );
  AND2X2 U283 ( .A(n1), .B(N32), .Y(\data_out<0> ) );
  MUX2X1 U284 ( .B(n160), .A(n161), .S(n1177), .Y(n159) );
  MUX2X1 U285 ( .B(n163), .A(n164), .S(n1177), .Y(n162) );
  MUX2X1 U286 ( .B(n166), .A(n167), .S(n1177), .Y(n165) );
  MUX2X1 U287 ( .B(n169), .A(n170), .S(n1177), .Y(n168) );
  MUX2X1 U288 ( .B(n172), .A(n173), .S(n1169), .Y(n171) );
  MUX2X1 U289 ( .B(n175), .A(n176), .S(n1177), .Y(n174) );
  MUX2X1 U290 ( .B(n178), .A(n179), .S(n1177), .Y(n177) );
  MUX2X1 U291 ( .B(n181), .A(n182), .S(n1177), .Y(n180) );
  MUX2X1 U292 ( .B(n184), .A(n185), .S(n1177), .Y(n183) );
  MUX2X1 U293 ( .B(n187), .A(n188), .S(n1169), .Y(n186) );
  MUX2X1 U294 ( .B(n190), .A(n191), .S(n1178), .Y(n189) );
  MUX2X1 U295 ( .B(n193), .A(n194), .S(n1178), .Y(n192) );
  MUX2X1 U296 ( .B(n196), .A(n197), .S(n1178), .Y(n195) );
  MUX2X1 U297 ( .B(n199), .A(n200), .S(n1178), .Y(n198) );
  MUX2X1 U298 ( .B(n202), .A(n203), .S(n1169), .Y(n201) );
  MUX2X1 U299 ( .B(n205), .A(n206), .S(n1178), .Y(n204) );
  MUX2X1 U300 ( .B(n208), .A(n209), .S(n1178), .Y(n207) );
  MUX2X1 U301 ( .B(n211), .A(n212), .S(n1178), .Y(n210) );
  MUX2X1 U302 ( .B(n215), .A(n216), .S(n1178), .Y(n213) );
  MUX2X1 U303 ( .B(n218), .A(n219), .S(n1169), .Y(n217) );
  MUX2X1 U304 ( .B(n221), .A(n222), .S(n1178), .Y(n220) );
  MUX2X1 U305 ( .B(n224), .A(n225), .S(n1178), .Y(n223) );
  MUX2X1 U306 ( .B(n227), .A(n228), .S(n1178), .Y(n226) );
  MUX2X1 U307 ( .B(n230), .A(n231), .S(n1178), .Y(n229) );
  MUX2X1 U308 ( .B(n233), .A(n234), .S(n1169), .Y(n232) );
  MUX2X1 U309 ( .B(n236), .A(n237), .S(n1179), .Y(n235) );
  MUX2X1 U310 ( .B(n239), .A(n240), .S(n1179), .Y(n238) );
  MUX2X1 U311 ( .B(n242), .A(n243), .S(n1179), .Y(n241) );
  MUX2X1 U312 ( .B(n245), .A(n246), .S(n1179), .Y(n244) );
  MUX2X1 U313 ( .B(n248), .A(n249), .S(n1169), .Y(n247) );
  MUX2X1 U314 ( .B(n251), .A(n252), .S(n1179), .Y(n250) );
  MUX2X1 U315 ( .B(n254), .A(n255), .S(n1179), .Y(n253) );
  MUX2X1 U316 ( .B(n257), .A(n258), .S(n1179), .Y(n256) );
  MUX2X1 U317 ( .B(n260), .A(n261), .S(n1179), .Y(n259) );
  MUX2X1 U318 ( .B(n263), .A(n264), .S(n1169), .Y(n262) );
  MUX2X1 U319 ( .B(n266), .A(n267), .S(n1179), .Y(n265) );
  MUX2X1 U320 ( .B(n269), .A(n270), .S(n1179), .Y(n268) );
  MUX2X1 U321 ( .B(n272), .A(n273), .S(n1179), .Y(n271) );
  MUX2X1 U322 ( .B(n275), .A(n276), .S(n1179), .Y(n274) );
  MUX2X1 U323 ( .B(n278), .A(n279), .S(n1169), .Y(n277) );
  MUX2X1 U324 ( .B(n281), .A(n282), .S(n1180), .Y(n280) );
  MUX2X1 U325 ( .B(n284), .A(n285), .S(n1180), .Y(n283) );
  MUX2X1 U326 ( .B(n287), .A(n288), .S(n1180), .Y(n286) );
  MUX2X1 U327 ( .B(n290), .A(n291), .S(n1180), .Y(n289) );
  MUX2X1 U328 ( .B(n293), .A(n294), .S(n1169), .Y(n292) );
  MUX2X1 U329 ( .B(n296), .A(n297), .S(n1180), .Y(n295) );
  MUX2X1 U330 ( .B(n299), .A(n300), .S(n1180), .Y(n298) );
  MUX2X1 U331 ( .B(n302), .A(n303), .S(n1180), .Y(n301) );
  MUX2X1 U332 ( .B(n305), .A(n306), .S(n1180), .Y(n304) );
  MUX2X1 U333 ( .B(n308), .A(n309), .S(n1169), .Y(n307) );
  MUX2X1 U334 ( .B(n311), .A(n312), .S(n1180), .Y(n310) );
  MUX2X1 U335 ( .B(n314), .A(n315), .S(n1180), .Y(n313) );
  MUX2X1 U336 ( .B(n317), .A(n318), .S(n1180), .Y(n316) );
  MUX2X1 U337 ( .B(n320), .A(n321), .S(n1180), .Y(n319) );
  MUX2X1 U338 ( .B(n323), .A(n324), .S(n1169), .Y(n322) );
  MUX2X1 U339 ( .B(n326), .A(n327), .S(n1181), .Y(n325) );
  MUX2X1 U340 ( .B(n329), .A(n330), .S(n1181), .Y(n328) );
  MUX2X1 U341 ( .B(n332), .A(n333), .S(n1181), .Y(n331) );
  MUX2X1 U342 ( .B(n335), .A(n336), .S(n1181), .Y(n334) );
  MUX2X1 U343 ( .B(n338), .A(n339), .S(n1169), .Y(n337) );
  MUX2X1 U344 ( .B(n341), .A(n342), .S(n1181), .Y(n340) );
  MUX2X1 U345 ( .B(n344), .A(n345), .S(n1181), .Y(n343) );
  MUX2X1 U346 ( .B(n347), .A(n348), .S(n1181), .Y(n346) );
  MUX2X1 U347 ( .B(n350), .A(n351), .S(n1181), .Y(n349) );
  MUX2X1 U348 ( .B(n353), .A(n354), .S(n1319), .Y(n352) );
  MUX2X1 U349 ( .B(n356), .A(n357), .S(n1181), .Y(n355) );
  MUX2X1 U350 ( .B(n359), .A(n360), .S(n1181), .Y(n358) );
  MUX2X1 U351 ( .B(n362), .A(n363), .S(n1181), .Y(n361) );
  MUX2X1 U352 ( .B(n365), .A(n366), .S(n1181), .Y(n364) );
  MUX2X1 U353 ( .B(n368), .A(n369), .S(n1319), .Y(n367) );
  MUX2X1 U354 ( .B(n371), .A(n372), .S(n1182), .Y(n370) );
  MUX2X1 U355 ( .B(n374), .A(n375), .S(n1182), .Y(n373) );
  MUX2X1 U356 ( .B(n377), .A(n378), .S(n1182), .Y(n376) );
  MUX2X1 U357 ( .B(n380), .A(n381), .S(n1182), .Y(n379) );
  MUX2X1 U358 ( .B(n383), .A(n384), .S(n1319), .Y(n382) );
  MUX2X1 U359 ( .B(n386), .A(n387), .S(n1182), .Y(n385) );
  MUX2X1 U360 ( .B(n389), .A(n390), .S(n1182), .Y(n388) );
  MUX2X1 U361 ( .B(n392), .A(n393), .S(n1182), .Y(n391) );
  MUX2X1 U362 ( .B(n395), .A(n396), .S(n1182), .Y(n394) );
  MUX2X1 U363 ( .B(n398), .A(n399), .S(n1319), .Y(n397) );
  MUX2X1 U364 ( .B(n401), .A(n402), .S(n1182), .Y(n400) );
  MUX2X1 U365 ( .B(n404), .A(n405), .S(n1182), .Y(n403) );
  MUX2X1 U366 ( .B(n407), .A(n408), .S(n1182), .Y(n406) );
  MUX2X1 U367 ( .B(n410), .A(n411), .S(n1182), .Y(n409) );
  MUX2X1 U368 ( .B(n413), .A(n414), .S(n1319), .Y(n412) );
  MUX2X1 U369 ( .B(n416), .A(n417), .S(n1183), .Y(n415) );
  MUX2X1 U370 ( .B(n419), .A(n420), .S(n1183), .Y(n418) );
  MUX2X1 U371 ( .B(n422), .A(n423), .S(n1183), .Y(n421) );
  MUX2X1 U372 ( .B(n425), .A(n426), .S(n1183), .Y(n424) );
  MUX2X1 U373 ( .B(n428), .A(n429), .S(n1319), .Y(n427) );
  MUX2X1 U374 ( .B(n431), .A(n432), .S(n1183), .Y(n430) );
  MUX2X1 U375 ( .B(n434), .A(n435), .S(n1183), .Y(n433) );
  MUX2X1 U376 ( .B(n437), .A(n438), .S(n1183), .Y(n436) );
  MUX2X1 U377 ( .B(n440), .A(n441), .S(n1183), .Y(n439) );
  MUX2X1 U378 ( .B(n443), .A(n444), .S(n1319), .Y(n442) );
  MUX2X1 U379 ( .B(n446), .A(n447), .S(n1183), .Y(n445) );
  MUX2X1 U380 ( .B(n449), .A(n450), .S(n1183), .Y(n448) );
  MUX2X1 U381 ( .B(n452), .A(n453), .S(n1183), .Y(n451) );
  MUX2X1 U382 ( .B(n455), .A(n456), .S(n1183), .Y(n454) );
  MUX2X1 U383 ( .B(n458), .A(n459), .S(n1319), .Y(n457) );
  MUX2X1 U384 ( .B(n461), .A(n462), .S(n1184), .Y(n460) );
  MUX2X1 U385 ( .B(n464), .A(n465), .S(n1184), .Y(n463) );
  MUX2X1 U386 ( .B(n467), .A(n468), .S(n1184), .Y(n466) );
  MUX2X1 U387 ( .B(n470), .A(n471), .S(n1184), .Y(n469) );
  MUX2X1 U388 ( .B(n473), .A(n474), .S(n1319), .Y(n472) );
  MUX2X1 U389 ( .B(n476), .A(n477), .S(n1184), .Y(n475) );
  MUX2X1 U390 ( .B(n479), .A(n480), .S(n1184), .Y(n478) );
  MUX2X1 U391 ( .B(n482), .A(n483), .S(n1184), .Y(n481) );
  MUX2X1 U392 ( .B(n485), .A(n486), .S(n1184), .Y(n484) );
  MUX2X1 U393 ( .B(n488), .A(n489), .S(n1319), .Y(n487) );
  MUX2X1 U394 ( .B(n491), .A(n492), .S(n1184), .Y(n490) );
  MUX2X1 U395 ( .B(n494), .A(n495), .S(n1184), .Y(n493) );
  MUX2X1 U396 ( .B(n497), .A(n498), .S(n1184), .Y(n496) );
  MUX2X1 U397 ( .B(n500), .A(n501), .S(n1184), .Y(n499) );
  MUX2X1 U398 ( .B(n503), .A(n504), .S(n1319), .Y(n502) );
  MUX2X1 U399 ( .B(n506), .A(n507), .S(n1185), .Y(n505) );
  MUX2X1 U400 ( .B(n509), .A(n510), .S(n1185), .Y(n508) );
  MUX2X1 U401 ( .B(n512), .A(n513), .S(n1185), .Y(n511) );
  MUX2X1 U402 ( .B(n515), .A(n516), .S(n1185), .Y(n514) );
  MUX2X1 U403 ( .B(n518), .A(n519), .S(n1319), .Y(n517) );
  MUX2X1 U404 ( .B(n521), .A(n522), .S(n1185), .Y(n520) );
  MUX2X1 U405 ( .B(n524), .A(n525), .S(n1185), .Y(n523) );
  MUX2X1 U406 ( .B(n527), .A(n528), .S(n1185), .Y(n526) );
  MUX2X1 U407 ( .B(n530), .A(n531), .S(n1185), .Y(n529) );
  MUX2X1 U408 ( .B(n533), .A(n534), .S(n1169), .Y(n532) );
  MUX2X1 U409 ( .B(n536), .A(n537), .S(n1185), .Y(n535) );
  MUX2X1 U410 ( .B(n539), .A(n540), .S(n1185), .Y(n538) );
  MUX2X1 U411 ( .B(n542), .A(n543), .S(n1185), .Y(n541) );
  MUX2X1 U412 ( .B(n545), .A(n546), .S(n1185), .Y(n544) );
  MUX2X1 U413 ( .B(n548), .A(n549), .S(n1169), .Y(n547) );
  MUX2X1 U414 ( .B(n551), .A(n552), .S(n1186), .Y(n550) );
  MUX2X1 U415 ( .B(n554), .A(n555), .S(n1186), .Y(n553) );
  MUX2X1 U416 ( .B(n557), .A(n558), .S(n1186), .Y(n556) );
  MUX2X1 U417 ( .B(n560), .A(n561), .S(n1186), .Y(n559) );
  MUX2X1 U418 ( .B(n563), .A(n564), .S(n1319), .Y(n562) );
  MUX2X1 U419 ( .B(n566), .A(n567), .S(n1186), .Y(n565) );
  MUX2X1 U420 ( .B(n569), .A(n570), .S(n1186), .Y(n568) );
  MUX2X1 U421 ( .B(n572), .A(n573), .S(n1186), .Y(n571) );
  MUX2X1 U422 ( .B(n575), .A(n576), .S(n1186), .Y(n574) );
  MUX2X1 U423 ( .B(n578), .A(n579), .S(n1169), .Y(n577) );
  MUX2X1 U424 ( .B(n581), .A(n582), .S(n1186), .Y(n580) );
  MUX2X1 U425 ( .B(n584), .A(n585), .S(n1186), .Y(n583) );
  MUX2X1 U426 ( .B(n587), .A(n588), .S(n1186), .Y(n586) );
  MUX2X1 U427 ( .B(n590), .A(n591), .S(n1186), .Y(n589) );
  MUX2X1 U428 ( .B(n593), .A(n594), .S(n1169), .Y(n592) );
  MUX2X1 U429 ( .B(n596), .A(n597), .S(n1187), .Y(n595) );
  MUX2X1 U430 ( .B(n599), .A(n600), .S(n1187), .Y(n598) );
  MUX2X1 U431 ( .B(n602), .A(n603), .S(n1187), .Y(n601) );
  MUX2X1 U432 ( .B(n605), .A(n606), .S(n1187), .Y(n604) );
  MUX2X1 U433 ( .B(n608), .A(n609), .S(n1169), .Y(n607) );
  MUX2X1 U434 ( .B(n611), .A(n612), .S(n1187), .Y(n610) );
  MUX2X1 U435 ( .B(n614), .A(n615), .S(n1187), .Y(n613) );
  MUX2X1 U436 ( .B(n617), .A(n618), .S(n1187), .Y(n616) );
  MUX2X1 U437 ( .B(n620), .A(n621), .S(n1187), .Y(n619) );
  MUX2X1 U438 ( .B(n623), .A(n624), .S(n1319), .Y(n622) );
  MUX2X1 U439 ( .B(n626), .A(n627), .S(n1187), .Y(n625) );
  MUX2X1 U440 ( .B(n629), .A(n630), .S(n1187), .Y(n628) );
  MUX2X1 U441 ( .B(n632), .A(n633), .S(n1187), .Y(n631) );
  MUX2X1 U442 ( .B(n635), .A(n636), .S(n1187), .Y(n634) );
  MUX2X1 U443 ( .B(n638), .A(n639), .S(n1319), .Y(n637) );
  MUX2X1 U444 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1193), .Y(n161) );
  MUX2X1 U445 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1193), .Y(n160) );
  MUX2X1 U446 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1193), .Y(n164) );
  MUX2X1 U447 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1193), .Y(n163) );
  MUX2X1 U448 ( .B(n162), .A(n159), .S(n1174), .Y(n173) );
  MUX2X1 U449 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1194), .Y(n167) );
  MUX2X1 U450 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1194), .Y(n166) );
  MUX2X1 U451 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1194), .Y(n170) );
  MUX2X1 U452 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1194), .Y(n169) );
  MUX2X1 U453 ( .B(n168), .A(n165), .S(n1174), .Y(n172) );
  MUX2X1 U454 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1194), .Y(n176) );
  MUX2X1 U455 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1194), .Y(n175) );
  MUX2X1 U456 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1194), .Y(n179) );
  MUX2X1 U457 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1194), .Y(n178) );
  MUX2X1 U458 ( .B(n177), .A(n174), .S(n1174), .Y(n188) );
  MUX2X1 U459 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1194), .Y(n182) );
  MUX2X1 U460 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1194), .Y(n181) );
  MUX2X1 U461 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1194), .Y(n185) );
  MUX2X1 U462 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1194), .Y(n184) );
  MUX2X1 U463 ( .B(n183), .A(n180), .S(n1174), .Y(n187) );
  MUX2X1 U464 ( .B(n186), .A(n171), .S(n1168), .Y(n640) );
  MUX2X1 U465 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1195), .Y(n191) );
  MUX2X1 U466 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1195), .Y(n190) );
  MUX2X1 U467 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1195), .Y(n194) );
  MUX2X1 U468 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1195), .Y(n193) );
  MUX2X1 U469 ( .B(n192), .A(n189), .S(n1174), .Y(n203) );
  MUX2X1 U470 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1195), .Y(n197) );
  MUX2X1 U471 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1195), .Y(n196) );
  MUX2X1 U472 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1195), .Y(n200) );
  MUX2X1 U473 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1195), .Y(n199) );
  MUX2X1 U474 ( .B(n198), .A(n195), .S(n1174), .Y(n202) );
  MUX2X1 U475 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1195), .Y(n206) );
  MUX2X1 U476 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1195), .Y(n205) );
  MUX2X1 U477 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1195), .Y(n209) );
  MUX2X1 U478 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1195), .Y(n208) );
  MUX2X1 U479 ( .B(n207), .A(n204), .S(n1174), .Y(n219) );
  MUX2X1 U480 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1196), .Y(n212) );
  MUX2X1 U481 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1196), .Y(n211) );
  MUX2X1 U482 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1196), .Y(n216) );
  MUX2X1 U483 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1196), .Y(n215) );
  MUX2X1 U484 ( .B(n213), .A(n210), .S(n1174), .Y(n218) );
  MUX2X1 U485 ( .B(n217), .A(n201), .S(n1168), .Y(n641) );
  MUX2X1 U486 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1196), .Y(n222) );
  MUX2X1 U487 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1196), .Y(n221) );
  MUX2X1 U488 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1196), .Y(n225) );
  MUX2X1 U489 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1196), .Y(n224) );
  MUX2X1 U490 ( .B(n223), .A(n220), .S(n1174), .Y(n234) );
  MUX2X1 U491 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1196), .Y(n228) );
  MUX2X1 U492 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1196), .Y(n227) );
  MUX2X1 U493 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1196), .Y(n231) );
  MUX2X1 U494 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1196), .Y(n230) );
  MUX2X1 U495 ( .B(n229), .A(n226), .S(n1174), .Y(n233) );
  MUX2X1 U496 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1197), .Y(n237) );
  MUX2X1 U497 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1197), .Y(n236) );
  MUX2X1 U498 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1197), .Y(n240) );
  MUX2X1 U499 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1197), .Y(n239) );
  MUX2X1 U500 ( .B(n238), .A(n235), .S(n1174), .Y(n249) );
  MUX2X1 U501 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1197), .Y(n243) );
  MUX2X1 U502 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1197), .Y(n242) );
  MUX2X1 U503 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1197), .Y(n246) );
  MUX2X1 U504 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1197), .Y(n245) );
  MUX2X1 U505 ( .B(n244), .A(n241), .S(n1174), .Y(n248) );
  MUX2X1 U506 ( .B(n247), .A(n232), .S(n1168), .Y(n642) );
  MUX2X1 U507 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1197), .Y(n252) );
  MUX2X1 U508 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1197), .Y(n251) );
  MUX2X1 U509 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1197), .Y(n255) );
  MUX2X1 U510 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1197), .Y(n254) );
  MUX2X1 U511 ( .B(n253), .A(n250), .S(n1173), .Y(n264) );
  MUX2X1 U512 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1198), .Y(n258) );
  MUX2X1 U513 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1198), .Y(n257) );
  MUX2X1 U514 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1198), .Y(n261) );
  MUX2X1 U515 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1198), .Y(n260) );
  MUX2X1 U516 ( .B(n259), .A(n256), .S(n1173), .Y(n263) );
  MUX2X1 U517 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1198), .Y(n267) );
  MUX2X1 U518 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1198), .Y(n266) );
  MUX2X1 U519 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1198), .Y(n270) );
  MUX2X1 U520 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1198), .Y(n269) );
  MUX2X1 U521 ( .B(n268), .A(n265), .S(n1173), .Y(n279) );
  MUX2X1 U522 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1198), .Y(n273) );
  MUX2X1 U523 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1198), .Y(n272) );
  MUX2X1 U524 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1198), .Y(n276) );
  MUX2X1 U525 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1198), .Y(n275) );
  MUX2X1 U526 ( .B(n274), .A(n271), .S(n1173), .Y(n278) );
  MUX2X1 U527 ( .B(n277), .A(n262), .S(n1168), .Y(n643) );
  MUX2X1 U528 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1199), .Y(n282) );
  MUX2X1 U529 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1199), .Y(n281) );
  MUX2X1 U530 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1199), .Y(n285) );
  MUX2X1 U531 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1199), .Y(n284) );
  MUX2X1 U532 ( .B(n283), .A(n280), .S(n1173), .Y(n294) );
  MUX2X1 U533 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1199), .Y(n288) );
  MUX2X1 U534 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1199), .Y(n287) );
  MUX2X1 U535 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1199), .Y(n291) );
  MUX2X1 U536 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1199), .Y(n290) );
  MUX2X1 U537 ( .B(n289), .A(n286), .S(n1173), .Y(n293) );
  MUX2X1 U538 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1199), .Y(n297) );
  MUX2X1 U539 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1199), .Y(n296) );
  MUX2X1 U540 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1199), .Y(n300) );
  MUX2X1 U541 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1199), .Y(n299) );
  MUX2X1 U542 ( .B(n298), .A(n295), .S(n1173), .Y(n309) );
  MUX2X1 U543 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1200), .Y(n303) );
  MUX2X1 U544 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1200), .Y(n302) );
  MUX2X1 U545 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1200), .Y(n306) );
  MUX2X1 U546 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1200), .Y(n305) );
  MUX2X1 U547 ( .B(n304), .A(n301), .S(n1173), .Y(n308) );
  MUX2X1 U548 ( .B(n307), .A(n292), .S(n1168), .Y(n644) );
  MUX2X1 U549 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1200), .Y(n312) );
  MUX2X1 U550 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1200), .Y(n311) );
  MUX2X1 U551 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1200), .Y(n315) );
  MUX2X1 U552 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1200), .Y(n314) );
  MUX2X1 U553 ( .B(n313), .A(n310), .S(n1173), .Y(n324) );
  MUX2X1 U554 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1200), .Y(n318) );
  MUX2X1 U555 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1200), .Y(n317) );
  MUX2X1 U556 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1200), .Y(n321) );
  MUX2X1 U557 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1200), .Y(n320) );
  MUX2X1 U558 ( .B(n319), .A(n316), .S(n1173), .Y(n323) );
  MUX2X1 U559 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1201), .Y(n327) );
  MUX2X1 U560 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1201), .Y(n326) );
  MUX2X1 U561 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1201), .Y(n330) );
  MUX2X1 U562 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1201), .Y(n329) );
  MUX2X1 U563 ( .B(n328), .A(n325), .S(n1173), .Y(n339) );
  MUX2X1 U564 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1201), .Y(n333) );
  MUX2X1 U565 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1201), .Y(n332) );
  MUX2X1 U566 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1201), .Y(n336) );
  MUX2X1 U567 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1201), .Y(n335) );
  MUX2X1 U568 ( .B(n334), .A(n331), .S(n1173), .Y(n338) );
  MUX2X1 U569 ( .B(n337), .A(n322), .S(n1168), .Y(n645) );
  MUX2X1 U570 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1201), .Y(n342) );
  MUX2X1 U571 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1201), .Y(n341) );
  MUX2X1 U572 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1201), .Y(n345) );
  MUX2X1 U573 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1201), .Y(n344) );
  MUX2X1 U574 ( .B(n343), .A(n340), .S(n1172), .Y(n354) );
  MUX2X1 U575 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1202), .Y(n348) );
  MUX2X1 U576 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1202), .Y(n347) );
  MUX2X1 U577 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1202), .Y(n351) );
  MUX2X1 U578 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1202), .Y(n350) );
  MUX2X1 U579 ( .B(n349), .A(n346), .S(n1172), .Y(n353) );
  MUX2X1 U580 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1202), .Y(n357) );
  MUX2X1 U581 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1202), .Y(n356) );
  MUX2X1 U582 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1202), .Y(n360) );
  MUX2X1 U583 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1202), .Y(n359) );
  MUX2X1 U584 ( .B(n358), .A(n355), .S(n1172), .Y(n369) );
  MUX2X1 U585 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1202), .Y(n363) );
  MUX2X1 U586 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1202), .Y(n362) );
  MUX2X1 U587 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1202), .Y(n366) );
  MUX2X1 U588 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1202), .Y(n365) );
  MUX2X1 U589 ( .B(n364), .A(n361), .S(n1172), .Y(n368) );
  MUX2X1 U590 ( .B(n367), .A(n352), .S(n1168), .Y(n646) );
  MUX2X1 U591 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1203), .Y(n372) );
  MUX2X1 U592 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1203), .Y(n371) );
  MUX2X1 U593 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1203), .Y(n375) );
  MUX2X1 U594 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1203), .Y(n374) );
  MUX2X1 U595 ( .B(n373), .A(n370), .S(n1172), .Y(n384) );
  MUX2X1 U596 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1203), .Y(n378) );
  MUX2X1 U597 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1203), .Y(n377) );
  MUX2X1 U598 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1203), .Y(n381) );
  MUX2X1 U599 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1203), .Y(n380) );
  MUX2X1 U600 ( .B(n379), .A(n376), .S(n1172), .Y(n383) );
  MUX2X1 U601 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1203), .Y(n387) );
  MUX2X1 U602 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1203), .Y(n386) );
  MUX2X1 U603 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1203), .Y(n390) );
  MUX2X1 U604 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1203), .Y(n389) );
  MUX2X1 U605 ( .B(n388), .A(n385), .S(n1172), .Y(n399) );
  MUX2X1 U606 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1204), .Y(n393) );
  MUX2X1 U607 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1204), .Y(n392) );
  MUX2X1 U608 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1204), .Y(n396) );
  MUX2X1 U609 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1204), .Y(n395) );
  MUX2X1 U610 ( .B(n394), .A(n391), .S(n1172), .Y(n398) );
  MUX2X1 U611 ( .B(n397), .A(n382), .S(n1168), .Y(n647) );
  MUX2X1 U612 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1204), .Y(n402) );
  MUX2X1 U613 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1204), .Y(n401) );
  MUX2X1 U614 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1204), .Y(n405) );
  MUX2X1 U615 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1204), .Y(n404) );
  MUX2X1 U616 ( .B(n403), .A(n400), .S(n1172), .Y(n414) );
  MUX2X1 U617 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1204), .Y(n408) );
  MUX2X1 U618 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1204), .Y(n407) );
  MUX2X1 U619 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1204), .Y(n411) );
  MUX2X1 U620 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1204), .Y(n410) );
  MUX2X1 U621 ( .B(n409), .A(n406), .S(n1172), .Y(n413) );
  MUX2X1 U622 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1205), .Y(n417) );
  MUX2X1 U623 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1205), .Y(n416) );
  MUX2X1 U624 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1205), .Y(n420) );
  MUX2X1 U625 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1205), .Y(n419) );
  MUX2X1 U626 ( .B(n418), .A(n415), .S(n1172), .Y(n429) );
  MUX2X1 U627 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1205), .Y(n423) );
  MUX2X1 U628 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1205), .Y(n422) );
  MUX2X1 U629 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1205), .Y(n426) );
  MUX2X1 U630 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1205), .Y(n425) );
  MUX2X1 U631 ( .B(n424), .A(n421), .S(n1172), .Y(n428) );
  MUX2X1 U632 ( .B(n427), .A(n412), .S(n1168), .Y(n648) );
  MUX2X1 U633 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1205), .Y(n432) );
  MUX2X1 U634 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1205), .Y(n431) );
  MUX2X1 U635 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1205), .Y(n435) );
  MUX2X1 U636 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1205), .Y(n434) );
  MUX2X1 U637 ( .B(n433), .A(n430), .S(n1171), .Y(n444) );
  MUX2X1 U638 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1206), .Y(n438) );
  MUX2X1 U639 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1206), .Y(n437) );
  MUX2X1 U640 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1206), .Y(n441) );
  MUX2X1 U641 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1206), .Y(n440) );
  MUX2X1 U642 ( .B(n439), .A(n436), .S(n1171), .Y(n443) );
  MUX2X1 U643 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1206), .Y(n447) );
  MUX2X1 U644 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1206), .Y(n446) );
  MUX2X1 U645 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1206), .Y(n450) );
  MUX2X1 U646 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1206), .Y(n449) );
  MUX2X1 U647 ( .B(n448), .A(n445), .S(n1171), .Y(n459) );
  MUX2X1 U648 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1206), .Y(n453) );
  MUX2X1 U649 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1206), .Y(n452) );
  MUX2X1 U650 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1206), .Y(n456) );
  MUX2X1 U651 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1206), .Y(n455) );
  MUX2X1 U652 ( .B(n454), .A(n451), .S(n1171), .Y(n458) );
  MUX2X1 U653 ( .B(n457), .A(n442), .S(n1168), .Y(n649) );
  MUX2X1 U654 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1207), .Y(n462) );
  MUX2X1 U655 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1207), .Y(n461) );
  MUX2X1 U656 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1207), .Y(n465) );
  MUX2X1 U657 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1207), .Y(n464) );
  MUX2X1 U658 ( .B(n463), .A(n460), .S(n1171), .Y(n474) );
  MUX2X1 U659 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1207), .Y(n468) );
  MUX2X1 U660 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1207), .Y(n467) );
  MUX2X1 U661 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1207), .Y(n471) );
  MUX2X1 U662 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1207), .Y(n470) );
  MUX2X1 U663 ( .B(n469), .A(n466), .S(n1171), .Y(n473) );
  MUX2X1 U664 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1207), .Y(n477) );
  MUX2X1 U665 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1207), .Y(n476) );
  MUX2X1 U666 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1207), .Y(n480) );
  MUX2X1 U667 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1207), .Y(n479) );
  MUX2X1 U668 ( .B(n478), .A(n475), .S(n1171), .Y(n489) );
  MUX2X1 U669 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1208), .Y(n483) );
  MUX2X1 U670 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1208), .Y(n482) );
  MUX2X1 U671 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1208), .Y(n486) );
  MUX2X1 U672 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1208), .Y(n485) );
  MUX2X1 U673 ( .B(n484), .A(n481), .S(n1171), .Y(n488) );
  MUX2X1 U674 ( .B(n487), .A(n472), .S(n1168), .Y(n650) );
  MUX2X1 U675 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1208), .Y(n492) );
  MUX2X1 U676 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1208), .Y(n491) );
  MUX2X1 U677 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1208), .Y(n495) );
  MUX2X1 U678 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1208), .Y(n494) );
  MUX2X1 U679 ( .B(n493), .A(n490), .S(n1171), .Y(n504) );
  MUX2X1 U680 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1208), .Y(n498) );
  MUX2X1 U681 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1208), .Y(n497) );
  MUX2X1 U682 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1208), .Y(n501) );
  MUX2X1 U683 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1208), .Y(n500) );
  MUX2X1 U684 ( .B(n499), .A(n496), .S(n1171), .Y(n503) );
  MUX2X1 U685 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1209), .Y(n507) );
  MUX2X1 U686 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1209), .Y(n506) );
  MUX2X1 U687 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1209), .Y(n510) );
  MUX2X1 U688 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1209), .Y(n509) );
  MUX2X1 U689 ( .B(n508), .A(n505), .S(n1171), .Y(n519) );
  MUX2X1 U690 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1209), .Y(n513) );
  MUX2X1 U691 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1209), .Y(n512) );
  MUX2X1 U692 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1209), .Y(n516) );
  MUX2X1 U693 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1209), .Y(n515) );
  MUX2X1 U694 ( .B(n514), .A(n511), .S(n1171), .Y(n518) );
  MUX2X1 U695 ( .B(n517), .A(n502), .S(n1168), .Y(n1163) );
  MUX2X1 U696 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1209), .Y(n522) );
  MUX2X1 U697 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1209), .Y(n521) );
  MUX2X1 U698 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1209), .Y(n525) );
  MUX2X1 U699 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1209), .Y(n524) );
  MUX2X1 U700 ( .B(n523), .A(n520), .S(n1170), .Y(n534) );
  MUX2X1 U701 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1210), .Y(n528) );
  MUX2X1 U702 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1210), .Y(n527) );
  MUX2X1 U703 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1210), .Y(n531) );
  MUX2X1 U704 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1210), .Y(n530) );
  MUX2X1 U705 ( .B(n529), .A(n526), .S(n1170), .Y(n533) );
  MUX2X1 U706 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1210), .Y(n537) );
  MUX2X1 U707 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1210), .Y(n536) );
  MUX2X1 U708 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1210), .Y(n540) );
  MUX2X1 U709 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1210), .Y(n539) );
  MUX2X1 U710 ( .B(n538), .A(n535), .S(n1170), .Y(n549) );
  MUX2X1 U711 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1210), .Y(n543) );
  MUX2X1 U712 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1210), .Y(n542) );
  MUX2X1 U713 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1210), .Y(n546) );
  MUX2X1 U714 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1210), .Y(n545) );
  MUX2X1 U715 ( .B(n544), .A(n541), .S(n1170), .Y(n548) );
  MUX2X1 U716 ( .B(n547), .A(n532), .S(n1168), .Y(n1164) );
  MUX2X1 U717 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1211), .Y(n552) );
  MUX2X1 U718 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1211), .Y(n551) );
  MUX2X1 U719 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1211), .Y(n555) );
  MUX2X1 U720 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1211), .Y(n554) );
  MUX2X1 U721 ( .B(n553), .A(n550), .S(n1170), .Y(n564) );
  MUX2X1 U722 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1211), .Y(n558) );
  MUX2X1 U723 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1211), .Y(n557) );
  MUX2X1 U724 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1211), .Y(n561) );
  MUX2X1 U725 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1211), .Y(n560) );
  MUX2X1 U726 ( .B(n559), .A(n556), .S(n1170), .Y(n563) );
  MUX2X1 U727 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1211), .Y(n567) );
  MUX2X1 U728 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1211), .Y(n566) );
  MUX2X1 U729 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1211), .Y(n570) );
  MUX2X1 U730 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1211), .Y(n569) );
  MUX2X1 U731 ( .B(n568), .A(n565), .S(n1170), .Y(n579) );
  MUX2X1 U732 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1212), .Y(n573) );
  MUX2X1 U733 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1212), .Y(n572) );
  MUX2X1 U734 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1212), .Y(n576) );
  MUX2X1 U735 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1212), .Y(n575) );
  MUX2X1 U736 ( .B(n574), .A(n571), .S(n1170), .Y(n578) );
  MUX2X1 U737 ( .B(n577), .A(n562), .S(n1168), .Y(n1165) );
  MUX2X1 U738 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1212), .Y(n582) );
  MUX2X1 U739 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1212), .Y(n581) );
  MUX2X1 U740 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1212), .Y(n585) );
  MUX2X1 U741 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1212), .Y(n584) );
  MUX2X1 U742 ( .B(n583), .A(n580), .S(n1170), .Y(n594) );
  MUX2X1 U743 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1212), .Y(n588) );
  MUX2X1 U744 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1212), .Y(n587) );
  MUX2X1 U745 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1212), .Y(n591) );
  MUX2X1 U746 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1212), .Y(n590) );
  MUX2X1 U747 ( .B(n589), .A(n586), .S(n1170), .Y(n593) );
  MUX2X1 U748 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1213), .Y(n597) );
  MUX2X1 U749 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1213), .Y(n596) );
  MUX2X1 U750 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1213), .Y(n600) );
  MUX2X1 U751 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1213), .Y(n599) );
  MUX2X1 U752 ( .B(n598), .A(n595), .S(n1170), .Y(n609) );
  MUX2X1 U753 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1213), .Y(n603) );
  MUX2X1 U754 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1213), .Y(n602) );
  MUX2X1 U755 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1213), .Y(n606) );
  MUX2X1 U756 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1213), .Y(n605) );
  MUX2X1 U757 ( .B(n604), .A(n601), .S(n1170), .Y(n608) );
  MUX2X1 U758 ( .B(n607), .A(n592), .S(n1168), .Y(n1166) );
  MUX2X1 U759 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1213), .Y(n612) );
  MUX2X1 U760 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1213), .Y(n611) );
  MUX2X1 U761 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1213), .Y(n615) );
  MUX2X1 U762 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1213), .Y(n614) );
  MUX2X1 U763 ( .B(n613), .A(n610), .S(n1170), .Y(n624) );
  MUX2X1 U764 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1193), .Y(n618) );
  MUX2X1 U765 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1215), .Y(n617) );
  MUX2X1 U766 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1215), .Y(n621) );
  MUX2X1 U767 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1215), .Y(n620) );
  MUX2X1 U768 ( .B(n619), .A(n616), .S(n1171), .Y(n623) );
  MUX2X1 U769 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1193), .Y(n627) );
  MUX2X1 U770 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1211), .Y(n626) );
  MUX2X1 U771 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1193), .Y(n630) );
  MUX2X1 U772 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1193), .Y(n629) );
  MUX2X1 U773 ( .B(n628), .A(n625), .S(n1170), .Y(n639) );
  MUX2X1 U774 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1213), .Y(n633) );
  MUX2X1 U775 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1193), .Y(n632) );
  MUX2X1 U776 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1212), .Y(n636) );
  MUX2X1 U777 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1212), .Y(n635) );
  MUX2X1 U778 ( .B(n634), .A(n631), .S(n1171), .Y(n638) );
  MUX2X1 U779 ( .B(n637), .A(n622), .S(n1168), .Y(n1167) );
  INVX8 U780 ( .A(n1192), .Y(n1193) );
  INVX8 U781 ( .A(n1192), .Y(n1194) );
  INVX8 U782 ( .A(n1192), .Y(n1195) );
  INVX8 U783 ( .A(n1191), .Y(n1196) );
  INVX8 U784 ( .A(n1191), .Y(n1197) );
  INVX8 U785 ( .A(n1191), .Y(n1198) );
  INVX8 U786 ( .A(n1192), .Y(n1199) );
  INVX8 U787 ( .A(n1191), .Y(n1200) );
  INVX8 U788 ( .A(n1191), .Y(n1201) );
  INVX8 U789 ( .A(n1190), .Y(n1202) );
  INVX8 U790 ( .A(n1190), .Y(n1203) );
  INVX8 U791 ( .A(n1190), .Y(n1204) );
  INVX8 U792 ( .A(n1189), .Y(n1205) );
  INVX8 U793 ( .A(n1189), .Y(n1206) );
  INVX8 U794 ( .A(n1189), .Y(n1207) );
  INVX8 U795 ( .A(n1190), .Y(n1208) );
  INVX8 U796 ( .A(n1189), .Y(n1209) );
  INVX8 U797 ( .A(n1189), .Y(n1210) );
  INVX8 U798 ( .A(n1192), .Y(n1211) );
  INVX8 U799 ( .A(n1190), .Y(n1213) );
  INVX1 U800 ( .A(N11), .Y(n1316) );
  INVX1 U801 ( .A(N10), .Y(n1314) );
  INVX8 U802 ( .A(n1280), .Y(n1278) );
  INVX8 U803 ( .A(n1280), .Y(n1279) );
  INVX8 U804 ( .A(n89), .Y(n1281) );
  INVX8 U805 ( .A(n89), .Y(n1282) );
  INVX8 U806 ( .A(n90), .Y(n1283) );
  INVX8 U807 ( .A(n90), .Y(n1284) );
  INVX8 U808 ( .A(n91), .Y(n1285) );
  INVX8 U809 ( .A(n91), .Y(n1286) );
  INVX8 U810 ( .A(n92), .Y(n1287) );
  INVX8 U811 ( .A(n92), .Y(n1288) );
  INVX8 U812 ( .A(n93), .Y(n1289) );
  INVX8 U813 ( .A(n93), .Y(n1290) );
  INVX8 U814 ( .A(n94), .Y(n1291) );
  INVX8 U815 ( .A(n94), .Y(n1292) );
  INVX8 U816 ( .A(n95), .Y(n1293) );
  INVX8 U817 ( .A(n95), .Y(n1294) );
  INVX8 U818 ( .A(n5), .Y(n1295) );
  INVX8 U819 ( .A(n5), .Y(n1296) );
  INVX8 U820 ( .A(n96), .Y(n1297) );
  INVX8 U821 ( .A(n96), .Y(n1298) );
  INVX8 U822 ( .A(n97), .Y(n1299) );
  INVX8 U823 ( .A(n97), .Y(n1300) );
  INVX8 U824 ( .A(n98), .Y(n1301) );
  INVX8 U825 ( .A(n98), .Y(n1302) );
  INVX8 U826 ( .A(n6), .Y(n1303) );
  INVX8 U827 ( .A(n6), .Y(n1304) );
  INVX8 U828 ( .A(n7), .Y(n1305) );
  INVX8 U829 ( .A(n8), .Y(n1306) );
  INVX8 U830 ( .A(n8), .Y(n1307) );
  INVX8 U831 ( .A(n9), .Y(n1308) );
  INVX8 U832 ( .A(n9), .Y(n1309) );
  INVX8 U833 ( .A(n10), .Y(n1310) );
  INVX8 U834 ( .A(n10), .Y(n1311) );
  AND2X2 U835 ( .A(n75), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U836 ( .A(n75), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U837 ( .A(n75), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U838 ( .A(n1), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U839 ( .A(n75), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U840 ( .A(n75), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U841 ( .A(n75), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U842 ( .A(n75), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U843 ( .A(n75), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U844 ( .A(n75), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U845 ( .A(n1), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U846 ( .A(n1), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U847 ( .A(n1), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U848 ( .A(n1), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U849 ( .A(n1), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U850 ( .A(\mem<31><0> ), .B(n4), .Y(n1323) );
  OAI21X1 U851 ( .A(n1219), .B(n1281), .C(n1323), .Y(n2361) );
  NAND2X1 U852 ( .A(\mem<31><1> ), .B(n4), .Y(n1324) );
  OAI21X1 U853 ( .A(n1284), .B(n1218), .C(n1324), .Y(n2360) );
  NAND2X1 U854 ( .A(\mem<31><2> ), .B(n4), .Y(n1325) );
  OAI21X1 U855 ( .A(n1286), .B(n1218), .C(n1325), .Y(n2359) );
  NAND2X1 U856 ( .A(\mem<31><3> ), .B(n4), .Y(n1326) );
  OAI21X1 U857 ( .A(n1288), .B(n1218), .C(n1326), .Y(n2358) );
  NAND2X1 U858 ( .A(\mem<31><4> ), .B(n4), .Y(n1327) );
  OAI21X1 U859 ( .A(n1290), .B(n1218), .C(n1327), .Y(n2357) );
  NAND2X1 U860 ( .A(\mem<31><5> ), .B(n4), .Y(n1328) );
  OAI21X1 U861 ( .A(n1292), .B(n1218), .C(n1328), .Y(n2356) );
  NAND2X1 U862 ( .A(\mem<31><6> ), .B(n4), .Y(n1329) );
  OAI21X1 U863 ( .A(n1294), .B(n1218), .C(n1329), .Y(n2355) );
  NAND2X1 U864 ( .A(\mem<31><7> ), .B(n4), .Y(n1330) );
  OAI21X1 U865 ( .A(n1296), .B(n1218), .C(n1330), .Y(n2354) );
  NAND2X1 U866 ( .A(\mem<31><8> ), .B(n4), .Y(n1331) );
  OAI21X1 U867 ( .A(n1298), .B(n1218), .C(n1331), .Y(n2353) );
  NAND2X1 U868 ( .A(\mem<31><9> ), .B(n4), .Y(n1332) );
  OAI21X1 U869 ( .A(n1300), .B(n1219), .C(n1332), .Y(n2352) );
  NAND2X1 U870 ( .A(\mem<31><10> ), .B(n4), .Y(n1333) );
  OAI21X1 U871 ( .A(n1302), .B(n1219), .C(n1333), .Y(n2351) );
  NAND2X1 U872 ( .A(\mem<31><11> ), .B(n4), .Y(n1334) );
  OAI21X1 U873 ( .A(n1304), .B(n1219), .C(n1334), .Y(n2350) );
  NAND2X1 U874 ( .A(\mem<31><12> ), .B(n4), .Y(n1335) );
  OAI21X1 U875 ( .A(n1305), .B(n1219), .C(n1335), .Y(n2349) );
  NAND2X1 U876 ( .A(\mem<31><13> ), .B(n4), .Y(n1336) );
  OAI21X1 U877 ( .A(n1307), .B(n1219), .C(n1336), .Y(n2348) );
  NAND2X1 U878 ( .A(\mem<31><14> ), .B(n4), .Y(n1337) );
  OAI21X1 U879 ( .A(n1309), .B(n1219), .C(n1337), .Y(n2347) );
  NAND2X1 U880 ( .A(\mem<31><15> ), .B(n4), .Y(n1338) );
  OAI21X1 U881 ( .A(n1311), .B(n1219), .C(n1338), .Y(n2346) );
  NAND2X1 U882 ( .A(\mem<30><0> ), .B(n12), .Y(n1339) );
  OAI21X1 U883 ( .A(n1220), .B(n1281), .C(n1339), .Y(n2345) );
  NAND2X1 U884 ( .A(\mem<30><1> ), .B(n12), .Y(n1340) );
  OAI21X1 U885 ( .A(n1220), .B(n1283), .C(n1340), .Y(n2344) );
  NAND2X1 U886 ( .A(\mem<30><2> ), .B(n12), .Y(n1341) );
  OAI21X1 U887 ( .A(n1220), .B(n1286), .C(n1341), .Y(n2343) );
  NAND2X1 U888 ( .A(\mem<30><3> ), .B(n12), .Y(n1342) );
  OAI21X1 U889 ( .A(n1220), .B(n1287), .C(n1342), .Y(n2342) );
  NAND2X1 U890 ( .A(\mem<30><4> ), .B(n12), .Y(n1343) );
  OAI21X1 U891 ( .A(n1220), .B(n1290), .C(n1343), .Y(n2341) );
  NAND2X1 U892 ( .A(\mem<30><5> ), .B(n12), .Y(n1344) );
  OAI21X1 U893 ( .A(n1220), .B(n1291), .C(n1344), .Y(n2340) );
  NAND2X1 U894 ( .A(\mem<30><6> ), .B(n12), .Y(n1345) );
  OAI21X1 U895 ( .A(n1220), .B(n1294), .C(n1345), .Y(n2339) );
  NAND2X1 U896 ( .A(\mem<30><7> ), .B(n12), .Y(n1346) );
  OAI21X1 U897 ( .A(n1220), .B(n1295), .C(n1346), .Y(n2338) );
  NAND2X1 U898 ( .A(\mem<30><8> ), .B(n12), .Y(n1347) );
  OAI21X1 U899 ( .A(n1221), .B(n1298), .C(n1347), .Y(n2337) );
  NAND2X1 U900 ( .A(\mem<30><9> ), .B(n12), .Y(n1348) );
  OAI21X1 U901 ( .A(n1221), .B(n1299), .C(n1348), .Y(n2336) );
  NAND2X1 U902 ( .A(\mem<30><10> ), .B(n12), .Y(n1349) );
  OAI21X1 U903 ( .A(n1221), .B(n1302), .C(n1349), .Y(n2335) );
  NAND2X1 U904 ( .A(\mem<30><11> ), .B(n12), .Y(n1350) );
  OAI21X1 U905 ( .A(n1221), .B(n1303), .C(n1350), .Y(n2334) );
  NAND2X1 U906 ( .A(\mem<30><12> ), .B(n12), .Y(n1351) );
  OAI21X1 U907 ( .A(n1221), .B(n1305), .C(n1351), .Y(n2333) );
  NAND2X1 U908 ( .A(\mem<30><13> ), .B(n12), .Y(n1352) );
  OAI21X1 U909 ( .A(n1221), .B(n1306), .C(n1352), .Y(n2332) );
  NAND2X1 U910 ( .A(\mem<30><14> ), .B(n12), .Y(n1353) );
  OAI21X1 U911 ( .A(n1221), .B(n1308), .C(n1353), .Y(n2331) );
  NAND2X1 U912 ( .A(\mem<30><15> ), .B(n12), .Y(n1354) );
  OAI21X1 U913 ( .A(n1221), .B(n1310), .C(n1354), .Y(n2330) );
  NAND3X1 U914 ( .A(n1313), .B(n1317), .C(n1316), .Y(n1355) );
  NAND2X1 U915 ( .A(\mem<29><0> ), .B(n14), .Y(n1356) );
  OAI21X1 U916 ( .A(n1222), .B(n1281), .C(n1356), .Y(n2329) );
  NAND2X1 U917 ( .A(\mem<29><1> ), .B(n14), .Y(n1357) );
  OAI21X1 U918 ( .A(n1222), .B(n1284), .C(n1357), .Y(n2328) );
  NAND2X1 U919 ( .A(\mem<29><2> ), .B(n14), .Y(n1358) );
  OAI21X1 U920 ( .A(n1222), .B(n1285), .C(n1358), .Y(n2327) );
  NAND2X1 U921 ( .A(\mem<29><3> ), .B(n14), .Y(n1359) );
  OAI21X1 U922 ( .A(n1222), .B(n1288), .C(n1359), .Y(n2326) );
  NAND2X1 U923 ( .A(\mem<29><4> ), .B(n14), .Y(n1360) );
  OAI21X1 U924 ( .A(n1222), .B(n1289), .C(n1360), .Y(n2325) );
  NAND2X1 U925 ( .A(\mem<29><5> ), .B(n14), .Y(n1361) );
  OAI21X1 U926 ( .A(n1222), .B(n1292), .C(n1361), .Y(n2324) );
  NAND2X1 U927 ( .A(\mem<29><6> ), .B(n14), .Y(n1362) );
  OAI21X1 U928 ( .A(n1222), .B(n1293), .C(n1362), .Y(n2323) );
  NAND2X1 U929 ( .A(\mem<29><7> ), .B(n14), .Y(n1363) );
  OAI21X1 U930 ( .A(n1222), .B(n1296), .C(n1363), .Y(n2322) );
  NAND2X1 U931 ( .A(\mem<29><8> ), .B(n14), .Y(n1364) );
  OAI21X1 U932 ( .A(n1223), .B(n1297), .C(n1364), .Y(n2321) );
  NAND2X1 U933 ( .A(\mem<29><9> ), .B(n14), .Y(n1365) );
  OAI21X1 U934 ( .A(n1223), .B(n1300), .C(n1365), .Y(n2320) );
  NAND2X1 U935 ( .A(\mem<29><10> ), .B(n14), .Y(n1366) );
  OAI21X1 U936 ( .A(n1223), .B(n1301), .C(n1366), .Y(n2319) );
  NAND2X1 U937 ( .A(\mem<29><11> ), .B(n14), .Y(n1367) );
  OAI21X1 U938 ( .A(n1223), .B(n1304), .C(n1367), .Y(n2318) );
  NAND2X1 U939 ( .A(\mem<29><12> ), .B(n14), .Y(n1368) );
  OAI21X1 U940 ( .A(n1223), .B(n1305), .C(n1368), .Y(n2317) );
  NAND2X1 U941 ( .A(\mem<29><13> ), .B(n14), .Y(n1369) );
  OAI21X1 U942 ( .A(n1223), .B(n1307), .C(n1369), .Y(n2316) );
  NAND2X1 U943 ( .A(\mem<29><14> ), .B(n14), .Y(n1370) );
  OAI21X1 U944 ( .A(n1223), .B(n1309), .C(n1370), .Y(n2315) );
  NAND2X1 U945 ( .A(\mem<29><15> ), .B(n14), .Y(n1371) );
  OAI21X1 U946 ( .A(n1223), .B(n1311), .C(n1371), .Y(n2314) );
  NAND3X1 U947 ( .A(n1317), .B(n1316), .C(n1314), .Y(n1372) );
  NAND2X1 U948 ( .A(\mem<28><0> ), .B(n16), .Y(n1373) );
  OAI21X1 U949 ( .A(n1224), .B(n1281), .C(n1373), .Y(n2313) );
  NAND2X1 U950 ( .A(\mem<28><1> ), .B(n16), .Y(n1374) );
  OAI21X1 U951 ( .A(n1224), .B(n1283), .C(n1374), .Y(n2312) );
  NAND2X1 U952 ( .A(\mem<28><2> ), .B(n16), .Y(n1375) );
  OAI21X1 U953 ( .A(n1224), .B(n1286), .C(n1375), .Y(n2311) );
  NAND2X1 U954 ( .A(\mem<28><3> ), .B(n16), .Y(n1376) );
  OAI21X1 U955 ( .A(n1224), .B(n1287), .C(n1376), .Y(n2310) );
  NAND2X1 U956 ( .A(\mem<28><4> ), .B(n16), .Y(n1377) );
  OAI21X1 U957 ( .A(n1224), .B(n1290), .C(n1377), .Y(n2309) );
  NAND2X1 U958 ( .A(\mem<28><5> ), .B(n16), .Y(n1378) );
  OAI21X1 U959 ( .A(n1224), .B(n1291), .C(n1378), .Y(n2308) );
  NAND2X1 U960 ( .A(\mem<28><6> ), .B(n16), .Y(n1379) );
  OAI21X1 U961 ( .A(n1224), .B(n1294), .C(n1379), .Y(n2307) );
  NAND2X1 U962 ( .A(\mem<28><7> ), .B(n16), .Y(n1380) );
  OAI21X1 U963 ( .A(n1224), .B(n1295), .C(n1380), .Y(n2306) );
  NAND2X1 U964 ( .A(\mem<28><8> ), .B(n16), .Y(n1381) );
  OAI21X1 U965 ( .A(n1225), .B(n1298), .C(n1381), .Y(n2305) );
  NAND2X1 U966 ( .A(\mem<28><9> ), .B(n16), .Y(n1382) );
  OAI21X1 U967 ( .A(n1225), .B(n1299), .C(n1382), .Y(n2304) );
  NAND2X1 U968 ( .A(\mem<28><10> ), .B(n16), .Y(n1383) );
  OAI21X1 U969 ( .A(n1225), .B(n1302), .C(n1383), .Y(n2303) );
  NAND2X1 U970 ( .A(\mem<28><11> ), .B(n16), .Y(n1384) );
  OAI21X1 U971 ( .A(n1225), .B(n1303), .C(n1384), .Y(n2302) );
  NAND2X1 U972 ( .A(\mem<28><12> ), .B(n16), .Y(n1385) );
  OAI21X1 U973 ( .A(n1225), .B(n1305), .C(n1385), .Y(n2301) );
  NAND2X1 U974 ( .A(\mem<28><13> ), .B(n16), .Y(n1386) );
  OAI21X1 U975 ( .A(n1225), .B(n1306), .C(n1386), .Y(n2300) );
  NAND2X1 U976 ( .A(\mem<28><14> ), .B(n16), .Y(n1387) );
  OAI21X1 U977 ( .A(n1225), .B(n1308), .C(n1387), .Y(n2299) );
  NAND2X1 U978 ( .A(\mem<28><15> ), .B(n16), .Y(n1388) );
  OAI21X1 U979 ( .A(n1225), .B(n1310), .C(n1388), .Y(n2298) );
  NAND3X1 U980 ( .A(n1313), .B(n1315), .C(n1318), .Y(n1389) );
  NAND2X1 U981 ( .A(\mem<27><0> ), .B(n18), .Y(n1390) );
  OAI21X1 U982 ( .A(n1226), .B(n1281), .C(n1390), .Y(n2297) );
  NAND2X1 U983 ( .A(\mem<27><1> ), .B(n18), .Y(n1391) );
  OAI21X1 U984 ( .A(n1226), .B(n1284), .C(n1391), .Y(n2296) );
  NAND2X1 U985 ( .A(\mem<27><2> ), .B(n18), .Y(n1392) );
  OAI21X1 U986 ( .A(n1226), .B(n1285), .C(n1392), .Y(n2295) );
  NAND2X1 U987 ( .A(\mem<27><3> ), .B(n18), .Y(n1393) );
  OAI21X1 U988 ( .A(n1226), .B(n1288), .C(n1393), .Y(n2294) );
  NAND2X1 U989 ( .A(\mem<27><4> ), .B(n18), .Y(n1394) );
  OAI21X1 U990 ( .A(n1226), .B(n1289), .C(n1394), .Y(n2293) );
  NAND2X1 U991 ( .A(\mem<27><5> ), .B(n18), .Y(n1395) );
  OAI21X1 U992 ( .A(n1226), .B(n1292), .C(n1395), .Y(n2292) );
  NAND2X1 U993 ( .A(\mem<27><6> ), .B(n18), .Y(n1396) );
  OAI21X1 U994 ( .A(n1226), .B(n1293), .C(n1396), .Y(n2291) );
  NAND2X1 U995 ( .A(\mem<27><7> ), .B(n18), .Y(n1397) );
  OAI21X1 U996 ( .A(n1226), .B(n1296), .C(n1397), .Y(n2290) );
  NAND2X1 U997 ( .A(\mem<27><8> ), .B(n18), .Y(n1398) );
  OAI21X1 U998 ( .A(n1227), .B(n1297), .C(n1398), .Y(n2289) );
  NAND2X1 U999 ( .A(\mem<27><9> ), .B(n18), .Y(n1399) );
  OAI21X1 U1000 ( .A(n1227), .B(n1300), .C(n1399), .Y(n2288) );
  NAND2X1 U1001 ( .A(\mem<27><10> ), .B(n18), .Y(n1400) );
  OAI21X1 U1002 ( .A(n1227), .B(n1301), .C(n1400), .Y(n2287) );
  NAND2X1 U1003 ( .A(\mem<27><11> ), .B(n18), .Y(n1401) );
  OAI21X1 U1004 ( .A(n1227), .B(n1304), .C(n1401), .Y(n2286) );
  NAND2X1 U1005 ( .A(\mem<27><12> ), .B(n18), .Y(n1402) );
  OAI21X1 U1006 ( .A(n1227), .B(n1305), .C(n1402), .Y(n2285) );
  NAND2X1 U1007 ( .A(\mem<27><13> ), .B(n18), .Y(n1403) );
  OAI21X1 U1008 ( .A(n1227), .B(n1307), .C(n1403), .Y(n2284) );
  NAND2X1 U1009 ( .A(\mem<27><14> ), .B(n18), .Y(n1404) );
  OAI21X1 U1010 ( .A(n1227), .B(n1309), .C(n1404), .Y(n2283) );
  NAND2X1 U1011 ( .A(\mem<27><15> ), .B(n18), .Y(n1405) );
  OAI21X1 U1012 ( .A(n1227), .B(n1311), .C(n1405), .Y(n2282) );
  NAND3X1 U1013 ( .A(n1318), .B(n1315), .C(n1314), .Y(n1406) );
  NAND2X1 U1014 ( .A(\mem<26><0> ), .B(n20), .Y(n1407) );
  OAI21X1 U1015 ( .A(n1228), .B(n1281), .C(n1407), .Y(n2281) );
  NAND2X1 U1016 ( .A(\mem<26><1> ), .B(n20), .Y(n1408) );
  OAI21X1 U1017 ( .A(n1228), .B(n1283), .C(n1408), .Y(n2280) );
  NAND2X1 U1018 ( .A(\mem<26><2> ), .B(n20), .Y(n1409) );
  OAI21X1 U1019 ( .A(n1228), .B(n1286), .C(n1409), .Y(n2279) );
  NAND2X1 U1020 ( .A(\mem<26><3> ), .B(n20), .Y(n1410) );
  OAI21X1 U1021 ( .A(n1228), .B(n1287), .C(n1410), .Y(n2278) );
  NAND2X1 U1022 ( .A(\mem<26><4> ), .B(n20), .Y(n1411) );
  OAI21X1 U1023 ( .A(n1228), .B(n1290), .C(n1411), .Y(n2277) );
  NAND2X1 U1024 ( .A(\mem<26><5> ), .B(n20), .Y(n1412) );
  OAI21X1 U1025 ( .A(n1228), .B(n1291), .C(n1412), .Y(n2276) );
  NAND2X1 U1026 ( .A(\mem<26><6> ), .B(n20), .Y(n1413) );
  OAI21X1 U1027 ( .A(n1228), .B(n1294), .C(n1413), .Y(n2275) );
  NAND2X1 U1028 ( .A(\mem<26><7> ), .B(n20), .Y(n1414) );
  OAI21X1 U1029 ( .A(n1228), .B(n1295), .C(n1414), .Y(n2274) );
  NAND2X1 U1030 ( .A(\mem<26><8> ), .B(n20), .Y(n1415) );
  OAI21X1 U1031 ( .A(n1229), .B(n1298), .C(n1415), .Y(n2273) );
  NAND2X1 U1032 ( .A(\mem<26><9> ), .B(n20), .Y(n1416) );
  OAI21X1 U1033 ( .A(n1229), .B(n1299), .C(n1416), .Y(n2272) );
  NAND2X1 U1034 ( .A(\mem<26><10> ), .B(n20), .Y(n1417) );
  OAI21X1 U1035 ( .A(n1229), .B(n1302), .C(n1417), .Y(n2271) );
  NAND2X1 U1036 ( .A(\mem<26><11> ), .B(n20), .Y(n1418) );
  OAI21X1 U1037 ( .A(n1229), .B(n1303), .C(n1418), .Y(n2270) );
  NAND2X1 U1038 ( .A(\mem<26><12> ), .B(n20), .Y(n1419) );
  OAI21X1 U1039 ( .A(n1229), .B(n1305), .C(n1419), .Y(n2269) );
  NAND2X1 U1040 ( .A(\mem<26><13> ), .B(n20), .Y(n1420) );
  OAI21X1 U1041 ( .A(n1229), .B(n1306), .C(n1420), .Y(n2268) );
  NAND2X1 U1042 ( .A(\mem<26><14> ), .B(n20), .Y(n1421) );
  OAI21X1 U1043 ( .A(n1229), .B(n1308), .C(n1421), .Y(n2267) );
  NAND2X1 U1044 ( .A(\mem<26><15> ), .B(n20), .Y(n1422) );
  OAI21X1 U1045 ( .A(n1229), .B(n1310), .C(n1422), .Y(n2266) );
  NAND3X1 U1046 ( .A(n1313), .B(n1318), .C(n1316), .Y(n1423) );
  NAND2X1 U1047 ( .A(\mem<25><0> ), .B(n22), .Y(n1424) );
  OAI21X1 U1048 ( .A(n1230), .B(n1281), .C(n1424), .Y(n2265) );
  NAND2X1 U1049 ( .A(\mem<25><1> ), .B(n22), .Y(n1425) );
  OAI21X1 U1050 ( .A(n1230), .B(n1284), .C(n1425), .Y(n2264) );
  NAND2X1 U1051 ( .A(\mem<25><2> ), .B(n22), .Y(n1426) );
  OAI21X1 U1052 ( .A(n1230), .B(n1285), .C(n1426), .Y(n2263) );
  NAND2X1 U1053 ( .A(\mem<25><3> ), .B(n22), .Y(n1427) );
  OAI21X1 U1054 ( .A(n1230), .B(n1288), .C(n1427), .Y(n2262) );
  NAND2X1 U1055 ( .A(\mem<25><4> ), .B(n22), .Y(n1428) );
  OAI21X1 U1056 ( .A(n1230), .B(n1289), .C(n1428), .Y(n2261) );
  NAND2X1 U1057 ( .A(\mem<25><5> ), .B(n22), .Y(n1429) );
  OAI21X1 U1058 ( .A(n1230), .B(n1292), .C(n1429), .Y(n2260) );
  NAND2X1 U1059 ( .A(\mem<25><6> ), .B(n22), .Y(n1430) );
  OAI21X1 U1060 ( .A(n1230), .B(n1293), .C(n1430), .Y(n2259) );
  NAND2X1 U1061 ( .A(\mem<25><7> ), .B(n22), .Y(n1431) );
  OAI21X1 U1062 ( .A(n1230), .B(n1296), .C(n1431), .Y(n2258) );
  NAND2X1 U1063 ( .A(\mem<25><8> ), .B(n22), .Y(n1432) );
  OAI21X1 U1064 ( .A(n1231), .B(n1297), .C(n1432), .Y(n2257) );
  NAND2X1 U1065 ( .A(\mem<25><9> ), .B(n22), .Y(n1433) );
  OAI21X1 U1066 ( .A(n1231), .B(n1300), .C(n1433), .Y(n2256) );
  NAND2X1 U1067 ( .A(\mem<25><10> ), .B(n22), .Y(n1434) );
  OAI21X1 U1068 ( .A(n1231), .B(n1301), .C(n1434), .Y(n2255) );
  NAND2X1 U1069 ( .A(\mem<25><11> ), .B(n22), .Y(n1435) );
  OAI21X1 U1070 ( .A(n1231), .B(n1304), .C(n1435), .Y(n2254) );
  NAND2X1 U1071 ( .A(\mem<25><12> ), .B(n22), .Y(n1436) );
  OAI21X1 U1072 ( .A(n1231), .B(n1305), .C(n1436), .Y(n2253) );
  NAND2X1 U1073 ( .A(\mem<25><13> ), .B(n22), .Y(n1437) );
  OAI21X1 U1074 ( .A(n1231), .B(n1307), .C(n1437), .Y(n2252) );
  NAND2X1 U1075 ( .A(\mem<25><14> ), .B(n22), .Y(n1438) );
  OAI21X1 U1076 ( .A(n1231), .B(n1309), .C(n1438), .Y(n2251) );
  NAND2X1 U1077 ( .A(\mem<25><15> ), .B(n22), .Y(n1439) );
  OAI21X1 U1078 ( .A(n1231), .B(n1311), .C(n1439), .Y(n2250) );
  NOR3X1 U1079 ( .A(n1313), .B(n1315), .C(n1317), .Y(n1833) );
  NAND2X1 U1080 ( .A(\mem<24><0> ), .B(n24), .Y(n1440) );
  OAI21X1 U1081 ( .A(n1232), .B(n1281), .C(n1440), .Y(n2249) );
  NAND2X1 U1082 ( .A(\mem<24><1> ), .B(n24), .Y(n1441) );
  OAI21X1 U1083 ( .A(n1232), .B(n1283), .C(n1441), .Y(n2248) );
  NAND2X1 U1084 ( .A(\mem<24><2> ), .B(n24), .Y(n1442) );
  OAI21X1 U1085 ( .A(n1232), .B(n1285), .C(n1442), .Y(n2247) );
  NAND2X1 U1086 ( .A(\mem<24><3> ), .B(n24), .Y(n1443) );
  OAI21X1 U1087 ( .A(n1232), .B(n1287), .C(n1443), .Y(n2246) );
  NAND2X1 U1088 ( .A(\mem<24><4> ), .B(n24), .Y(n1444) );
  OAI21X1 U1089 ( .A(n1232), .B(n1289), .C(n1444), .Y(n2245) );
  NAND2X1 U1090 ( .A(\mem<24><5> ), .B(n24), .Y(n1445) );
  OAI21X1 U1091 ( .A(n1232), .B(n1291), .C(n1445), .Y(n2244) );
  NAND2X1 U1092 ( .A(\mem<24><6> ), .B(n24), .Y(n1446) );
  OAI21X1 U1093 ( .A(n1232), .B(n1293), .C(n1446), .Y(n2243) );
  NAND2X1 U1094 ( .A(\mem<24><7> ), .B(n24), .Y(n1447) );
  OAI21X1 U1095 ( .A(n1232), .B(n1295), .C(n1447), .Y(n2242) );
  NAND2X1 U1096 ( .A(\mem<24><8> ), .B(n24), .Y(n1448) );
  OAI21X1 U1097 ( .A(n1232), .B(n1297), .C(n1448), .Y(n2241) );
  NAND2X1 U1098 ( .A(\mem<24><9> ), .B(n24), .Y(n1449) );
  OAI21X1 U1099 ( .A(n1232), .B(n1299), .C(n1449), .Y(n2240) );
  NAND2X1 U1100 ( .A(\mem<24><10> ), .B(n24), .Y(n1450) );
  OAI21X1 U1101 ( .A(n1232), .B(n1301), .C(n1450), .Y(n2239) );
  NAND2X1 U1102 ( .A(\mem<24><11> ), .B(n24), .Y(n1451) );
  OAI21X1 U1103 ( .A(n1232), .B(n1303), .C(n1451), .Y(n2238) );
  NAND2X1 U1104 ( .A(\mem<24><12> ), .B(n24), .Y(n1452) );
  OAI21X1 U1105 ( .A(n1232), .B(n1305), .C(n1452), .Y(n2237) );
  NAND2X1 U1106 ( .A(\mem<24><13> ), .B(n24), .Y(n1453) );
  OAI21X1 U1107 ( .A(n1232), .B(n1306), .C(n1453), .Y(n2236) );
  NAND2X1 U1108 ( .A(\mem<24><14> ), .B(n24), .Y(n1454) );
  OAI21X1 U1109 ( .A(n1232), .B(n1308), .C(n1454), .Y(n2235) );
  NAND2X1 U1110 ( .A(\mem<24><15> ), .B(n24), .Y(n1455) );
  OAI21X1 U1111 ( .A(n1232), .B(n1310), .C(n1455), .Y(n2234) );
  NAND2X1 U1112 ( .A(\mem<23><0> ), .B(n26), .Y(n1456) );
  OAI21X1 U1113 ( .A(n1233), .B(n1281), .C(n1456), .Y(n2233) );
  NAND2X1 U1114 ( .A(\mem<23><1> ), .B(n26), .Y(n1457) );
  OAI21X1 U1115 ( .A(n1233), .B(n1284), .C(n1457), .Y(n2232) );
  NAND2X1 U1116 ( .A(\mem<23><2> ), .B(n26), .Y(n1458) );
  OAI21X1 U1117 ( .A(n1233), .B(n1286), .C(n1458), .Y(n2231) );
  NAND2X1 U1118 ( .A(\mem<23><3> ), .B(n26), .Y(n1459) );
  OAI21X1 U1119 ( .A(n1233), .B(n1288), .C(n1459), .Y(n2230) );
  NAND2X1 U1120 ( .A(\mem<23><4> ), .B(n26), .Y(n1460) );
  OAI21X1 U1121 ( .A(n1233), .B(n1290), .C(n1460), .Y(n2229) );
  NAND2X1 U1122 ( .A(\mem<23><5> ), .B(n26), .Y(n1461) );
  OAI21X1 U1123 ( .A(n1233), .B(n1292), .C(n1461), .Y(n2228) );
  NAND2X1 U1124 ( .A(\mem<23><6> ), .B(n26), .Y(n1462) );
  OAI21X1 U1125 ( .A(n1233), .B(n1294), .C(n1462), .Y(n2227) );
  NAND2X1 U1126 ( .A(\mem<23><7> ), .B(n26), .Y(n1463) );
  OAI21X1 U1127 ( .A(n1233), .B(n1296), .C(n1463), .Y(n2226) );
  NAND2X1 U1128 ( .A(\mem<23><8> ), .B(n26), .Y(n1464) );
  OAI21X1 U1129 ( .A(n1234), .B(n1298), .C(n1464), .Y(n2225) );
  NAND2X1 U1130 ( .A(\mem<23><9> ), .B(n26), .Y(n1465) );
  OAI21X1 U1131 ( .A(n1234), .B(n1300), .C(n1465), .Y(n2224) );
  NAND2X1 U1132 ( .A(\mem<23><10> ), .B(n26), .Y(n1466) );
  OAI21X1 U1133 ( .A(n1234), .B(n1302), .C(n1466), .Y(n2223) );
  NAND2X1 U1134 ( .A(\mem<23><11> ), .B(n26), .Y(n1467) );
  OAI21X1 U1135 ( .A(n1234), .B(n1304), .C(n1467), .Y(n2222) );
  NAND2X1 U1136 ( .A(\mem<23><12> ), .B(n26), .Y(n1468) );
  OAI21X1 U1137 ( .A(n1234), .B(n1305), .C(n1468), .Y(n2221) );
  NAND2X1 U1138 ( .A(\mem<23><13> ), .B(n26), .Y(n1469) );
  OAI21X1 U1139 ( .A(n1234), .B(n1307), .C(n1469), .Y(n2220) );
  NAND2X1 U1140 ( .A(\mem<23><14> ), .B(n26), .Y(n1470) );
  OAI21X1 U1141 ( .A(n1234), .B(n1309), .C(n1470), .Y(n2219) );
  NAND2X1 U1142 ( .A(\mem<23><15> ), .B(n26), .Y(n1471) );
  OAI21X1 U1143 ( .A(n1234), .B(n1311), .C(n1471), .Y(n2218) );
  NAND2X1 U1144 ( .A(\mem<22><0> ), .B(n28), .Y(n1472) );
  OAI21X1 U1145 ( .A(n1235), .B(n1281), .C(n1472), .Y(n2217) );
  NAND2X1 U1146 ( .A(\mem<22><1> ), .B(n28), .Y(n1473) );
  OAI21X1 U1147 ( .A(n1235), .B(n1284), .C(n1473), .Y(n2216) );
  NAND2X1 U1148 ( .A(\mem<22><2> ), .B(n28), .Y(n1474) );
  OAI21X1 U1149 ( .A(n1235), .B(n1286), .C(n1474), .Y(n2215) );
  NAND2X1 U1150 ( .A(\mem<22><3> ), .B(n28), .Y(n1475) );
  OAI21X1 U1151 ( .A(n1235), .B(n1288), .C(n1475), .Y(n2214) );
  NAND2X1 U1152 ( .A(\mem<22><4> ), .B(n28), .Y(n1476) );
  OAI21X1 U1153 ( .A(n1235), .B(n1290), .C(n1476), .Y(n2213) );
  NAND2X1 U1154 ( .A(\mem<22><5> ), .B(n28), .Y(n1477) );
  OAI21X1 U1155 ( .A(n1235), .B(n1292), .C(n1477), .Y(n2212) );
  NAND2X1 U1156 ( .A(\mem<22><6> ), .B(n28), .Y(n1478) );
  OAI21X1 U1157 ( .A(n1235), .B(n1294), .C(n1478), .Y(n2211) );
  NAND2X1 U1158 ( .A(\mem<22><7> ), .B(n28), .Y(n1479) );
  OAI21X1 U1159 ( .A(n1235), .B(n1296), .C(n1479), .Y(n2210) );
  NAND2X1 U1160 ( .A(\mem<22><8> ), .B(n28), .Y(n1480) );
  OAI21X1 U1161 ( .A(n1236), .B(n1298), .C(n1480), .Y(n2209) );
  NAND2X1 U1162 ( .A(\mem<22><9> ), .B(n28), .Y(n1481) );
  OAI21X1 U1163 ( .A(n1236), .B(n1300), .C(n1481), .Y(n2208) );
  NAND2X1 U1164 ( .A(\mem<22><10> ), .B(n28), .Y(n1482) );
  OAI21X1 U1165 ( .A(n1236), .B(n1302), .C(n1482), .Y(n2207) );
  NAND2X1 U1166 ( .A(\mem<22><11> ), .B(n28), .Y(n1483) );
  OAI21X1 U1167 ( .A(n1236), .B(n1304), .C(n1483), .Y(n2206) );
  NAND2X1 U1168 ( .A(\mem<22><12> ), .B(n28), .Y(n1484) );
  OAI21X1 U1169 ( .A(n1236), .B(n1305), .C(n1484), .Y(n2205) );
  NAND2X1 U1170 ( .A(\mem<22><13> ), .B(n28), .Y(n1485) );
  OAI21X1 U1171 ( .A(n1236), .B(n1307), .C(n1485), .Y(n2204) );
  NAND2X1 U1172 ( .A(\mem<22><14> ), .B(n28), .Y(n1486) );
  OAI21X1 U1173 ( .A(n1236), .B(n1309), .C(n1486), .Y(n2203) );
  NAND2X1 U1174 ( .A(\mem<22><15> ), .B(n28), .Y(n1487) );
  OAI21X1 U1175 ( .A(n1236), .B(n1311), .C(n1487), .Y(n2202) );
  NAND2X1 U1177 ( .A(\mem<21><0> ), .B(n30), .Y(n1488) );
  OAI21X1 U1178 ( .A(n1237), .B(n1281), .C(n1488), .Y(n2201) );
  NAND2X1 U1179 ( .A(\mem<21><1> ), .B(n30), .Y(n1489) );
  OAI21X1 U1180 ( .A(n1237), .B(n1284), .C(n1489), .Y(n2200) );
  NAND2X1 U1181 ( .A(\mem<21><2> ), .B(n30), .Y(n1490) );
  OAI21X1 U1182 ( .A(n1237), .B(n1286), .C(n1490), .Y(n2199) );
  NAND2X1 U1183 ( .A(\mem<21><3> ), .B(n30), .Y(n1491) );
  OAI21X1 U1184 ( .A(n1237), .B(n1288), .C(n1491), .Y(n2198) );
  NAND2X1 U1185 ( .A(\mem<21><4> ), .B(n30), .Y(n1492) );
  OAI21X1 U1186 ( .A(n1237), .B(n1290), .C(n1492), .Y(n2197) );
  NAND2X1 U1187 ( .A(\mem<21><5> ), .B(n30), .Y(n1493) );
  OAI21X1 U1188 ( .A(n1237), .B(n1292), .C(n1493), .Y(n2196) );
  NAND2X1 U1189 ( .A(\mem<21><6> ), .B(n30), .Y(n1494) );
  OAI21X1 U1190 ( .A(n1237), .B(n1294), .C(n1494), .Y(n2195) );
  NAND2X1 U1191 ( .A(\mem<21><7> ), .B(n30), .Y(n1495) );
  OAI21X1 U1192 ( .A(n1237), .B(n1296), .C(n1495), .Y(n2194) );
  NAND2X1 U1193 ( .A(\mem<21><8> ), .B(n30), .Y(n1496) );
  OAI21X1 U1194 ( .A(n1238), .B(n1298), .C(n1496), .Y(n2193) );
  NAND2X1 U1195 ( .A(\mem<21><9> ), .B(n30), .Y(n1497) );
  OAI21X1 U1196 ( .A(n1238), .B(n1300), .C(n1497), .Y(n2192) );
  NAND2X1 U1197 ( .A(\mem<21><10> ), .B(n30), .Y(n1498) );
  OAI21X1 U1198 ( .A(n1238), .B(n1302), .C(n1498), .Y(n2191) );
  NAND2X1 U1199 ( .A(\mem<21><11> ), .B(n30), .Y(n1499) );
  OAI21X1 U1200 ( .A(n1238), .B(n1304), .C(n1499), .Y(n2190) );
  NAND2X1 U1201 ( .A(\mem<21><12> ), .B(n30), .Y(n1500) );
  OAI21X1 U1202 ( .A(n1238), .B(n1305), .C(n1500), .Y(n2189) );
  NAND2X1 U1203 ( .A(\mem<21><13> ), .B(n30), .Y(n1501) );
  OAI21X1 U1204 ( .A(n1238), .B(n1307), .C(n1501), .Y(n2188) );
  NAND2X1 U1205 ( .A(\mem<21><14> ), .B(n30), .Y(n1502) );
  OAI21X1 U1206 ( .A(n1238), .B(n1309), .C(n1502), .Y(n2187) );
  NAND2X1 U1207 ( .A(\mem<21><15> ), .B(n30), .Y(n1503) );
  OAI21X1 U1208 ( .A(n1238), .B(n1311), .C(n1503), .Y(n2186) );
  NAND2X1 U1209 ( .A(\mem<20><0> ), .B(n32), .Y(n1504) );
  OAI21X1 U1210 ( .A(n1239), .B(n1281), .C(n1504), .Y(n2185) );
  NAND2X1 U1211 ( .A(\mem<20><1> ), .B(n32), .Y(n1505) );
  OAI21X1 U1212 ( .A(n1239), .B(n1284), .C(n1505), .Y(n2184) );
  NAND2X1 U1213 ( .A(\mem<20><2> ), .B(n32), .Y(n1506) );
  OAI21X1 U1214 ( .A(n1239), .B(n1286), .C(n1506), .Y(n2183) );
  NAND2X1 U1215 ( .A(\mem<20><3> ), .B(n32), .Y(n1507) );
  OAI21X1 U1216 ( .A(n1239), .B(n1288), .C(n1507), .Y(n2182) );
  NAND2X1 U1217 ( .A(\mem<20><4> ), .B(n32), .Y(n1508) );
  OAI21X1 U1218 ( .A(n1239), .B(n1290), .C(n1508), .Y(n2181) );
  NAND2X1 U1219 ( .A(\mem<20><5> ), .B(n32), .Y(n1509) );
  OAI21X1 U1220 ( .A(n1239), .B(n1292), .C(n1509), .Y(n2180) );
  NAND2X1 U1221 ( .A(\mem<20><6> ), .B(n32), .Y(n1510) );
  OAI21X1 U1222 ( .A(n1239), .B(n1294), .C(n1510), .Y(n2179) );
  NAND2X1 U1223 ( .A(\mem<20><7> ), .B(n32), .Y(n1511) );
  OAI21X1 U1224 ( .A(n1239), .B(n1296), .C(n1511), .Y(n2178) );
  NAND2X1 U1225 ( .A(\mem<20><8> ), .B(n32), .Y(n1512) );
  OAI21X1 U1226 ( .A(n1240), .B(n1298), .C(n1512), .Y(n2177) );
  NAND2X1 U1227 ( .A(\mem<20><9> ), .B(n32), .Y(n1513) );
  OAI21X1 U1228 ( .A(n1240), .B(n1300), .C(n1513), .Y(n2176) );
  NAND2X1 U1229 ( .A(\mem<20><10> ), .B(n32), .Y(n1514) );
  OAI21X1 U1230 ( .A(n1240), .B(n1302), .C(n1514), .Y(n2175) );
  NAND2X1 U1231 ( .A(\mem<20><11> ), .B(n32), .Y(n1515) );
  OAI21X1 U1232 ( .A(n1240), .B(n1304), .C(n1515), .Y(n2174) );
  NAND2X1 U1233 ( .A(\mem<20><12> ), .B(n32), .Y(n1516) );
  OAI21X1 U1234 ( .A(n1240), .B(n1305), .C(n1516), .Y(n2173) );
  NAND2X1 U1235 ( .A(\mem<20><13> ), .B(n32), .Y(n1517) );
  OAI21X1 U1236 ( .A(n1240), .B(n1307), .C(n1517), .Y(n2172) );
  NAND2X1 U1237 ( .A(\mem<20><14> ), .B(n32), .Y(n1518) );
  OAI21X1 U1238 ( .A(n1240), .B(n1309), .C(n1518), .Y(n2171) );
  NAND2X1 U1239 ( .A(\mem<20><15> ), .B(n32), .Y(n1519) );
  OAI21X1 U1240 ( .A(n1240), .B(n1311), .C(n1519), .Y(n2170) );
  NAND2X1 U1241 ( .A(\mem<19><0> ), .B(n34), .Y(n1520) );
  OAI21X1 U1242 ( .A(n1241), .B(n1282), .C(n1520), .Y(n2169) );
  NAND2X1 U1243 ( .A(\mem<19><1> ), .B(n34), .Y(n1521) );
  OAI21X1 U1244 ( .A(n1241), .B(n1284), .C(n1521), .Y(n2168) );
  NAND2X1 U1245 ( .A(\mem<19><2> ), .B(n34), .Y(n1522) );
  OAI21X1 U1246 ( .A(n1241), .B(n1286), .C(n1522), .Y(n2167) );
  NAND2X1 U1247 ( .A(\mem<19><3> ), .B(n34), .Y(n1523) );
  OAI21X1 U1248 ( .A(n1241), .B(n1288), .C(n1523), .Y(n2166) );
  NAND2X1 U1249 ( .A(\mem<19><4> ), .B(n34), .Y(n1524) );
  OAI21X1 U1250 ( .A(n1241), .B(n1290), .C(n1524), .Y(n2165) );
  NAND2X1 U1251 ( .A(\mem<19><5> ), .B(n34), .Y(n1525) );
  OAI21X1 U1252 ( .A(n1241), .B(n1292), .C(n1525), .Y(n2164) );
  NAND2X1 U1253 ( .A(\mem<19><6> ), .B(n34), .Y(n1526) );
  OAI21X1 U1254 ( .A(n1241), .B(n1294), .C(n1526), .Y(n2163) );
  NAND2X1 U1255 ( .A(\mem<19><7> ), .B(n34), .Y(n1527) );
  OAI21X1 U1256 ( .A(n1241), .B(n1296), .C(n1527), .Y(n2162) );
  NAND2X1 U1257 ( .A(\mem<19><8> ), .B(n34), .Y(n1528) );
  OAI21X1 U1258 ( .A(n1242), .B(n1298), .C(n1528), .Y(n2161) );
  NAND2X1 U1259 ( .A(\mem<19><9> ), .B(n34), .Y(n1529) );
  OAI21X1 U1260 ( .A(n1242), .B(n1300), .C(n1529), .Y(n2160) );
  NAND2X1 U1261 ( .A(\mem<19><10> ), .B(n34), .Y(n1530) );
  OAI21X1 U1262 ( .A(n1242), .B(n1302), .C(n1530), .Y(n2159) );
  NAND2X1 U1263 ( .A(\mem<19><11> ), .B(n34), .Y(n1531) );
  OAI21X1 U1264 ( .A(n1242), .B(n1304), .C(n1531), .Y(n2158) );
  NAND2X1 U1265 ( .A(\mem<19><12> ), .B(n34), .Y(n1532) );
  OAI21X1 U1266 ( .A(n1242), .B(n1305), .C(n1532), .Y(n2157) );
  NAND2X1 U1267 ( .A(\mem<19><13> ), .B(n34), .Y(n1533) );
  OAI21X1 U1268 ( .A(n1242), .B(n1307), .C(n1533), .Y(n2156) );
  NAND2X1 U1269 ( .A(\mem<19><14> ), .B(n34), .Y(n1534) );
  OAI21X1 U1270 ( .A(n1242), .B(n1309), .C(n1534), .Y(n2155) );
  NAND2X1 U1271 ( .A(\mem<19><15> ), .B(n34), .Y(n1535) );
  OAI21X1 U1272 ( .A(n1242), .B(n1311), .C(n1535), .Y(n2154) );
  NAND2X1 U1273 ( .A(\mem<18><0> ), .B(n36), .Y(n1536) );
  OAI21X1 U1274 ( .A(n1243), .B(n1282), .C(n1536), .Y(n2153) );
  NAND2X1 U1275 ( .A(\mem<18><1> ), .B(n36), .Y(n1537) );
  OAI21X1 U1276 ( .A(n1243), .B(n1284), .C(n1537), .Y(n2152) );
  NAND2X1 U1277 ( .A(\mem<18><2> ), .B(n36), .Y(n1538) );
  OAI21X1 U1278 ( .A(n1243), .B(n1286), .C(n1538), .Y(n2151) );
  NAND2X1 U1279 ( .A(\mem<18><3> ), .B(n36), .Y(n1539) );
  OAI21X1 U1280 ( .A(n1243), .B(n1288), .C(n1539), .Y(n2150) );
  NAND2X1 U1281 ( .A(\mem<18><4> ), .B(n36), .Y(n1540) );
  OAI21X1 U1282 ( .A(n1243), .B(n1290), .C(n1540), .Y(n2149) );
  NAND2X1 U1283 ( .A(\mem<18><5> ), .B(n36), .Y(n1541) );
  OAI21X1 U1284 ( .A(n1243), .B(n1292), .C(n1541), .Y(n2148) );
  NAND2X1 U1285 ( .A(\mem<18><6> ), .B(n36), .Y(n1542) );
  OAI21X1 U1286 ( .A(n1243), .B(n1294), .C(n1542), .Y(n2147) );
  NAND2X1 U1287 ( .A(\mem<18><7> ), .B(n36), .Y(n1543) );
  OAI21X1 U1288 ( .A(n1243), .B(n1296), .C(n1543), .Y(n2146) );
  NAND2X1 U1289 ( .A(\mem<18><8> ), .B(n36), .Y(n1544) );
  OAI21X1 U1290 ( .A(n1244), .B(n1298), .C(n1544), .Y(n2145) );
  NAND2X1 U1291 ( .A(\mem<18><9> ), .B(n36), .Y(n1545) );
  OAI21X1 U1292 ( .A(n1244), .B(n1300), .C(n1545), .Y(n2144) );
  NAND2X1 U1293 ( .A(\mem<18><10> ), .B(n36), .Y(n1546) );
  OAI21X1 U1294 ( .A(n1244), .B(n1302), .C(n1546), .Y(n2143) );
  NAND2X1 U1295 ( .A(\mem<18><11> ), .B(n36), .Y(n1547) );
  OAI21X1 U1296 ( .A(n1244), .B(n1304), .C(n1547), .Y(n2142) );
  NAND2X1 U1297 ( .A(\mem<18><12> ), .B(n36), .Y(n1548) );
  OAI21X1 U1298 ( .A(n1244), .B(n1305), .C(n1548), .Y(n2141) );
  NAND2X1 U1299 ( .A(\mem<18><13> ), .B(n36), .Y(n1549) );
  OAI21X1 U1300 ( .A(n1244), .B(n1307), .C(n1549), .Y(n2140) );
  NAND2X1 U1301 ( .A(\mem<18><14> ), .B(n36), .Y(n1550) );
  OAI21X1 U1302 ( .A(n1244), .B(n1309), .C(n1550), .Y(n2139) );
  NAND2X1 U1303 ( .A(\mem<18><15> ), .B(n36), .Y(n1551) );
  OAI21X1 U1304 ( .A(n1244), .B(n1311), .C(n1551), .Y(n2138) );
  NAND2X1 U1305 ( .A(\mem<17><0> ), .B(n38), .Y(n1552) );
  OAI21X1 U1306 ( .A(n1245), .B(n1282), .C(n1552), .Y(n2137) );
  NAND2X1 U1307 ( .A(\mem<17><1> ), .B(n38), .Y(n1553) );
  OAI21X1 U1308 ( .A(n1245), .B(n1284), .C(n1553), .Y(n2136) );
  NAND2X1 U1309 ( .A(\mem<17><2> ), .B(n38), .Y(n1554) );
  OAI21X1 U1310 ( .A(n1245), .B(n1286), .C(n1554), .Y(n2135) );
  NAND2X1 U1311 ( .A(\mem<17><3> ), .B(n38), .Y(n1555) );
  OAI21X1 U1312 ( .A(n1245), .B(n1288), .C(n1555), .Y(n2134) );
  NAND2X1 U1313 ( .A(\mem<17><4> ), .B(n38), .Y(n1556) );
  OAI21X1 U1314 ( .A(n1245), .B(n1290), .C(n1556), .Y(n2133) );
  NAND2X1 U1315 ( .A(\mem<17><5> ), .B(n38), .Y(n1557) );
  OAI21X1 U1316 ( .A(n1245), .B(n1292), .C(n1557), .Y(n2132) );
  NAND2X1 U1317 ( .A(\mem<17><6> ), .B(n38), .Y(n1558) );
  OAI21X1 U1318 ( .A(n1245), .B(n1294), .C(n1558), .Y(n2131) );
  NAND2X1 U1319 ( .A(\mem<17><7> ), .B(n38), .Y(n1559) );
  OAI21X1 U1320 ( .A(n1245), .B(n1296), .C(n1559), .Y(n2130) );
  NAND2X1 U1321 ( .A(\mem<17><8> ), .B(n38), .Y(n1560) );
  OAI21X1 U1322 ( .A(n1246), .B(n1298), .C(n1560), .Y(n2129) );
  NAND2X1 U1323 ( .A(\mem<17><9> ), .B(n38), .Y(n1561) );
  OAI21X1 U1324 ( .A(n1246), .B(n1300), .C(n1561), .Y(n2128) );
  NAND2X1 U1325 ( .A(\mem<17><10> ), .B(n38), .Y(n1562) );
  OAI21X1 U1326 ( .A(n1246), .B(n1302), .C(n1562), .Y(n2127) );
  NAND2X1 U1327 ( .A(\mem<17><11> ), .B(n38), .Y(n1563) );
  OAI21X1 U1328 ( .A(n1246), .B(n1304), .C(n1563), .Y(n2126) );
  NAND2X1 U1329 ( .A(\mem<17><12> ), .B(n38), .Y(n1564) );
  OAI21X1 U1330 ( .A(n1246), .B(n1305), .C(n1564), .Y(n2125) );
  NAND2X1 U1331 ( .A(\mem<17><13> ), .B(n38), .Y(n1565) );
  OAI21X1 U1332 ( .A(n1246), .B(n1307), .C(n1565), .Y(n2124) );
  NAND2X1 U1333 ( .A(\mem<17><14> ), .B(n38), .Y(n1566) );
  OAI21X1 U1334 ( .A(n1246), .B(n1309), .C(n1566), .Y(n2123) );
  NAND2X1 U1335 ( .A(\mem<17><15> ), .B(n38), .Y(n1567) );
  OAI21X1 U1336 ( .A(n1246), .B(n1311), .C(n1567), .Y(n2122) );
  NAND2X1 U1337 ( .A(\mem<16><0> ), .B(n40), .Y(n1568) );
  OAI21X1 U1338 ( .A(n1247), .B(n1282), .C(n1568), .Y(n2121) );
  NAND2X1 U1339 ( .A(\mem<16><1> ), .B(n40), .Y(n1569) );
  OAI21X1 U1340 ( .A(n1247), .B(n1284), .C(n1569), .Y(n2120) );
  NAND2X1 U1341 ( .A(\mem<16><2> ), .B(n40), .Y(n1570) );
  OAI21X1 U1342 ( .A(n1247), .B(n1286), .C(n1570), .Y(n2119) );
  NAND2X1 U1343 ( .A(\mem<16><3> ), .B(n40), .Y(n1571) );
  OAI21X1 U1344 ( .A(n1247), .B(n1288), .C(n1571), .Y(n2118) );
  NAND2X1 U1345 ( .A(\mem<16><4> ), .B(n40), .Y(n1572) );
  OAI21X1 U1346 ( .A(n1247), .B(n1290), .C(n1572), .Y(n2117) );
  NAND2X1 U1347 ( .A(\mem<16><5> ), .B(n40), .Y(n1573) );
  OAI21X1 U1348 ( .A(n1247), .B(n1292), .C(n1573), .Y(n2116) );
  NAND2X1 U1349 ( .A(\mem<16><6> ), .B(n40), .Y(n1574) );
  OAI21X1 U1350 ( .A(n1247), .B(n1294), .C(n1574), .Y(n2115) );
  NAND2X1 U1351 ( .A(\mem<16><7> ), .B(n40), .Y(n1575) );
  OAI21X1 U1352 ( .A(n1247), .B(n1296), .C(n1575), .Y(n2114) );
  NAND2X1 U1353 ( .A(\mem<16><8> ), .B(n40), .Y(n1576) );
  OAI21X1 U1354 ( .A(n1247), .B(n1298), .C(n1576), .Y(n2113) );
  NAND2X1 U1355 ( .A(\mem<16><9> ), .B(n40), .Y(n1577) );
  OAI21X1 U1356 ( .A(n1247), .B(n1300), .C(n1577), .Y(n2112) );
  NAND2X1 U1357 ( .A(\mem<16><10> ), .B(n40), .Y(n1578) );
  OAI21X1 U1358 ( .A(n1247), .B(n1302), .C(n1578), .Y(n2111) );
  NAND2X1 U1359 ( .A(\mem<16><11> ), .B(n40), .Y(n1579) );
  OAI21X1 U1360 ( .A(n1247), .B(n1304), .C(n1579), .Y(n2110) );
  NAND2X1 U1361 ( .A(\mem<16><12> ), .B(n40), .Y(n1580) );
  OAI21X1 U1362 ( .A(n1247), .B(n1305), .C(n1580), .Y(n2109) );
  NAND2X1 U1363 ( .A(\mem<16><13> ), .B(n40), .Y(n1581) );
  OAI21X1 U1364 ( .A(n1247), .B(n1307), .C(n1581), .Y(n2108) );
  NAND2X1 U1365 ( .A(\mem<16><14> ), .B(n40), .Y(n1582) );
  OAI21X1 U1366 ( .A(n1247), .B(n1309), .C(n1582), .Y(n2107) );
  NAND2X1 U1367 ( .A(\mem<16><15> ), .B(n40), .Y(n1583) );
  OAI21X1 U1368 ( .A(n1247), .B(n1311), .C(n1583), .Y(n2106) );
  NAND3X1 U1369 ( .A(n1319), .B(n2362), .C(n1322), .Y(n1584) );
  NAND2X1 U1370 ( .A(\mem<15><0> ), .B(n42), .Y(n1585) );
  OAI21X1 U1371 ( .A(n1248), .B(n1282), .C(n1585), .Y(n2105) );
  NAND2X1 U1372 ( .A(\mem<15><1> ), .B(n42), .Y(n1586) );
  OAI21X1 U1373 ( .A(n1248), .B(n1284), .C(n1586), .Y(n2104) );
  NAND2X1 U1374 ( .A(\mem<15><2> ), .B(n42), .Y(n1587) );
  OAI21X1 U1375 ( .A(n1248), .B(n1286), .C(n1587), .Y(n2103) );
  NAND2X1 U1376 ( .A(\mem<15><3> ), .B(n42), .Y(n1588) );
  OAI21X1 U1377 ( .A(n1248), .B(n1288), .C(n1588), .Y(n2102) );
  NAND2X1 U1378 ( .A(\mem<15><4> ), .B(n42), .Y(n1589) );
  OAI21X1 U1379 ( .A(n1248), .B(n1290), .C(n1589), .Y(n2101) );
  NAND2X1 U1380 ( .A(\mem<15><5> ), .B(n42), .Y(n1590) );
  OAI21X1 U1381 ( .A(n1248), .B(n1292), .C(n1590), .Y(n2100) );
  NAND2X1 U1382 ( .A(\mem<15><6> ), .B(n42), .Y(n1591) );
  OAI21X1 U1383 ( .A(n1248), .B(n1294), .C(n1591), .Y(n2099) );
  NAND2X1 U1384 ( .A(\mem<15><7> ), .B(n42), .Y(n1592) );
  OAI21X1 U1385 ( .A(n1248), .B(n1296), .C(n1592), .Y(n2098) );
  NAND2X1 U1386 ( .A(\mem<15><8> ), .B(n42), .Y(n1593) );
  OAI21X1 U1387 ( .A(n1249), .B(n1298), .C(n1593), .Y(n2097) );
  NAND2X1 U1388 ( .A(\mem<15><9> ), .B(n42), .Y(n1594) );
  OAI21X1 U1389 ( .A(n1249), .B(n1300), .C(n1594), .Y(n2096) );
  NAND2X1 U1390 ( .A(\mem<15><10> ), .B(n42), .Y(n1595) );
  OAI21X1 U1391 ( .A(n1249), .B(n1302), .C(n1595), .Y(n2095) );
  NAND2X1 U1392 ( .A(\mem<15><11> ), .B(n42), .Y(n1596) );
  OAI21X1 U1393 ( .A(n1249), .B(n1304), .C(n1596), .Y(n2094) );
  NAND2X1 U1394 ( .A(\mem<15><12> ), .B(n42), .Y(n1597) );
  OAI21X1 U1395 ( .A(n1249), .B(n1305), .C(n1597), .Y(n2093) );
  NAND2X1 U1396 ( .A(\mem<15><13> ), .B(n42), .Y(n1598) );
  OAI21X1 U1397 ( .A(n1249), .B(n1307), .C(n1598), .Y(n2092) );
  NAND2X1 U1398 ( .A(\mem<15><14> ), .B(n42), .Y(n1599) );
  OAI21X1 U1399 ( .A(n1249), .B(n1309), .C(n1599), .Y(n2091) );
  NAND2X1 U1400 ( .A(\mem<15><15> ), .B(n42), .Y(n1600) );
  OAI21X1 U1401 ( .A(n1249), .B(n1311), .C(n1600), .Y(n2090) );
  NAND2X1 U1402 ( .A(\mem<14><0> ), .B(n44), .Y(n1601) );
  OAI21X1 U1403 ( .A(n1250), .B(n1282), .C(n1601), .Y(n2089) );
  NAND2X1 U1404 ( .A(\mem<14><1> ), .B(n44), .Y(n1602) );
  OAI21X1 U1405 ( .A(n1250), .B(n1284), .C(n1602), .Y(n2088) );
  NAND2X1 U1406 ( .A(\mem<14><2> ), .B(n44), .Y(n1603) );
  OAI21X1 U1407 ( .A(n1250), .B(n1286), .C(n1603), .Y(n2087) );
  NAND2X1 U1408 ( .A(\mem<14><3> ), .B(n44), .Y(n1604) );
  OAI21X1 U1409 ( .A(n1250), .B(n1288), .C(n1604), .Y(n2086) );
  NAND2X1 U1410 ( .A(\mem<14><4> ), .B(n44), .Y(n1605) );
  OAI21X1 U1411 ( .A(n1250), .B(n1290), .C(n1605), .Y(n2085) );
  NAND2X1 U1412 ( .A(\mem<14><5> ), .B(n44), .Y(n1606) );
  OAI21X1 U1413 ( .A(n1250), .B(n1292), .C(n1606), .Y(n2084) );
  NAND2X1 U1414 ( .A(\mem<14><6> ), .B(n44), .Y(n1607) );
  OAI21X1 U1415 ( .A(n1250), .B(n1294), .C(n1607), .Y(n2083) );
  NAND2X1 U1416 ( .A(\mem<14><7> ), .B(n44), .Y(n1608) );
  OAI21X1 U1417 ( .A(n1250), .B(n1296), .C(n1608), .Y(n2082) );
  NAND2X1 U1418 ( .A(\mem<14><8> ), .B(n44), .Y(n1609) );
  OAI21X1 U1419 ( .A(n1251), .B(n1298), .C(n1609), .Y(n2081) );
  NAND2X1 U1420 ( .A(\mem<14><9> ), .B(n44), .Y(n1610) );
  OAI21X1 U1421 ( .A(n1251), .B(n1300), .C(n1610), .Y(n2080) );
  NAND2X1 U1422 ( .A(\mem<14><10> ), .B(n44), .Y(n1611) );
  OAI21X1 U1423 ( .A(n1251), .B(n1302), .C(n1611), .Y(n2079) );
  NAND2X1 U1424 ( .A(\mem<14><11> ), .B(n44), .Y(n1612) );
  OAI21X1 U1425 ( .A(n1251), .B(n1304), .C(n1612), .Y(n2078) );
  NAND2X1 U1426 ( .A(\mem<14><12> ), .B(n44), .Y(n1613) );
  OAI21X1 U1427 ( .A(n1251), .B(n1305), .C(n1613), .Y(n2077) );
  NAND2X1 U1428 ( .A(\mem<14><13> ), .B(n44), .Y(n1614) );
  OAI21X1 U1429 ( .A(n1251), .B(n1307), .C(n1614), .Y(n2076) );
  NAND2X1 U1430 ( .A(\mem<14><14> ), .B(n44), .Y(n1615) );
  OAI21X1 U1431 ( .A(n1251), .B(n1309), .C(n1615), .Y(n2075) );
  NAND2X1 U1432 ( .A(\mem<14><15> ), .B(n44), .Y(n1616) );
  OAI21X1 U1433 ( .A(n1251), .B(n1311), .C(n1616), .Y(n2074) );
  NAND2X1 U1434 ( .A(\mem<13><0> ), .B(n46), .Y(n1617) );
  OAI21X1 U1435 ( .A(n1252), .B(n1282), .C(n1617), .Y(n2073) );
  NAND2X1 U1436 ( .A(\mem<13><1> ), .B(n46), .Y(n1618) );
  OAI21X1 U1437 ( .A(n1252), .B(n1284), .C(n1618), .Y(n2072) );
  NAND2X1 U1438 ( .A(\mem<13><2> ), .B(n46), .Y(n1619) );
  OAI21X1 U1439 ( .A(n1252), .B(n1286), .C(n1619), .Y(n2071) );
  NAND2X1 U1440 ( .A(\mem<13><3> ), .B(n46), .Y(n1620) );
  OAI21X1 U1441 ( .A(n1252), .B(n1288), .C(n1620), .Y(n2070) );
  NAND2X1 U1442 ( .A(\mem<13><4> ), .B(n46), .Y(n1621) );
  OAI21X1 U1443 ( .A(n1252), .B(n1290), .C(n1621), .Y(n2069) );
  NAND2X1 U1444 ( .A(\mem<13><5> ), .B(n46), .Y(n1622) );
  OAI21X1 U1445 ( .A(n1252), .B(n1292), .C(n1622), .Y(n2068) );
  NAND2X1 U1446 ( .A(\mem<13><6> ), .B(n46), .Y(n1623) );
  OAI21X1 U1447 ( .A(n1252), .B(n1294), .C(n1623), .Y(n2067) );
  NAND2X1 U1448 ( .A(\mem<13><7> ), .B(n46), .Y(n1624) );
  OAI21X1 U1449 ( .A(n1252), .B(n1296), .C(n1624), .Y(n2066) );
  NAND2X1 U1450 ( .A(\mem<13><8> ), .B(n46), .Y(n1625) );
  OAI21X1 U1451 ( .A(n1253), .B(n1298), .C(n1625), .Y(n2065) );
  NAND2X1 U1452 ( .A(\mem<13><9> ), .B(n46), .Y(n1626) );
  OAI21X1 U1453 ( .A(n1253), .B(n1300), .C(n1626), .Y(n2064) );
  NAND2X1 U1454 ( .A(\mem<13><10> ), .B(n46), .Y(n1627) );
  OAI21X1 U1455 ( .A(n1253), .B(n1302), .C(n1627), .Y(n2063) );
  NAND2X1 U1456 ( .A(\mem<13><11> ), .B(n46), .Y(n1628) );
  OAI21X1 U1457 ( .A(n1253), .B(n1304), .C(n1628), .Y(n2062) );
  NAND2X1 U1458 ( .A(\mem<13><12> ), .B(n46), .Y(n1629) );
  OAI21X1 U1459 ( .A(n1253), .B(n1305), .C(n1629), .Y(n2061) );
  NAND2X1 U1460 ( .A(\mem<13><13> ), .B(n46), .Y(n1630) );
  OAI21X1 U1461 ( .A(n1253), .B(n1307), .C(n1630), .Y(n2060) );
  NAND2X1 U1462 ( .A(\mem<13><14> ), .B(n46), .Y(n1631) );
  OAI21X1 U1463 ( .A(n1253), .B(n1309), .C(n1631), .Y(n2059) );
  NAND2X1 U1464 ( .A(\mem<13><15> ), .B(n46), .Y(n1632) );
  OAI21X1 U1465 ( .A(n1253), .B(n1311), .C(n1632), .Y(n2058) );
  NAND2X1 U1466 ( .A(\mem<12><0> ), .B(n48), .Y(n1633) );
  OAI21X1 U1467 ( .A(n1254), .B(n1282), .C(n1633), .Y(n2057) );
  NAND2X1 U1468 ( .A(\mem<12><1> ), .B(n48), .Y(n1634) );
  OAI21X1 U1469 ( .A(n1254), .B(n1284), .C(n1634), .Y(n2056) );
  NAND2X1 U1470 ( .A(\mem<12><2> ), .B(n48), .Y(n1635) );
  OAI21X1 U1471 ( .A(n1254), .B(n1286), .C(n1635), .Y(n2055) );
  NAND2X1 U1472 ( .A(\mem<12><3> ), .B(n48), .Y(n1636) );
  OAI21X1 U1473 ( .A(n1254), .B(n1288), .C(n1636), .Y(n2054) );
  NAND2X1 U1474 ( .A(\mem<12><4> ), .B(n48), .Y(n1637) );
  OAI21X1 U1475 ( .A(n1254), .B(n1290), .C(n1637), .Y(n2053) );
  NAND2X1 U1476 ( .A(\mem<12><5> ), .B(n48), .Y(n1638) );
  OAI21X1 U1477 ( .A(n1254), .B(n1292), .C(n1638), .Y(n2052) );
  NAND2X1 U1478 ( .A(\mem<12><6> ), .B(n48), .Y(n1639) );
  OAI21X1 U1479 ( .A(n1254), .B(n1294), .C(n1639), .Y(n2051) );
  NAND2X1 U1480 ( .A(\mem<12><7> ), .B(n48), .Y(n1640) );
  OAI21X1 U1481 ( .A(n1254), .B(n1296), .C(n1640), .Y(n2050) );
  NAND2X1 U1482 ( .A(\mem<12><8> ), .B(n48), .Y(n1641) );
  OAI21X1 U1483 ( .A(n1255), .B(n1298), .C(n1641), .Y(n2049) );
  NAND2X1 U1484 ( .A(\mem<12><9> ), .B(n48), .Y(n1642) );
  OAI21X1 U1485 ( .A(n1255), .B(n1300), .C(n1642), .Y(n2048) );
  NAND2X1 U1486 ( .A(\mem<12><10> ), .B(n48), .Y(n1643) );
  OAI21X1 U1487 ( .A(n1255), .B(n1302), .C(n1643), .Y(n2047) );
  NAND2X1 U1488 ( .A(\mem<12><11> ), .B(n48), .Y(n1644) );
  OAI21X1 U1489 ( .A(n1255), .B(n1304), .C(n1644), .Y(n2046) );
  NAND2X1 U1490 ( .A(\mem<12><12> ), .B(n48), .Y(n1645) );
  OAI21X1 U1491 ( .A(n1255), .B(n1305), .C(n1645), .Y(n2045) );
  NAND2X1 U1492 ( .A(\mem<12><13> ), .B(n48), .Y(n1646) );
  OAI21X1 U1493 ( .A(n1255), .B(n1307), .C(n1646), .Y(n2044) );
  NAND2X1 U1494 ( .A(\mem<12><14> ), .B(n48), .Y(n1647) );
  OAI21X1 U1495 ( .A(n1255), .B(n1309), .C(n1647), .Y(n2043) );
  NAND2X1 U1496 ( .A(\mem<12><15> ), .B(n48), .Y(n1648) );
  OAI21X1 U1497 ( .A(n1255), .B(n1311), .C(n1648), .Y(n2042) );
  NAND2X1 U1498 ( .A(\mem<11><0> ), .B(n50), .Y(n1649) );
  OAI21X1 U1499 ( .A(n1256), .B(n1282), .C(n1649), .Y(n2041) );
  NAND2X1 U1500 ( .A(\mem<11><1> ), .B(n50), .Y(n1650) );
  OAI21X1 U1501 ( .A(n1256), .B(n1283), .C(n1650), .Y(n2040) );
  NAND2X1 U1502 ( .A(\mem<11><2> ), .B(n50), .Y(n1651) );
  OAI21X1 U1503 ( .A(n1256), .B(n1285), .C(n1651), .Y(n2039) );
  NAND2X1 U1504 ( .A(\mem<11><3> ), .B(n50), .Y(n1652) );
  OAI21X1 U1505 ( .A(n1256), .B(n1287), .C(n1652), .Y(n2038) );
  NAND2X1 U1506 ( .A(\mem<11><4> ), .B(n50), .Y(n1653) );
  OAI21X1 U1507 ( .A(n1256), .B(n1289), .C(n1653), .Y(n2037) );
  NAND2X1 U1508 ( .A(\mem<11><5> ), .B(n50), .Y(n1654) );
  OAI21X1 U1509 ( .A(n1256), .B(n1291), .C(n1654), .Y(n2036) );
  NAND2X1 U1510 ( .A(\mem<11><6> ), .B(n50), .Y(n1655) );
  OAI21X1 U1511 ( .A(n1256), .B(n1293), .C(n1655), .Y(n2035) );
  NAND2X1 U1512 ( .A(\mem<11><7> ), .B(n50), .Y(n1656) );
  OAI21X1 U1513 ( .A(n1256), .B(n1295), .C(n1656), .Y(n2034) );
  NAND2X1 U1514 ( .A(\mem<11><8> ), .B(n50), .Y(n1657) );
  OAI21X1 U1515 ( .A(n1257), .B(n1297), .C(n1657), .Y(n2033) );
  NAND2X1 U1516 ( .A(\mem<11><9> ), .B(n50), .Y(n1658) );
  OAI21X1 U1517 ( .A(n1257), .B(n1299), .C(n1658), .Y(n2032) );
  NAND2X1 U1518 ( .A(\mem<11><10> ), .B(n50), .Y(n1659) );
  OAI21X1 U1519 ( .A(n1257), .B(n1301), .C(n1659), .Y(n2031) );
  NAND2X1 U1520 ( .A(\mem<11><11> ), .B(n50), .Y(n1660) );
  OAI21X1 U1521 ( .A(n1257), .B(n1303), .C(n1660), .Y(n2030) );
  NAND2X1 U1522 ( .A(\mem<11><12> ), .B(n50), .Y(n1661) );
  OAI21X1 U1523 ( .A(n1257), .B(n1305), .C(n1661), .Y(n2029) );
  NAND2X1 U1524 ( .A(\mem<11><13> ), .B(n50), .Y(n1662) );
  OAI21X1 U1525 ( .A(n1257), .B(n1306), .C(n1662), .Y(n2028) );
  NAND2X1 U1526 ( .A(\mem<11><14> ), .B(n50), .Y(n1663) );
  OAI21X1 U1527 ( .A(n1257), .B(n1308), .C(n1663), .Y(n2027) );
  NAND2X1 U1528 ( .A(\mem<11><15> ), .B(n50), .Y(n1664) );
  OAI21X1 U1529 ( .A(n1257), .B(n1310), .C(n1664), .Y(n2026) );
  NAND2X1 U1530 ( .A(\mem<10><0> ), .B(n52), .Y(n1665) );
  OAI21X1 U1531 ( .A(n1258), .B(n1282), .C(n1665), .Y(n2025) );
  NAND2X1 U1532 ( .A(\mem<10><1> ), .B(n52), .Y(n1666) );
  OAI21X1 U1533 ( .A(n1258), .B(n1283), .C(n1666), .Y(n2024) );
  NAND2X1 U1534 ( .A(\mem<10><2> ), .B(n52), .Y(n1667) );
  OAI21X1 U1535 ( .A(n1258), .B(n1285), .C(n1667), .Y(n2023) );
  NAND2X1 U1536 ( .A(\mem<10><3> ), .B(n52), .Y(n1668) );
  OAI21X1 U1537 ( .A(n1258), .B(n1287), .C(n1668), .Y(n2022) );
  NAND2X1 U1538 ( .A(\mem<10><4> ), .B(n52), .Y(n1669) );
  OAI21X1 U1539 ( .A(n1258), .B(n1289), .C(n1669), .Y(n2021) );
  NAND2X1 U1540 ( .A(\mem<10><5> ), .B(n52), .Y(n1670) );
  OAI21X1 U1541 ( .A(n1258), .B(n1291), .C(n1670), .Y(n2020) );
  NAND2X1 U1542 ( .A(\mem<10><6> ), .B(n52), .Y(n1671) );
  OAI21X1 U1543 ( .A(n1258), .B(n1293), .C(n1671), .Y(n2019) );
  NAND2X1 U1544 ( .A(\mem<10><7> ), .B(n52), .Y(n1672) );
  OAI21X1 U1545 ( .A(n1258), .B(n1295), .C(n1672), .Y(n2018) );
  NAND2X1 U1546 ( .A(\mem<10><8> ), .B(n52), .Y(n1673) );
  OAI21X1 U1547 ( .A(n1259), .B(n1297), .C(n1673), .Y(n2017) );
  NAND2X1 U1548 ( .A(\mem<10><9> ), .B(n52), .Y(n1674) );
  OAI21X1 U1549 ( .A(n1259), .B(n1299), .C(n1674), .Y(n2016) );
  NAND2X1 U1550 ( .A(\mem<10><10> ), .B(n52), .Y(n1675) );
  OAI21X1 U1551 ( .A(n1259), .B(n1301), .C(n1675), .Y(n2015) );
  NAND2X1 U1552 ( .A(\mem<10><11> ), .B(n52), .Y(n1676) );
  OAI21X1 U1553 ( .A(n1259), .B(n1303), .C(n1676), .Y(n2014) );
  NAND2X1 U1554 ( .A(\mem<10><12> ), .B(n52), .Y(n1677) );
  OAI21X1 U1555 ( .A(n1259), .B(n1305), .C(n1677), .Y(n2013) );
  NAND2X1 U1556 ( .A(\mem<10><13> ), .B(n52), .Y(n1678) );
  OAI21X1 U1557 ( .A(n1259), .B(n1306), .C(n1678), .Y(n2012) );
  NAND2X1 U1558 ( .A(\mem<10><14> ), .B(n52), .Y(n1679) );
  OAI21X1 U1559 ( .A(n1259), .B(n1308), .C(n1679), .Y(n2011) );
  NAND2X1 U1560 ( .A(\mem<10><15> ), .B(n52), .Y(n1680) );
  OAI21X1 U1561 ( .A(n1259), .B(n1310), .C(n1680), .Y(n2010) );
  NAND2X1 U1562 ( .A(\mem<9><0> ), .B(n54), .Y(n1681) );
  OAI21X1 U1563 ( .A(n1260), .B(n1282), .C(n1681), .Y(n2009) );
  NAND2X1 U1564 ( .A(\mem<9><1> ), .B(n54), .Y(n1682) );
  OAI21X1 U1565 ( .A(n1260), .B(n1283), .C(n1682), .Y(n2008) );
  NAND2X1 U1566 ( .A(\mem<9><2> ), .B(n54), .Y(n1683) );
  OAI21X1 U1567 ( .A(n1260), .B(n1285), .C(n1683), .Y(n2007) );
  NAND2X1 U1568 ( .A(\mem<9><3> ), .B(n54), .Y(n1684) );
  OAI21X1 U1569 ( .A(n1260), .B(n1287), .C(n1684), .Y(n2006) );
  NAND2X1 U1570 ( .A(\mem<9><4> ), .B(n54), .Y(n1685) );
  OAI21X1 U1571 ( .A(n1260), .B(n1289), .C(n1685), .Y(n2005) );
  NAND2X1 U1572 ( .A(\mem<9><5> ), .B(n54), .Y(n1686) );
  OAI21X1 U1573 ( .A(n1260), .B(n1291), .C(n1686), .Y(n2004) );
  NAND2X1 U1574 ( .A(\mem<9><6> ), .B(n54), .Y(n1687) );
  OAI21X1 U1575 ( .A(n1260), .B(n1293), .C(n1687), .Y(n2003) );
  NAND2X1 U1576 ( .A(\mem<9><7> ), .B(n54), .Y(n1688) );
  OAI21X1 U1577 ( .A(n1260), .B(n1295), .C(n1688), .Y(n2002) );
  NAND2X1 U1578 ( .A(\mem<9><8> ), .B(n54), .Y(n1689) );
  OAI21X1 U1579 ( .A(n1261), .B(n1297), .C(n1689), .Y(n2001) );
  NAND2X1 U1580 ( .A(\mem<9><9> ), .B(n54), .Y(n1690) );
  OAI21X1 U1581 ( .A(n1261), .B(n1299), .C(n1690), .Y(n2000) );
  NAND2X1 U1582 ( .A(\mem<9><10> ), .B(n54), .Y(n1691) );
  OAI21X1 U1583 ( .A(n1261), .B(n1301), .C(n1691), .Y(n1999) );
  NAND2X1 U1584 ( .A(\mem<9><11> ), .B(n54), .Y(n1692) );
  OAI21X1 U1585 ( .A(n1261), .B(n1303), .C(n1692), .Y(n1998) );
  NAND2X1 U1586 ( .A(\mem<9><12> ), .B(n54), .Y(n1693) );
  OAI21X1 U1587 ( .A(n1261), .B(n1305), .C(n1693), .Y(n1997) );
  NAND2X1 U1588 ( .A(\mem<9><13> ), .B(n54), .Y(n1694) );
  OAI21X1 U1589 ( .A(n1261), .B(n1306), .C(n1694), .Y(n1996) );
  NAND2X1 U1590 ( .A(\mem<9><14> ), .B(n54), .Y(n1695) );
  OAI21X1 U1591 ( .A(n1261), .B(n1308), .C(n1695), .Y(n1995) );
  NAND2X1 U1592 ( .A(\mem<9><15> ), .B(n54), .Y(n1696) );
  OAI21X1 U1593 ( .A(n1261), .B(n1310), .C(n1696), .Y(n1994) );
  NAND2X1 U1594 ( .A(\mem<8><0> ), .B(n56), .Y(n1698) );
  OAI21X1 U1595 ( .A(n1262), .B(n1282), .C(n1698), .Y(n1993) );
  NAND2X1 U1596 ( .A(\mem<8><1> ), .B(n56), .Y(n1699) );
  OAI21X1 U1597 ( .A(n1262), .B(n1283), .C(n1699), .Y(n1992) );
  NAND2X1 U1598 ( .A(\mem<8><2> ), .B(n56), .Y(n1700) );
  OAI21X1 U1599 ( .A(n1262), .B(n1285), .C(n1700), .Y(n1991) );
  NAND2X1 U1600 ( .A(\mem<8><3> ), .B(n56), .Y(n1701) );
  OAI21X1 U1601 ( .A(n1262), .B(n1287), .C(n1701), .Y(n1990) );
  NAND2X1 U1602 ( .A(\mem<8><4> ), .B(n56), .Y(n1702) );
  OAI21X1 U1603 ( .A(n1262), .B(n1289), .C(n1702), .Y(n1989) );
  NAND2X1 U1604 ( .A(\mem<8><5> ), .B(n56), .Y(n1703) );
  OAI21X1 U1605 ( .A(n1262), .B(n1291), .C(n1703), .Y(n1988) );
  NAND2X1 U1606 ( .A(\mem<8><6> ), .B(n56), .Y(n1704) );
  OAI21X1 U1607 ( .A(n1262), .B(n1293), .C(n1704), .Y(n1987) );
  NAND2X1 U1608 ( .A(\mem<8><7> ), .B(n56), .Y(n1705) );
  OAI21X1 U1609 ( .A(n1262), .B(n1295), .C(n1705), .Y(n1986) );
  NAND2X1 U1610 ( .A(\mem<8><8> ), .B(n56), .Y(n1706) );
  OAI21X1 U1611 ( .A(n1262), .B(n1297), .C(n1706), .Y(n1985) );
  NAND2X1 U1612 ( .A(\mem<8><9> ), .B(n56), .Y(n1707) );
  OAI21X1 U1613 ( .A(n1262), .B(n1299), .C(n1707), .Y(n1984) );
  NAND2X1 U1614 ( .A(\mem<8><10> ), .B(n56), .Y(n1708) );
  OAI21X1 U1615 ( .A(n1262), .B(n1301), .C(n1708), .Y(n1983) );
  NAND2X1 U1616 ( .A(\mem<8><11> ), .B(n56), .Y(n1709) );
  OAI21X1 U1617 ( .A(n1262), .B(n1303), .C(n1709), .Y(n1982) );
  NAND2X1 U1618 ( .A(\mem<8><12> ), .B(n56), .Y(n1710) );
  OAI21X1 U1619 ( .A(n1262), .B(n1305), .C(n1710), .Y(n1981) );
  NAND2X1 U1620 ( .A(\mem<8><13> ), .B(n56), .Y(n1711) );
  OAI21X1 U1621 ( .A(n1262), .B(n1306), .C(n1711), .Y(n1980) );
  NAND2X1 U1622 ( .A(\mem<8><14> ), .B(n56), .Y(n1712) );
  OAI21X1 U1623 ( .A(n1262), .B(n1308), .C(n1712), .Y(n1979) );
  NAND2X1 U1624 ( .A(\mem<8><15> ), .B(n56), .Y(n1713) );
  OAI21X1 U1625 ( .A(n1262), .B(n1310), .C(n1713), .Y(n1978) );
  NAND3X1 U1626 ( .A(n1320), .B(n2362), .C(n1322), .Y(n1714) );
  NAND2X1 U1627 ( .A(\mem<7><0> ), .B(n58), .Y(n1715) );
  OAI21X1 U1628 ( .A(n1263), .B(n1281), .C(n1715), .Y(n1977) );
  NAND2X1 U1629 ( .A(\mem<7><1> ), .B(n58), .Y(n1716) );
  OAI21X1 U1630 ( .A(n1263), .B(n1283), .C(n1716), .Y(n1976) );
  NAND2X1 U1631 ( .A(\mem<7><2> ), .B(n58), .Y(n1717) );
  OAI21X1 U1632 ( .A(n1263), .B(n1285), .C(n1717), .Y(n1975) );
  NAND2X1 U1633 ( .A(\mem<7><3> ), .B(n58), .Y(n1718) );
  OAI21X1 U1634 ( .A(n1263), .B(n1287), .C(n1718), .Y(n1974) );
  NAND2X1 U1635 ( .A(\mem<7><4> ), .B(n58), .Y(n1719) );
  OAI21X1 U1636 ( .A(n1263), .B(n1289), .C(n1719), .Y(n1973) );
  NAND2X1 U1637 ( .A(\mem<7><5> ), .B(n58), .Y(n1720) );
  OAI21X1 U1638 ( .A(n1263), .B(n1291), .C(n1720), .Y(n1972) );
  NAND2X1 U1639 ( .A(\mem<7><6> ), .B(n58), .Y(n1721) );
  OAI21X1 U1640 ( .A(n1263), .B(n1293), .C(n1721), .Y(n1971) );
  NAND2X1 U1641 ( .A(\mem<7><7> ), .B(n58), .Y(n1722) );
  OAI21X1 U1642 ( .A(n1263), .B(n1295), .C(n1722), .Y(n1970) );
  NAND2X1 U1643 ( .A(\mem<7><8> ), .B(n58), .Y(n1723) );
  OAI21X1 U1644 ( .A(n1264), .B(n1297), .C(n1723), .Y(n1969) );
  NAND2X1 U1645 ( .A(\mem<7><9> ), .B(n58), .Y(n1724) );
  OAI21X1 U1646 ( .A(n1264), .B(n1299), .C(n1724), .Y(n1968) );
  NAND2X1 U1647 ( .A(\mem<7><10> ), .B(n58), .Y(n1725) );
  OAI21X1 U1648 ( .A(n1264), .B(n1301), .C(n1725), .Y(n1967) );
  NAND2X1 U1649 ( .A(\mem<7><11> ), .B(n58), .Y(n1726) );
  OAI21X1 U1650 ( .A(n1264), .B(n1303), .C(n1726), .Y(n1966) );
  NAND2X1 U1651 ( .A(\mem<7><12> ), .B(n58), .Y(n1727) );
  OAI21X1 U1652 ( .A(n1264), .B(n1305), .C(n1727), .Y(n1965) );
  NAND2X1 U1653 ( .A(\mem<7><13> ), .B(n58), .Y(n1728) );
  OAI21X1 U1654 ( .A(n1264), .B(n1306), .C(n1728), .Y(n1964) );
  NAND2X1 U1655 ( .A(\mem<7><14> ), .B(n58), .Y(n1729) );
  OAI21X1 U1656 ( .A(n1264), .B(n1308), .C(n1729), .Y(n1963) );
  NAND2X1 U1657 ( .A(\mem<7><15> ), .B(n58), .Y(n1730) );
  OAI21X1 U1658 ( .A(n1264), .B(n1310), .C(n1730), .Y(n1962) );
  NAND2X1 U1659 ( .A(\mem<6><0> ), .B(n60), .Y(n1731) );
  OAI21X1 U1660 ( .A(n1265), .B(n1281), .C(n1731), .Y(n1961) );
  NAND2X1 U1661 ( .A(\mem<6><1> ), .B(n60), .Y(n1732) );
  OAI21X1 U1662 ( .A(n1265), .B(n1283), .C(n1732), .Y(n1960) );
  NAND2X1 U1663 ( .A(\mem<6><2> ), .B(n60), .Y(n1733) );
  OAI21X1 U1664 ( .A(n1265), .B(n1285), .C(n1733), .Y(n1959) );
  NAND2X1 U1665 ( .A(\mem<6><3> ), .B(n60), .Y(n1734) );
  OAI21X1 U1666 ( .A(n1265), .B(n1287), .C(n1734), .Y(n1958) );
  NAND2X1 U1667 ( .A(\mem<6><4> ), .B(n60), .Y(n1735) );
  OAI21X1 U1668 ( .A(n1265), .B(n1289), .C(n1735), .Y(n1957) );
  NAND2X1 U1669 ( .A(\mem<6><5> ), .B(n60), .Y(n1736) );
  OAI21X1 U1670 ( .A(n1265), .B(n1291), .C(n1736), .Y(n1956) );
  NAND2X1 U1671 ( .A(\mem<6><6> ), .B(n60), .Y(n1737) );
  OAI21X1 U1672 ( .A(n1265), .B(n1293), .C(n1737), .Y(n1955) );
  NAND2X1 U1673 ( .A(\mem<6><7> ), .B(n60), .Y(n1738) );
  OAI21X1 U1674 ( .A(n1265), .B(n1295), .C(n1738), .Y(n1954) );
  NAND2X1 U1675 ( .A(\mem<6><8> ), .B(n60), .Y(n1739) );
  OAI21X1 U1676 ( .A(n1266), .B(n1297), .C(n1739), .Y(n1953) );
  NAND2X1 U1677 ( .A(\mem<6><9> ), .B(n60), .Y(n1740) );
  OAI21X1 U1678 ( .A(n1266), .B(n1299), .C(n1740), .Y(n1952) );
  NAND2X1 U1679 ( .A(\mem<6><10> ), .B(n60), .Y(n1741) );
  OAI21X1 U1680 ( .A(n1266), .B(n1301), .C(n1741), .Y(n1951) );
  NAND2X1 U1681 ( .A(\mem<6><11> ), .B(n60), .Y(n1742) );
  OAI21X1 U1682 ( .A(n1266), .B(n1303), .C(n1742), .Y(n1950) );
  NAND2X1 U1683 ( .A(\mem<6><12> ), .B(n60), .Y(n1743) );
  OAI21X1 U1684 ( .A(n1266), .B(n1305), .C(n1743), .Y(n1949) );
  NAND2X1 U1685 ( .A(\mem<6><13> ), .B(n60), .Y(n1744) );
  OAI21X1 U1686 ( .A(n1266), .B(n1306), .C(n1744), .Y(n1948) );
  NAND2X1 U1687 ( .A(\mem<6><14> ), .B(n60), .Y(n1745) );
  OAI21X1 U1688 ( .A(n1266), .B(n1308), .C(n1745), .Y(n1947) );
  NAND2X1 U1689 ( .A(\mem<6><15> ), .B(n60), .Y(n1746) );
  OAI21X1 U1690 ( .A(n1266), .B(n1310), .C(n1746), .Y(n1946) );
  NAND2X1 U1691 ( .A(\mem<5><0> ), .B(n62), .Y(n1748) );
  OAI21X1 U1692 ( .A(n1267), .B(n1282), .C(n1748), .Y(n1945) );
  NAND2X1 U1693 ( .A(\mem<5><1> ), .B(n62), .Y(n1749) );
  OAI21X1 U1694 ( .A(n1267), .B(n1283), .C(n1749), .Y(n1944) );
  NAND2X1 U1695 ( .A(\mem<5><2> ), .B(n62), .Y(n1750) );
  OAI21X1 U1696 ( .A(n1267), .B(n1285), .C(n1750), .Y(n1943) );
  NAND2X1 U1697 ( .A(\mem<5><3> ), .B(n62), .Y(n1751) );
  OAI21X1 U1698 ( .A(n1267), .B(n1287), .C(n1751), .Y(n1942) );
  NAND2X1 U1699 ( .A(\mem<5><4> ), .B(n62), .Y(n1752) );
  OAI21X1 U1700 ( .A(n1267), .B(n1289), .C(n1752), .Y(n1941) );
  NAND2X1 U1701 ( .A(\mem<5><5> ), .B(n62), .Y(n1753) );
  OAI21X1 U1702 ( .A(n1267), .B(n1291), .C(n1753), .Y(n1940) );
  NAND2X1 U1703 ( .A(\mem<5><6> ), .B(n62), .Y(n1754) );
  OAI21X1 U1704 ( .A(n1267), .B(n1293), .C(n1754), .Y(n1939) );
  NAND2X1 U1705 ( .A(\mem<5><7> ), .B(n62), .Y(n1755) );
  OAI21X1 U1706 ( .A(n1267), .B(n1295), .C(n1755), .Y(n1938) );
  NAND2X1 U1707 ( .A(\mem<5><8> ), .B(n62), .Y(n1756) );
  OAI21X1 U1708 ( .A(n1268), .B(n1297), .C(n1756), .Y(n1937) );
  NAND2X1 U1709 ( .A(\mem<5><9> ), .B(n62), .Y(n1757) );
  OAI21X1 U1710 ( .A(n1268), .B(n1299), .C(n1757), .Y(n1936) );
  NAND2X1 U1711 ( .A(\mem<5><10> ), .B(n62), .Y(n1758) );
  OAI21X1 U1712 ( .A(n1268), .B(n1301), .C(n1758), .Y(n1935) );
  NAND2X1 U1713 ( .A(\mem<5><11> ), .B(n62), .Y(n1759) );
  OAI21X1 U1714 ( .A(n1268), .B(n1303), .C(n1759), .Y(n1934) );
  NAND2X1 U1715 ( .A(\mem<5><12> ), .B(n62), .Y(n1760) );
  OAI21X1 U1716 ( .A(n1268), .B(n1305), .C(n1760), .Y(n1933) );
  NAND2X1 U1717 ( .A(\mem<5><13> ), .B(n62), .Y(n1761) );
  OAI21X1 U1718 ( .A(n1268), .B(n1306), .C(n1761), .Y(n1932) );
  NAND2X1 U1719 ( .A(\mem<5><14> ), .B(n62), .Y(n1762) );
  OAI21X1 U1720 ( .A(n1268), .B(n1308), .C(n1762), .Y(n1931) );
  NAND2X1 U1721 ( .A(\mem<5><15> ), .B(n62), .Y(n1763) );
  OAI21X1 U1722 ( .A(n1268), .B(n1310), .C(n1763), .Y(n1930) );
  NAND2X1 U1723 ( .A(\mem<4><0> ), .B(n64), .Y(n1765) );
  OAI21X1 U1724 ( .A(n1269), .B(n1281), .C(n1765), .Y(n1929) );
  NAND2X1 U1725 ( .A(\mem<4><1> ), .B(n64), .Y(n1766) );
  OAI21X1 U1726 ( .A(n1269), .B(n1283), .C(n1766), .Y(n1928) );
  NAND2X1 U1727 ( .A(\mem<4><2> ), .B(n64), .Y(n1767) );
  OAI21X1 U1728 ( .A(n1269), .B(n1285), .C(n1767), .Y(n1927) );
  NAND2X1 U1729 ( .A(\mem<4><3> ), .B(n64), .Y(n1768) );
  OAI21X1 U1730 ( .A(n1269), .B(n1287), .C(n1768), .Y(n1926) );
  NAND2X1 U1731 ( .A(\mem<4><4> ), .B(n64), .Y(n1769) );
  OAI21X1 U1732 ( .A(n1269), .B(n1289), .C(n1769), .Y(n1925) );
  NAND2X1 U1733 ( .A(\mem<4><5> ), .B(n64), .Y(n1770) );
  OAI21X1 U1734 ( .A(n1269), .B(n1291), .C(n1770), .Y(n1924) );
  NAND2X1 U1735 ( .A(\mem<4><6> ), .B(n64), .Y(n1771) );
  OAI21X1 U1736 ( .A(n1269), .B(n1293), .C(n1771), .Y(n1923) );
  NAND2X1 U1737 ( .A(\mem<4><7> ), .B(n64), .Y(n1772) );
  OAI21X1 U1738 ( .A(n1269), .B(n1295), .C(n1772), .Y(n1922) );
  NAND2X1 U1739 ( .A(\mem<4><8> ), .B(n64), .Y(n1773) );
  OAI21X1 U1740 ( .A(n1270), .B(n1297), .C(n1773), .Y(n1921) );
  NAND2X1 U1741 ( .A(\mem<4><9> ), .B(n64), .Y(n1774) );
  OAI21X1 U1742 ( .A(n1270), .B(n1299), .C(n1774), .Y(n1920) );
  NAND2X1 U1743 ( .A(\mem<4><10> ), .B(n64), .Y(n1775) );
  OAI21X1 U1744 ( .A(n1270), .B(n1301), .C(n1775), .Y(n1919) );
  NAND2X1 U1745 ( .A(\mem<4><11> ), .B(n64), .Y(n1776) );
  OAI21X1 U1746 ( .A(n1270), .B(n1303), .C(n1776), .Y(n1918) );
  NAND2X1 U1747 ( .A(\mem<4><12> ), .B(n64), .Y(n1777) );
  OAI21X1 U1748 ( .A(n1270), .B(n1305), .C(n1777), .Y(n1917) );
  NAND2X1 U1749 ( .A(\mem<4><13> ), .B(n64), .Y(n1778) );
  OAI21X1 U1750 ( .A(n1270), .B(n1306), .C(n1778), .Y(n1916) );
  NAND2X1 U1751 ( .A(\mem<4><14> ), .B(n64), .Y(n1779) );
  OAI21X1 U1752 ( .A(n1270), .B(n1308), .C(n1779), .Y(n1915) );
  NAND2X1 U1753 ( .A(\mem<4><15> ), .B(n64), .Y(n1780) );
  OAI21X1 U1754 ( .A(n1270), .B(n1310), .C(n1780), .Y(n1914) );
  NAND2X1 U1755 ( .A(\mem<3><0> ), .B(n66), .Y(n1782) );
  OAI21X1 U1756 ( .A(n1271), .B(n1282), .C(n1782), .Y(n1913) );
  NAND2X1 U1757 ( .A(\mem<3><1> ), .B(n66), .Y(n1783) );
  OAI21X1 U1758 ( .A(n1271), .B(n1283), .C(n1783), .Y(n1912) );
  NAND2X1 U1759 ( .A(\mem<3><2> ), .B(n66), .Y(n1784) );
  OAI21X1 U1760 ( .A(n1271), .B(n1285), .C(n1784), .Y(n1911) );
  NAND2X1 U1761 ( .A(\mem<3><3> ), .B(n66), .Y(n1785) );
  OAI21X1 U1762 ( .A(n1271), .B(n1287), .C(n1785), .Y(n1910) );
  NAND2X1 U1763 ( .A(\mem<3><4> ), .B(n66), .Y(n1786) );
  OAI21X1 U1764 ( .A(n1271), .B(n1289), .C(n1786), .Y(n1909) );
  NAND2X1 U1765 ( .A(\mem<3><5> ), .B(n66), .Y(n1787) );
  OAI21X1 U1766 ( .A(n1271), .B(n1291), .C(n1787), .Y(n1908) );
  NAND2X1 U1767 ( .A(\mem<3><6> ), .B(n66), .Y(n1788) );
  OAI21X1 U1768 ( .A(n1271), .B(n1293), .C(n1788), .Y(n1907) );
  NAND2X1 U1769 ( .A(\mem<3><7> ), .B(n66), .Y(n1789) );
  OAI21X1 U1770 ( .A(n1271), .B(n1295), .C(n1789), .Y(n1906) );
  NAND2X1 U1771 ( .A(\mem<3><8> ), .B(n66), .Y(n1790) );
  OAI21X1 U1772 ( .A(n1272), .B(n1297), .C(n1790), .Y(n1905) );
  NAND2X1 U1773 ( .A(\mem<3><9> ), .B(n66), .Y(n1791) );
  OAI21X1 U1774 ( .A(n1272), .B(n1299), .C(n1791), .Y(n1904) );
  NAND2X1 U1775 ( .A(\mem<3><10> ), .B(n66), .Y(n1792) );
  OAI21X1 U1776 ( .A(n1272), .B(n1301), .C(n1792), .Y(n1903) );
  NAND2X1 U1777 ( .A(\mem<3><11> ), .B(n66), .Y(n1793) );
  OAI21X1 U1778 ( .A(n1272), .B(n1303), .C(n1793), .Y(n1902) );
  NAND2X1 U1779 ( .A(\mem<3><12> ), .B(n66), .Y(n1794) );
  OAI21X1 U1780 ( .A(n1272), .B(n1305), .C(n1794), .Y(n1901) );
  NAND2X1 U1781 ( .A(\mem<3><13> ), .B(n66), .Y(n1795) );
  OAI21X1 U1782 ( .A(n1272), .B(n1306), .C(n1795), .Y(n1900) );
  NAND2X1 U1783 ( .A(\mem<3><14> ), .B(n66), .Y(n1796) );
  OAI21X1 U1784 ( .A(n1272), .B(n1308), .C(n1796), .Y(n1899) );
  NAND2X1 U1785 ( .A(\mem<3><15> ), .B(n66), .Y(n1797) );
  OAI21X1 U1786 ( .A(n1272), .B(n1310), .C(n1797), .Y(n1898) );
  NAND2X1 U1787 ( .A(\mem<2><0> ), .B(n68), .Y(n1799) );
  OAI21X1 U1788 ( .A(n1273), .B(n1281), .C(n1799), .Y(n1897) );
  NAND2X1 U1789 ( .A(\mem<2><1> ), .B(n68), .Y(n1800) );
  OAI21X1 U1790 ( .A(n1273), .B(n1283), .C(n1800), .Y(n1896) );
  NAND2X1 U1791 ( .A(\mem<2><2> ), .B(n68), .Y(n1801) );
  OAI21X1 U1792 ( .A(n1273), .B(n1285), .C(n1801), .Y(n1895) );
  NAND2X1 U1793 ( .A(\mem<2><3> ), .B(n68), .Y(n1802) );
  OAI21X1 U1794 ( .A(n1273), .B(n1287), .C(n1802), .Y(n1894) );
  NAND2X1 U1795 ( .A(\mem<2><4> ), .B(n68), .Y(n1803) );
  OAI21X1 U1796 ( .A(n1273), .B(n1289), .C(n1803), .Y(n1893) );
  NAND2X1 U1797 ( .A(\mem<2><5> ), .B(n68), .Y(n1804) );
  OAI21X1 U1798 ( .A(n1273), .B(n1291), .C(n1804), .Y(n1892) );
  NAND2X1 U1799 ( .A(\mem<2><6> ), .B(n68), .Y(n1805) );
  OAI21X1 U1800 ( .A(n1273), .B(n1293), .C(n1805), .Y(n1891) );
  NAND2X1 U1801 ( .A(\mem<2><7> ), .B(n68), .Y(n1806) );
  OAI21X1 U1802 ( .A(n1273), .B(n1295), .C(n1806), .Y(n1890) );
  NAND2X1 U1803 ( .A(\mem<2><8> ), .B(n68), .Y(n1807) );
  OAI21X1 U1804 ( .A(n1274), .B(n1297), .C(n1807), .Y(n1889) );
  NAND2X1 U1805 ( .A(\mem<2><9> ), .B(n68), .Y(n1808) );
  OAI21X1 U1806 ( .A(n1274), .B(n1299), .C(n1808), .Y(n1888) );
  NAND2X1 U1807 ( .A(\mem<2><10> ), .B(n68), .Y(n1809) );
  OAI21X1 U1808 ( .A(n1274), .B(n1301), .C(n1809), .Y(n1887) );
  NAND2X1 U1809 ( .A(\mem<2><11> ), .B(n68), .Y(n1810) );
  OAI21X1 U1810 ( .A(n1274), .B(n1303), .C(n1810), .Y(n1886) );
  NAND2X1 U1811 ( .A(\mem<2><12> ), .B(n68), .Y(n1811) );
  OAI21X1 U1812 ( .A(n1274), .B(n1305), .C(n1811), .Y(n1885) );
  NAND2X1 U1813 ( .A(\mem<2><13> ), .B(n68), .Y(n1812) );
  OAI21X1 U1814 ( .A(n1274), .B(n1306), .C(n1812), .Y(n1884) );
  NAND2X1 U1815 ( .A(\mem<2><14> ), .B(n68), .Y(n1813) );
  OAI21X1 U1816 ( .A(n1274), .B(n1308), .C(n1813), .Y(n1883) );
  NAND2X1 U1817 ( .A(\mem<2><15> ), .B(n68), .Y(n1814) );
  OAI21X1 U1818 ( .A(n1274), .B(n1310), .C(n1814), .Y(n1882) );
  NAND2X1 U1819 ( .A(\mem<1><0> ), .B(n70), .Y(n1816) );
  OAI21X1 U1820 ( .A(n1275), .B(n1282), .C(n1816), .Y(n1881) );
  NAND2X1 U1821 ( .A(\mem<1><1> ), .B(n70), .Y(n1817) );
  OAI21X1 U1822 ( .A(n1275), .B(n1283), .C(n1817), .Y(n1880) );
  NAND2X1 U1823 ( .A(\mem<1><2> ), .B(n70), .Y(n1818) );
  OAI21X1 U1824 ( .A(n1275), .B(n1285), .C(n1818), .Y(n1879) );
  NAND2X1 U1825 ( .A(\mem<1><3> ), .B(n70), .Y(n1819) );
  OAI21X1 U1826 ( .A(n1275), .B(n1287), .C(n1819), .Y(n1878) );
  NAND2X1 U1827 ( .A(\mem<1><4> ), .B(n70), .Y(n1820) );
  OAI21X1 U1828 ( .A(n1275), .B(n1289), .C(n1820), .Y(n1877) );
  NAND2X1 U1829 ( .A(\mem<1><5> ), .B(n70), .Y(n1821) );
  OAI21X1 U1830 ( .A(n1275), .B(n1291), .C(n1821), .Y(n1876) );
  NAND2X1 U1831 ( .A(\mem<1><6> ), .B(n70), .Y(n1822) );
  OAI21X1 U1832 ( .A(n1275), .B(n1293), .C(n1822), .Y(n1875) );
  NAND2X1 U1833 ( .A(\mem<1><7> ), .B(n70), .Y(n1823) );
  OAI21X1 U1834 ( .A(n1275), .B(n1295), .C(n1823), .Y(n1874) );
  NAND2X1 U1835 ( .A(\mem<1><8> ), .B(n70), .Y(n1824) );
  OAI21X1 U1836 ( .A(n1276), .B(n1297), .C(n1824), .Y(n1873) );
  NAND2X1 U1837 ( .A(\mem<1><9> ), .B(n70), .Y(n1825) );
  OAI21X1 U1838 ( .A(n1276), .B(n1299), .C(n1825), .Y(n1872) );
  NAND2X1 U1839 ( .A(\mem<1><10> ), .B(n70), .Y(n1826) );
  OAI21X1 U1840 ( .A(n1276), .B(n1301), .C(n1826), .Y(n1871) );
  NAND2X1 U1841 ( .A(\mem<1><11> ), .B(n70), .Y(n1827) );
  OAI21X1 U1842 ( .A(n1276), .B(n1303), .C(n1827), .Y(n1870) );
  NAND2X1 U1843 ( .A(\mem<1><12> ), .B(n70), .Y(n1828) );
  OAI21X1 U1844 ( .A(n1276), .B(n1305), .C(n1828), .Y(n1869) );
  NAND2X1 U1845 ( .A(\mem<1><13> ), .B(n70), .Y(n1829) );
  OAI21X1 U1846 ( .A(n1276), .B(n1306), .C(n1829), .Y(n1868) );
  NAND2X1 U1847 ( .A(\mem<1><14> ), .B(n70), .Y(n1830) );
  OAI21X1 U1848 ( .A(n1276), .B(n1308), .C(n1830), .Y(n1867) );
  NAND2X1 U1849 ( .A(\mem<1><15> ), .B(n70), .Y(n1831) );
  OAI21X1 U1850 ( .A(n1276), .B(n1310), .C(n1831), .Y(n1866) );
  NAND2X1 U1851 ( .A(\mem<0><0> ), .B(n72), .Y(n1834) );
  OAI21X1 U1852 ( .A(n1277), .B(n1282), .C(n1834), .Y(n1865) );
  NAND2X1 U1853 ( .A(\mem<0><1> ), .B(n72), .Y(n1835) );
  OAI21X1 U1854 ( .A(n1277), .B(n1283), .C(n1835), .Y(n1864) );
  NAND2X1 U1855 ( .A(\mem<0><2> ), .B(n72), .Y(n1836) );
  OAI21X1 U1856 ( .A(n1277), .B(n1285), .C(n1836), .Y(n1863) );
  NAND2X1 U1857 ( .A(\mem<0><3> ), .B(n72), .Y(n1837) );
  OAI21X1 U1858 ( .A(n1277), .B(n1287), .C(n1837), .Y(n1862) );
  NAND2X1 U1859 ( .A(\mem<0><4> ), .B(n72), .Y(n1838) );
  OAI21X1 U1860 ( .A(n1277), .B(n1289), .C(n1838), .Y(n1861) );
  NAND2X1 U1861 ( .A(\mem<0><5> ), .B(n72), .Y(n1839) );
  OAI21X1 U1862 ( .A(n1277), .B(n1291), .C(n1839), .Y(n1860) );
  NAND2X1 U1863 ( .A(\mem<0><6> ), .B(n72), .Y(n1840) );
  OAI21X1 U1864 ( .A(n1277), .B(n1293), .C(n1840), .Y(n1859) );
  NAND2X1 U1865 ( .A(\mem<0><7> ), .B(n72), .Y(n1841) );
  OAI21X1 U1866 ( .A(n1277), .B(n1295), .C(n1841), .Y(n1858) );
  NAND2X1 U1867 ( .A(\mem<0><8> ), .B(n72), .Y(n1842) );
  OAI21X1 U1868 ( .A(n1277), .B(n1297), .C(n1842), .Y(n1857) );
  NAND2X1 U1869 ( .A(\mem<0><9> ), .B(n72), .Y(n1843) );
  OAI21X1 U1870 ( .A(n1277), .B(n1299), .C(n1843), .Y(n1856) );
  NAND2X1 U1871 ( .A(\mem<0><10> ), .B(n72), .Y(n1844) );
  OAI21X1 U1872 ( .A(n1277), .B(n1301), .C(n1844), .Y(n1855) );
  NAND2X1 U1873 ( .A(\mem<0><11> ), .B(n72), .Y(n1845) );
  OAI21X1 U1874 ( .A(n1277), .B(n1303), .C(n1845), .Y(n1854) );
  NAND2X1 U1875 ( .A(\mem<0><12> ), .B(n72), .Y(n1846) );
  OAI21X1 U1876 ( .A(n1277), .B(n1305), .C(n1846), .Y(n1853) );
  NAND2X1 U1877 ( .A(\mem<0><13> ), .B(n72), .Y(n1847) );
  OAI21X1 U1878 ( .A(n1277), .B(n1306), .C(n1847), .Y(n1852) );
  NAND2X1 U1879 ( .A(\mem<0><14> ), .B(n72), .Y(n1848) );
  OAI21X1 U1880 ( .A(n1277), .B(n1308), .C(n1848), .Y(n1851) );
  NAND2X1 U1881 ( .A(\mem<0><15> ), .B(n72), .Y(n1849) );
  OAI21X1 U1882 ( .A(n1277), .B(n1310), .C(n1849), .Y(n1850) );
endmodule


module memc_Size16_4 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1911), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1912), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1913), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1914), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1915), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1916), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1917), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1918), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1919), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1920), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1921), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1922), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1923), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1924), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1925), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1926), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1927), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1928), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1929), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1930), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1931), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1932), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1933), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1934), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1935), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1936), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1937), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1938), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1939), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1940), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1941), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1942), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1943), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1944), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1945), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1946), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1947), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1948), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1949), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1950), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1951), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1952), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1953), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1954), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1955), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1956), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1957), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1958), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1959), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1960), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1961), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1962), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1963), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1964), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1965), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1966), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1967), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1968), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1969), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1970), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1971), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1972), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1973), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1974), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1975), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1976), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1977), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1978), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1979), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1980), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1981), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1982), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1983), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1984), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1985), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1986), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1987), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1988), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1989), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1990), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1991), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1992), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1993), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1994), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1995), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1996), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1997), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1998), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1999), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2000), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2001), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2002), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2003), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2004), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2005), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2006), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2007), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2008), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2009), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2010), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2011), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2012), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2013), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2014), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2015), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2016), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2017), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2018), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2019), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2020), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2021), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2022), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2023), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2024), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2025), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2026), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2027), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2028), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2029), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2030), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2031), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2032), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2033), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2034), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2035), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2036), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2037), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2038), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2039), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2040), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2041), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2042), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2043), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2044), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2045), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2046), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2047), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2048), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2049), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2050), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2051), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2052), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2053), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2054), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2055), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2056), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2057), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2058), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2059), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2060), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2061), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2062), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2063), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2064), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2065), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2066), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2067), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2068), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2069), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2070), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2071), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2072), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2073), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2074), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2075), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2076), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2077), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2078), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2079), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2080), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2081), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2082), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2083), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2084), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2085), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2086), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2087), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2088), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2089), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2090), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2091), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2092), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2093), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2094), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2095), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2096), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2097), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2098), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2099), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2100), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2101), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2102), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2103), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2104), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2105), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2106), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2107), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2108), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2109), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2110), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2111), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2112), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2113), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2114), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2115), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2116), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2117), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2118), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2119), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2120), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2121), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2122), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2123), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2124), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2125), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2126), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2127), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2128), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2129), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2130), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2131), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2132), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2133), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2134), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2135), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2136), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2137), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2138), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2139), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2140), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2141), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2142), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2143), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2144), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2145), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2146), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2147), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2148), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2149), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2150), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2151), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2152), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2153), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2154), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2155), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2156), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2157), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2158), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2159), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2160), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2161), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2162), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2163), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2164), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2165), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2166), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2167), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2168), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2169), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2170), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2171), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2172), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2173), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2174), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2175), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2176), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2177), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2178), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2179), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2180), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2181), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2182), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2183), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2184), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2185), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2186), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2187), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2188), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2189), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2190), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2191), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2192), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2193), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2194), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2195), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2196), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2197), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2198), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2199), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2200), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2201), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2202), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2203), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2204), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2205), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2206), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2207), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2208), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2209), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2210), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2211), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2212), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2213), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2214), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2215), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2216), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2217), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2218), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2219), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2220), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2221), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2222), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2223), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2224), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2225), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2226), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2227), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2228), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2229), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2230), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2231), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2232), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2233), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2234), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2235), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2236), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2237), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2238), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2239), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2240), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2241), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2242), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2243), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2244), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2245), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2246), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2247), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2248), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2249), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2250), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2251), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2252), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2253), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2254), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2255), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2256), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2257), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2258), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2259), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2260), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2261), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2262), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2263), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2264), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2265), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2266), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2267), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2268), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2269), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2270), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2271), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2272), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2273), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2274), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2275), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2276), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2277), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2278), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2279), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2280), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2281), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2282), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2283), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2284), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2285), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2286), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2287), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2288), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2289), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2290), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2291), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2292), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2293), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2294), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2295), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2296), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2297), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2298), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2299), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2300), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2301), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2302), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2303), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2304), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2305), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2306), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2307), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2308), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2309), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2310), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2311), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2312), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2313), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2314), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2315), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2316), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2317), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2318), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2319), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2320), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2321), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2322), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2323), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2324), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2325), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2326), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2327), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2328), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2329), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2330), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2331), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2332), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2333), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2334), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2335), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2336), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2337), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2338), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2339), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2340), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2341), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2342), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2343), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2344), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2345), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2346), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2347), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2348), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2349), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2350), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2351), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2352), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2353), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2354), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2355), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2356), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2357), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2358), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2359), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2360), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2361), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2362), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2363), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2364), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2365), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2366), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2367), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2368), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2369), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2370), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2371), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2372), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2373), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2374), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2375), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2376), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2377), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2378), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2379), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2380), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2381), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2382), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2383), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2384), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2385), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2386), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2387), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2388), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2389), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2390), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2391), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2392), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2393), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2394), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2395), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2396), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2397), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2398), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2399), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2400), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2401), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2402), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2403), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2404), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2405), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2406), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2407), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2408), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2409), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2410), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2411), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2412), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2413), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2414), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2415), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2416), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2417), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2418), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2419), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2420), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2421), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2422), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2423) );
  OR2X2 U2 ( .A(n1338), .B(n1319), .Y(n92) );
  INVX1 U3 ( .A(n1214), .Y(n1216) );
  INVX1 U4 ( .A(n1216), .Y(n1191) );
  INVX1 U5 ( .A(n1216), .Y(n1190) );
  INVX1 U6 ( .A(n1216), .Y(n1189) );
  INVX1 U7 ( .A(n1215), .Y(n1188) );
  INVX2 U8 ( .A(n1215), .Y(n1187) );
  INVX1 U9 ( .A(n1191), .Y(n1192) );
  INVX2 U10 ( .A(n1191), .Y(n1193) );
  INVX1 U11 ( .A(n1185), .Y(n1174) );
  INVX2 U12 ( .A(n1191), .Y(n1194) );
  INVX2 U13 ( .A(n1190), .Y(n1195) );
  INVX1 U14 ( .A(n1185), .Y(n1175) );
  INVX2 U15 ( .A(n1190), .Y(n1197) );
  INVX2 U16 ( .A(n1190), .Y(n1196) );
  INVX1 U17 ( .A(n1185), .Y(n1176) );
  INVX2 U18 ( .A(n1189), .Y(n1198) );
  INVX2 U19 ( .A(n1189), .Y(n1199) );
  INVX1 U20 ( .A(n1173), .Y(n1177) );
  INVX2 U21 ( .A(n1189), .Y(n1200) );
  INVX1 U22 ( .A(n1173), .Y(n1178) );
  INVX2 U23 ( .A(n1173), .Y(n1179) );
  INVX1 U24 ( .A(n1172), .Y(n1180) );
  INVX1 U25 ( .A(n1172), .Y(n1181) );
  INVX2 U26 ( .A(n1172), .Y(n1182) );
  INVX2 U27 ( .A(n1173), .Y(n1183) );
  INVX2 U28 ( .A(n1172), .Y(n1184) );
  INVX1 U29 ( .A(n1377), .Y(n1171) );
  INVX1 U30 ( .A(n1377), .Y(n1170) );
  INVX1 U31 ( .A(n1377), .Y(n1169) );
  INVX1 U32 ( .A(n636), .Y(N32) );
  INVX1 U33 ( .A(n637), .Y(N31) );
  INVX1 U34 ( .A(n638), .Y(N30) );
  INVX1 U35 ( .A(n639), .Y(N29) );
  INVX1 U36 ( .A(n640), .Y(N28) );
  INVX1 U37 ( .A(n641), .Y(N27) );
  INVX1 U38 ( .A(n642), .Y(N26) );
  INVX1 U39 ( .A(n643), .Y(N25) );
  INVX1 U40 ( .A(n644), .Y(N24) );
  INVX1 U41 ( .A(n645), .Y(N23) );
  INVX1 U42 ( .A(n646), .Y(N22) );
  INVX1 U43 ( .A(n647), .Y(N21) );
  INVX1 U44 ( .A(n648), .Y(N20) );
  INVX1 U45 ( .A(n649), .Y(N19) );
  INVX1 U46 ( .A(n650), .Y(N18) );
  INVX1 U47 ( .A(n1163), .Y(N17) );
  BUFX2 U48 ( .A(n98), .Y(n1217) );
  BUFX2 U49 ( .A(n100), .Y(n1221) );
  BUFX2 U50 ( .A(n102), .Y(n1225) );
  BUFX2 U51 ( .A(n104), .Y(n1229) );
  BUFX2 U52 ( .A(n106), .Y(n1233) );
  BUFX2 U53 ( .A(n108), .Y(n1237) );
  BUFX2 U54 ( .A(n110), .Y(n1241) );
  BUFX2 U55 ( .A(n112), .Y(n1248) );
  BUFX2 U56 ( .A(n114), .Y(n1252) );
  BUFX2 U57 ( .A(n116), .Y(n1256) );
  BUFX2 U58 ( .A(n118), .Y(n1260) );
  BUFX2 U59 ( .A(n120), .Y(n1264) );
  BUFX2 U60 ( .A(n122), .Y(n1268) );
  BUFX2 U61 ( .A(n124), .Y(n1272) );
  BUFX2 U62 ( .A(n126), .Y(n1277) );
  BUFX2 U63 ( .A(n128), .Y(n1281) );
  BUFX2 U64 ( .A(n130), .Y(n1285) );
  BUFX2 U65 ( .A(n132), .Y(n1289) );
  BUFX2 U66 ( .A(n134), .Y(n1291) );
  BUFX2 U67 ( .A(n136), .Y(n1295) );
  BUFX2 U68 ( .A(n138), .Y(n1299) );
  BUFX2 U69 ( .A(n140), .Y(n1306) );
  BUFX2 U70 ( .A(n142), .Y(n1310) );
  BUFX2 U71 ( .A(n144), .Y(n1314) );
  BUFX2 U72 ( .A(n146), .Y(n1318) );
  BUFX2 U73 ( .A(n146), .Y(n1319) );
  BUFX2 U74 ( .A(n148), .Y(n1320) );
  BUFX2 U75 ( .A(n150), .Y(n1324) );
  BUFX2 U76 ( .A(n152), .Y(n1328) );
  INVX1 U77 ( .A(n1214), .Y(n1215) );
  INVX1 U78 ( .A(n1374), .Y(n1185) );
  INVX1 U79 ( .A(n1379), .Y(n1166) );
  INVX1 U80 ( .A(n1379), .Y(n1165) );
  INVX1 U81 ( .A(n1381), .Y(n1380) );
  INVX1 U82 ( .A(N14), .Y(n1381) );
  INVX1 U83 ( .A(N12), .Y(n1377) );
  INVX1 U84 ( .A(n1377), .Y(n1167) );
  INVX1 U85 ( .A(n1377), .Y(n1168) );
  INVX1 U86 ( .A(n1372), .Y(n1214) );
  INVX2 U87 ( .A(n1372), .Y(n1186) );
  BUFX2 U88 ( .A(n98), .Y(n1218) );
  BUFX2 U89 ( .A(n112), .Y(n1249) );
  INVX1 U90 ( .A(n1379), .Y(n1378) );
  INVX1 U91 ( .A(N13), .Y(n1379) );
  INVX1 U92 ( .A(n94), .Y(n1274) );
  INVX1 U93 ( .A(n95), .Y(n1303) );
  INVX1 U94 ( .A(n96), .Y(n1332) );
  INVX1 U95 ( .A(n93), .Y(n1245) );
  BUFX2 U96 ( .A(n100), .Y(n1222) );
  BUFX2 U97 ( .A(n114), .Y(n1253) );
  BUFX2 U98 ( .A(n116), .Y(n1257) );
  BUFX2 U99 ( .A(n118), .Y(n1261) );
  BUFX2 U100 ( .A(n120), .Y(n1265) );
  BUFX2 U101 ( .A(n122), .Y(n1269) );
  BUFX2 U102 ( .A(n102), .Y(n1226) );
  BUFX2 U103 ( .A(n104), .Y(n1230) );
  BUFX2 U104 ( .A(n106), .Y(n1234) );
  BUFX2 U105 ( .A(n108), .Y(n1238) );
  BUFX2 U106 ( .A(n110), .Y(n1242) );
  BUFX2 U107 ( .A(n128), .Y(n1282) );
  BUFX2 U108 ( .A(n130), .Y(n1286) );
  BUFX2 U109 ( .A(n134), .Y(n1292) );
  BUFX2 U110 ( .A(n136), .Y(n1296) );
  BUFX2 U111 ( .A(n138), .Y(n1300) );
  BUFX2 U112 ( .A(n142), .Y(n1311) );
  BUFX2 U113 ( .A(n144), .Y(n1315) );
  BUFX2 U114 ( .A(n148), .Y(n1321) );
  BUFX2 U115 ( .A(n150), .Y(n1325) );
  BUFX2 U116 ( .A(n152), .Y(n1329) );
  BUFX2 U117 ( .A(n126), .Y(n1278) );
  BUFX2 U118 ( .A(n140), .Y(n1307) );
  INVX1 U119 ( .A(n1374), .Y(n1172) );
  INVX1 U120 ( .A(n1374), .Y(n1173) );
  INVX1 U121 ( .A(n1381), .Y(n1164) );
  BUFX2 U122 ( .A(n132), .Y(n1290) );
  BUFX2 U123 ( .A(n124), .Y(n1273) );
  INVX1 U124 ( .A(rst), .Y(n1371) );
  INVX2 U125 ( .A(n3), .Y(n1) );
  INVX2 U126 ( .A(n3), .Y(n2) );
  OR2X2 U127 ( .A(write), .B(rst), .Y(n3) );
  AND2X2 U128 ( .A(\data_in<0> ), .B(n1337), .Y(n4) );
  AND2X2 U129 ( .A(n1335), .B(n97), .Y(n5) );
  INVX1 U130 ( .A(n5), .Y(n6) );
  AND2X2 U131 ( .A(\data_in<1> ), .B(n1337), .Y(n7) );
  AND2X2 U132 ( .A(\data_in<2> ), .B(n1337), .Y(n8) );
  AND2X2 U133 ( .A(\data_in<3> ), .B(n1337), .Y(n9) );
  AND2X2 U134 ( .A(\data_in<4> ), .B(n1337), .Y(n10) );
  AND2X2 U135 ( .A(\data_in<5> ), .B(n1337), .Y(n11) );
  AND2X2 U136 ( .A(\data_in<6> ), .B(n1337), .Y(n12) );
  AND2X2 U137 ( .A(\data_in<7> ), .B(n1337), .Y(n13) );
  AND2X2 U138 ( .A(\data_in<8> ), .B(n1337), .Y(n14) );
  AND2X2 U139 ( .A(\data_in<9> ), .B(n1337), .Y(n15) );
  AND2X2 U140 ( .A(\data_in<10> ), .B(n1337), .Y(n16) );
  AND2X2 U141 ( .A(\data_in<11> ), .B(n1336), .Y(n17) );
  AND2X2 U142 ( .A(\data_in<12> ), .B(n1336), .Y(n18) );
  AND2X2 U143 ( .A(\data_in<13> ), .B(n1336), .Y(n19) );
  AND2X2 U144 ( .A(\data_in<14> ), .B(n1336), .Y(n20) );
  AND2X2 U145 ( .A(\data_in<15> ), .B(n1336), .Y(n21) );
  AND2X2 U146 ( .A(n1337), .B(n99), .Y(n22) );
  INVX1 U147 ( .A(n22), .Y(n23) );
  AND2X2 U148 ( .A(n1336), .B(n101), .Y(n24) );
  INVX1 U149 ( .A(n24), .Y(n25) );
  AND2X2 U150 ( .A(n1335), .B(n103), .Y(n26) );
  INVX1 U151 ( .A(n26), .Y(n27) );
  AND2X2 U152 ( .A(n1337), .B(n105), .Y(n28) );
  INVX1 U153 ( .A(n28), .Y(n29) );
  AND2X2 U154 ( .A(n1336), .B(n107), .Y(n30) );
  INVX1 U155 ( .A(n30), .Y(n31) );
  AND2X2 U156 ( .A(n1335), .B(n109), .Y(n32) );
  INVX1 U157 ( .A(n32), .Y(n33) );
  AND2X2 U158 ( .A(n1337), .B(n93), .Y(n34) );
  INVX1 U159 ( .A(n34), .Y(n35) );
  AND2X2 U160 ( .A(n1337), .B(n111), .Y(n36) );
  INVX1 U161 ( .A(n36), .Y(n37) );
  AND2X2 U162 ( .A(n1336), .B(n113), .Y(n38) );
  INVX1 U163 ( .A(n38), .Y(n39) );
  AND2X2 U164 ( .A(n1335), .B(n115), .Y(n40) );
  INVX1 U165 ( .A(n40), .Y(n41) );
  AND2X2 U166 ( .A(n1337), .B(n117), .Y(n42) );
  INVX1 U167 ( .A(n42), .Y(n43) );
  AND2X2 U168 ( .A(n1335), .B(n119), .Y(n44) );
  INVX1 U169 ( .A(n44), .Y(n45) );
  AND2X2 U170 ( .A(n1335), .B(n121), .Y(n46) );
  INVX1 U171 ( .A(n46), .Y(n47) );
  AND2X2 U172 ( .A(n1335), .B(n94), .Y(n48) );
  INVX1 U173 ( .A(n48), .Y(n49) );
  AND2X2 U174 ( .A(n1335), .B(n125), .Y(n50) );
  INVX1 U175 ( .A(n50), .Y(n51) );
  AND2X2 U176 ( .A(n1335), .B(n127), .Y(n52) );
  INVX1 U177 ( .A(n52), .Y(n53) );
  AND2X2 U178 ( .A(n1335), .B(n129), .Y(n54) );
  INVX1 U179 ( .A(n54), .Y(n55) );
  AND2X2 U180 ( .A(n1335), .B(n133), .Y(n56) );
  INVX1 U181 ( .A(n56), .Y(n57) );
  AND2X2 U182 ( .A(n1335), .B(n135), .Y(n58) );
  INVX1 U183 ( .A(n58), .Y(n59) );
  AND2X2 U184 ( .A(n1335), .B(n137), .Y(n60) );
  INVX1 U185 ( .A(n60), .Y(n61) );
  AND2X2 U186 ( .A(n1336), .B(n95), .Y(n62) );
  INVX1 U187 ( .A(n62), .Y(n63) );
  AND2X2 U188 ( .A(n1336), .B(n139), .Y(n64) );
  INVX1 U189 ( .A(n64), .Y(n65) );
  AND2X2 U190 ( .A(n1336), .B(n141), .Y(n66) );
  INVX1 U191 ( .A(n66), .Y(n67) );
  AND2X2 U192 ( .A(n1336), .B(n143), .Y(n68) );
  INVX1 U193 ( .A(n68), .Y(n69) );
  AND2X2 U194 ( .A(n1336), .B(n147), .Y(n70) );
  INVX1 U195 ( .A(n70), .Y(n71) );
  AND2X2 U196 ( .A(n1336), .B(n149), .Y(n72) );
  INVX1 U197 ( .A(n72), .Y(n73) );
  AND2X2 U198 ( .A(n1336), .B(n151), .Y(n74) );
  INVX1 U199 ( .A(n74), .Y(n75) );
  AND2X2 U200 ( .A(n1335), .B(n96), .Y(n76) );
  INVX1 U201 ( .A(n76), .Y(n77) );
  BUFX2 U202 ( .A(n6), .Y(n1219) );
  BUFX2 U203 ( .A(n6), .Y(n1220) );
  BUFX2 U204 ( .A(n23), .Y(n1223) );
  BUFX2 U205 ( .A(n23), .Y(n1224) );
  BUFX2 U206 ( .A(n25), .Y(n1227) );
  BUFX2 U207 ( .A(n25), .Y(n1228) );
  BUFX2 U208 ( .A(n27), .Y(n1231) );
  BUFX2 U209 ( .A(n27), .Y(n1232) );
  BUFX2 U210 ( .A(n29), .Y(n1235) );
  BUFX2 U211 ( .A(n29), .Y(n1236) );
  BUFX2 U212 ( .A(n31), .Y(n1239) );
  BUFX2 U213 ( .A(n31), .Y(n1240) );
  BUFX2 U214 ( .A(n33), .Y(n1243) );
  BUFX2 U215 ( .A(n33), .Y(n1244) );
  BUFX2 U216 ( .A(n35), .Y(n1246) );
  BUFX2 U217 ( .A(n35), .Y(n1247) );
  BUFX2 U218 ( .A(n37), .Y(n1250) );
  BUFX2 U219 ( .A(n37), .Y(n1251) );
  BUFX2 U220 ( .A(n39), .Y(n1254) );
  BUFX2 U221 ( .A(n39), .Y(n1255) );
  BUFX2 U222 ( .A(n41), .Y(n1258) );
  BUFX2 U223 ( .A(n41), .Y(n1259) );
  BUFX2 U224 ( .A(n43), .Y(n1262) );
  BUFX2 U225 ( .A(n43), .Y(n1263) );
  AND2X2 U226 ( .A(n1371), .B(write), .Y(n78) );
  INVX1 U227 ( .A(n1377), .Y(n1376) );
  INVX1 U228 ( .A(n1373), .Y(n1372) );
  AND2X1 U229 ( .A(n1376), .B(n1374), .Y(n79) );
  INVX1 U230 ( .A(n1375), .Y(n1374) );
  AND2X1 U231 ( .A(n2423), .B(n1380), .Y(n80) );
  INVX2 U232 ( .A(n154), .Y(n1626) );
  INVX2 U233 ( .A(n153), .Y(n1708) );
  BUFX2 U234 ( .A(n1414), .Y(n81) );
  INVX1 U235 ( .A(n81), .Y(n1808) );
  BUFX2 U236 ( .A(n1431), .Y(n82) );
  INVX1 U237 ( .A(n82), .Y(n1825) );
  BUFX2 U238 ( .A(n1448), .Y(n83) );
  INVX1 U239 ( .A(n83), .Y(n1842) );
  BUFX2 U240 ( .A(n1465), .Y(n84) );
  INVX1 U241 ( .A(n84), .Y(n1859) );
  BUFX2 U242 ( .A(n1482), .Y(n85) );
  INVX1 U243 ( .A(n85), .Y(n1876) );
  BUFX2 U244 ( .A(n1644), .Y(n86) );
  INVX1 U245 ( .A(n86), .Y(n1758) );
  BUFX2 U246 ( .A(n1775), .Y(n87) );
  INVX1 U247 ( .A(n87), .Y(n1893) );
  AND2X1 U248 ( .A(n1372), .B(n79), .Y(n88) );
  AND2X1 U249 ( .A(n1378), .B(n80), .Y(n89) );
  AND2X1 U250 ( .A(n1373), .B(n79), .Y(n90) );
  AND2X1 U251 ( .A(n1379), .B(n80), .Y(n91) );
  AND2X1 U252 ( .A(n89), .B(n1894), .Y(n93) );
  AND2X1 U253 ( .A(n1894), .B(n91), .Y(n94) );
  AND2X1 U254 ( .A(n1894), .B(n1758), .Y(n95) );
  AND2X1 U255 ( .A(n1894), .B(n1893), .Y(n96) );
  AND2X1 U256 ( .A(n88), .B(n89), .Y(n97) );
  INVX1 U257 ( .A(n97), .Y(n98) );
  AND2X1 U258 ( .A(n89), .B(n90), .Y(n99) );
  INVX1 U259 ( .A(n99), .Y(n100) );
  AND2X1 U260 ( .A(n89), .B(n1808), .Y(n101) );
  INVX1 U261 ( .A(n101), .Y(n102) );
  AND2X1 U262 ( .A(n89), .B(n1825), .Y(n103) );
  INVX1 U263 ( .A(n103), .Y(n104) );
  AND2X1 U264 ( .A(n89), .B(n1842), .Y(n105) );
  INVX1 U265 ( .A(n105), .Y(n106) );
  AND2X1 U266 ( .A(n89), .B(n1859), .Y(n107) );
  INVX1 U267 ( .A(n107), .Y(n108) );
  AND2X1 U268 ( .A(n89), .B(n1876), .Y(n109) );
  INVX1 U269 ( .A(n109), .Y(n110) );
  AND2X1 U270 ( .A(n88), .B(n91), .Y(n111) );
  INVX1 U271 ( .A(n111), .Y(n112) );
  AND2X1 U272 ( .A(n90), .B(n91), .Y(n113) );
  INVX1 U273 ( .A(n113), .Y(n114) );
  AND2X1 U274 ( .A(n1808), .B(n91), .Y(n115) );
  INVX1 U275 ( .A(n115), .Y(n116) );
  AND2X1 U276 ( .A(n1825), .B(n91), .Y(n117) );
  INVX1 U277 ( .A(n117), .Y(n118) );
  AND2X1 U278 ( .A(n1842), .B(n91), .Y(n119) );
  INVX1 U279 ( .A(n119), .Y(n120) );
  AND2X1 U280 ( .A(n1859), .B(n91), .Y(n121) );
  INVX1 U281 ( .A(n121), .Y(n122) );
  AND2X1 U282 ( .A(n1876), .B(n91), .Y(n123) );
  INVX1 U283 ( .A(n123), .Y(n124) );
  AND2X1 U284 ( .A(n88), .B(n1758), .Y(n125) );
  INVX1 U285 ( .A(n125), .Y(n126) );
  AND2X1 U286 ( .A(n90), .B(n1758), .Y(n127) );
  INVX1 U287 ( .A(n127), .Y(n128) );
  AND2X1 U288 ( .A(n1808), .B(n1758), .Y(n129) );
  INVX1 U289 ( .A(n129), .Y(n130) );
  AND2X1 U290 ( .A(n1825), .B(n1758), .Y(n131) );
  INVX1 U291 ( .A(n131), .Y(n132) );
  AND2X1 U292 ( .A(n1842), .B(n1758), .Y(n133) );
  INVX1 U293 ( .A(n133), .Y(n134) );
  AND2X1 U294 ( .A(n1859), .B(n1758), .Y(n135) );
  INVX1 U295 ( .A(n135), .Y(n136) );
  AND2X1 U296 ( .A(n1876), .B(n1758), .Y(n137) );
  INVX1 U297 ( .A(n137), .Y(n138) );
  AND2X1 U298 ( .A(n88), .B(n1893), .Y(n139) );
  INVX1 U299 ( .A(n139), .Y(n140) );
  AND2X1 U300 ( .A(n90), .B(n1893), .Y(n141) );
  INVX1 U301 ( .A(n141), .Y(n142) );
  AND2X1 U302 ( .A(n1808), .B(n1893), .Y(n143) );
  INVX1 U303 ( .A(n143), .Y(n144) );
  AND2X1 U304 ( .A(n1825), .B(n1893), .Y(n145) );
  INVX1 U305 ( .A(n145), .Y(n146) );
  AND2X1 U306 ( .A(n1842), .B(n1893), .Y(n147) );
  INVX1 U307 ( .A(n147), .Y(n148) );
  AND2X1 U308 ( .A(n1859), .B(n1893), .Y(n149) );
  INVX1 U309 ( .A(n149), .Y(n150) );
  AND2X1 U310 ( .A(n1876), .B(n1893), .Y(n151) );
  INVX1 U311 ( .A(n151), .Y(n152) );
  INVX4 U312 ( .A(n78), .Y(n1338) );
  BUFX2 U313 ( .A(n59), .Y(n1297) );
  BUFX2 U314 ( .A(n73), .Y(n1326) );
  AND2X2 U315 ( .A(n1335), .B(n131), .Y(n153) );
  BUFX2 U316 ( .A(n53), .Y(n1283) );
  AND2X2 U317 ( .A(n1335), .B(n123), .Y(n154) );
  BUFX2 U318 ( .A(n45), .Y(n1266) );
  BUFX2 U319 ( .A(n67), .Y(n1312) );
  BUFX2 U320 ( .A(n77), .Y(n1333) );
  BUFX2 U321 ( .A(n77), .Y(n1334) );
  BUFX2 U322 ( .A(n49), .Y(n1276) );
  BUFX2 U323 ( .A(n49), .Y(n1275) );
  BUFX2 U324 ( .A(n61), .Y(n1301) );
  BUFX2 U325 ( .A(n61), .Y(n1302) );
  BUFX2 U326 ( .A(n59), .Y(n1298) );
  BUFX2 U327 ( .A(n57), .Y(n1293) );
  BUFX2 U328 ( .A(n57), .Y(n1294) );
  BUFX2 U329 ( .A(n55), .Y(n1287) );
  BUFX2 U330 ( .A(n55), .Y(n1288) );
  BUFX2 U331 ( .A(n53), .Y(n1284) );
  BUFX2 U332 ( .A(n51), .Y(n1279) );
  BUFX2 U333 ( .A(n51), .Y(n1280) );
  BUFX2 U334 ( .A(n47), .Y(n1270) );
  BUFX2 U335 ( .A(n47), .Y(n1271) );
  BUFX2 U336 ( .A(n45), .Y(n1267) );
  BUFX2 U337 ( .A(n63), .Y(n1304) );
  BUFX2 U338 ( .A(n63), .Y(n1305) );
  BUFX2 U339 ( .A(n75), .Y(n1330) );
  BUFX2 U340 ( .A(n75), .Y(n1331) );
  BUFX2 U341 ( .A(n73), .Y(n1327) );
  BUFX2 U342 ( .A(n71), .Y(n1322) );
  BUFX2 U343 ( .A(n71), .Y(n1323) );
  BUFX2 U344 ( .A(n69), .Y(n1316) );
  BUFX2 U345 ( .A(n69), .Y(n1317) );
  BUFX2 U346 ( .A(n67), .Y(n1313) );
  BUFX2 U347 ( .A(n65), .Y(n1308) );
  BUFX2 U348 ( .A(n65), .Y(n1309) );
  MUX2X1 U349 ( .B(n156), .A(n157), .S(n1174), .Y(n155) );
  MUX2X1 U350 ( .B(n159), .A(n160), .S(n1174), .Y(n158) );
  MUX2X1 U351 ( .B(n162), .A(n163), .S(n1174), .Y(n161) );
  MUX2X1 U352 ( .B(n165), .A(n166), .S(n1174), .Y(n164) );
  MUX2X1 U353 ( .B(n168), .A(n169), .S(n1166), .Y(n167) );
  MUX2X1 U354 ( .B(n171), .A(n172), .S(n1174), .Y(n170) );
  MUX2X1 U355 ( .B(n174), .A(n175), .S(n1174), .Y(n173) );
  MUX2X1 U356 ( .B(n177), .A(n178), .S(n1174), .Y(n176) );
  MUX2X1 U357 ( .B(n180), .A(n181), .S(n1174), .Y(n179) );
  MUX2X1 U358 ( .B(n183), .A(n184), .S(n1166), .Y(n182) );
  MUX2X1 U359 ( .B(n186), .A(n187), .S(n1175), .Y(n185) );
  MUX2X1 U360 ( .B(n189), .A(n190), .S(n1175), .Y(n188) );
  MUX2X1 U361 ( .B(n192), .A(n193), .S(n1175), .Y(n191) );
  MUX2X1 U362 ( .B(n195), .A(n196), .S(n1175), .Y(n194) );
  MUX2X1 U363 ( .B(n198), .A(n199), .S(n1166), .Y(n197) );
  MUX2X1 U364 ( .B(n201), .A(n202), .S(n1175), .Y(n200) );
  MUX2X1 U365 ( .B(n204), .A(n205), .S(n1175), .Y(n203) );
  MUX2X1 U366 ( .B(n207), .A(n208), .S(n1175), .Y(n206) );
  MUX2X1 U367 ( .B(n210), .A(n211), .S(n1175), .Y(n209) );
  MUX2X1 U368 ( .B(n213), .A(n215), .S(n1166), .Y(n212) );
  MUX2X1 U369 ( .B(n217), .A(n218), .S(n1175), .Y(n216) );
  MUX2X1 U370 ( .B(n220), .A(n221), .S(n1175), .Y(n219) );
  MUX2X1 U371 ( .B(n223), .A(n224), .S(n1175), .Y(n222) );
  MUX2X1 U372 ( .B(n226), .A(n227), .S(n1175), .Y(n225) );
  MUX2X1 U373 ( .B(n229), .A(n230), .S(n1166), .Y(n228) );
  MUX2X1 U374 ( .B(n232), .A(n233), .S(n1176), .Y(n231) );
  MUX2X1 U375 ( .B(n235), .A(n236), .S(n1176), .Y(n234) );
  MUX2X1 U376 ( .B(n238), .A(n239), .S(n1176), .Y(n237) );
  MUX2X1 U377 ( .B(n241), .A(n242), .S(n1176), .Y(n240) );
  MUX2X1 U378 ( .B(n244), .A(n245), .S(n1166), .Y(n243) );
  MUX2X1 U379 ( .B(n247), .A(n248), .S(n1176), .Y(n246) );
  MUX2X1 U380 ( .B(n250), .A(n251), .S(n1176), .Y(n249) );
  MUX2X1 U381 ( .B(n253), .A(n254), .S(n1176), .Y(n252) );
  MUX2X1 U382 ( .B(n256), .A(n257), .S(n1176), .Y(n255) );
  MUX2X1 U383 ( .B(n259), .A(n260), .S(n1166), .Y(n258) );
  MUX2X1 U384 ( .B(n262), .A(n263), .S(n1176), .Y(n261) );
  MUX2X1 U385 ( .B(n265), .A(n266), .S(n1176), .Y(n264) );
  MUX2X1 U386 ( .B(n268), .A(n269), .S(n1176), .Y(n267) );
  MUX2X1 U387 ( .B(n271), .A(n272), .S(n1176), .Y(n270) );
  MUX2X1 U388 ( .B(n274), .A(n275), .S(n1166), .Y(n273) );
  MUX2X1 U389 ( .B(n277), .A(n278), .S(n1177), .Y(n276) );
  MUX2X1 U390 ( .B(n280), .A(n281), .S(n1177), .Y(n279) );
  MUX2X1 U391 ( .B(n283), .A(n284), .S(n1177), .Y(n282) );
  MUX2X1 U392 ( .B(n286), .A(n287), .S(n1177), .Y(n285) );
  MUX2X1 U393 ( .B(n289), .A(n290), .S(n1166), .Y(n288) );
  MUX2X1 U394 ( .B(n292), .A(n293), .S(n1177), .Y(n291) );
  MUX2X1 U395 ( .B(n295), .A(n296), .S(n1177), .Y(n294) );
  MUX2X1 U396 ( .B(n298), .A(n299), .S(n1177), .Y(n297) );
  MUX2X1 U397 ( .B(n301), .A(n302), .S(n1177), .Y(n300) );
  MUX2X1 U398 ( .B(n304), .A(n305), .S(n1166), .Y(n303) );
  MUX2X1 U399 ( .B(n307), .A(n308), .S(n1177), .Y(n306) );
  MUX2X1 U400 ( .B(n310), .A(n311), .S(n1177), .Y(n309) );
  MUX2X1 U401 ( .B(n313), .A(n314), .S(n1177), .Y(n312) );
  MUX2X1 U402 ( .B(n316), .A(n317), .S(n1177), .Y(n315) );
  MUX2X1 U403 ( .B(n319), .A(n320), .S(n1166), .Y(n318) );
  MUX2X1 U404 ( .B(n322), .A(n323), .S(n1178), .Y(n321) );
  MUX2X1 U405 ( .B(n325), .A(n326), .S(n1178), .Y(n324) );
  MUX2X1 U406 ( .B(n328), .A(n329), .S(n1178), .Y(n327) );
  MUX2X1 U407 ( .B(n331), .A(n332), .S(n1178), .Y(n330) );
  MUX2X1 U408 ( .B(n334), .A(n335), .S(n1166), .Y(n333) );
  MUX2X1 U409 ( .B(n337), .A(n338), .S(n1178), .Y(n336) );
  MUX2X1 U410 ( .B(n340), .A(n341), .S(n1178), .Y(n339) );
  MUX2X1 U411 ( .B(n343), .A(n344), .S(n1178), .Y(n342) );
  MUX2X1 U412 ( .B(n346), .A(n347), .S(n1178), .Y(n345) );
  MUX2X1 U413 ( .B(n349), .A(n350), .S(n1165), .Y(n348) );
  MUX2X1 U414 ( .B(n352), .A(n353), .S(n1178), .Y(n351) );
  MUX2X1 U415 ( .B(n355), .A(n356), .S(n1178), .Y(n354) );
  MUX2X1 U416 ( .B(n358), .A(n359), .S(n1178), .Y(n357) );
  MUX2X1 U417 ( .B(n361), .A(n362), .S(n1178), .Y(n360) );
  MUX2X1 U418 ( .B(n364), .A(n365), .S(n1165), .Y(n363) );
  MUX2X1 U419 ( .B(n367), .A(n368), .S(n1179), .Y(n366) );
  MUX2X1 U420 ( .B(n370), .A(n371), .S(n1179), .Y(n369) );
  MUX2X1 U421 ( .B(n373), .A(n374), .S(n1179), .Y(n372) );
  MUX2X1 U422 ( .B(n376), .A(n377), .S(n1179), .Y(n375) );
  MUX2X1 U423 ( .B(n379), .A(n380), .S(n1165), .Y(n378) );
  MUX2X1 U424 ( .B(n382), .A(n383), .S(n1179), .Y(n381) );
  MUX2X1 U425 ( .B(n385), .A(n386), .S(n1179), .Y(n384) );
  MUX2X1 U426 ( .B(n388), .A(n389), .S(n1179), .Y(n387) );
  MUX2X1 U427 ( .B(n391), .A(n392), .S(n1179), .Y(n390) );
  MUX2X1 U428 ( .B(n394), .A(n395), .S(n1165), .Y(n393) );
  MUX2X1 U429 ( .B(n397), .A(n398), .S(n1179), .Y(n396) );
  MUX2X1 U430 ( .B(n400), .A(n401), .S(n1179), .Y(n399) );
  MUX2X1 U431 ( .B(n403), .A(n404), .S(n1179), .Y(n402) );
  MUX2X1 U432 ( .B(n406), .A(n407), .S(n1179), .Y(n405) );
  MUX2X1 U433 ( .B(n409), .A(n410), .S(n1165), .Y(n408) );
  MUX2X1 U434 ( .B(n412), .A(n413), .S(n1180), .Y(n411) );
  MUX2X1 U435 ( .B(n415), .A(n416), .S(n1180), .Y(n414) );
  MUX2X1 U436 ( .B(n418), .A(n419), .S(n1180), .Y(n417) );
  MUX2X1 U437 ( .B(n421), .A(n422), .S(n1180), .Y(n420) );
  MUX2X1 U438 ( .B(n424), .A(n425), .S(n1165), .Y(n423) );
  MUX2X1 U439 ( .B(n427), .A(n428), .S(n1180), .Y(n426) );
  MUX2X1 U440 ( .B(n430), .A(n431), .S(n1180), .Y(n429) );
  MUX2X1 U441 ( .B(n433), .A(n434), .S(n1180), .Y(n432) );
  MUX2X1 U442 ( .B(n436), .A(n437), .S(n1180), .Y(n435) );
  MUX2X1 U443 ( .B(n439), .A(n440), .S(n1165), .Y(n438) );
  MUX2X1 U444 ( .B(n442), .A(n443), .S(n1180), .Y(n441) );
  MUX2X1 U445 ( .B(n445), .A(n446), .S(n1180), .Y(n444) );
  MUX2X1 U446 ( .B(n448), .A(n449), .S(n1180), .Y(n447) );
  MUX2X1 U447 ( .B(n451), .A(n452), .S(n1180), .Y(n450) );
  MUX2X1 U448 ( .B(n454), .A(n455), .S(n1165), .Y(n453) );
  MUX2X1 U449 ( .B(n457), .A(n458), .S(n1181), .Y(n456) );
  MUX2X1 U450 ( .B(n460), .A(n461), .S(n1181), .Y(n459) );
  MUX2X1 U451 ( .B(n463), .A(n464), .S(n1181), .Y(n462) );
  MUX2X1 U452 ( .B(n466), .A(n467), .S(n1181), .Y(n465) );
  MUX2X1 U453 ( .B(n469), .A(n470), .S(n1165), .Y(n468) );
  MUX2X1 U454 ( .B(n472), .A(n473), .S(n1181), .Y(n471) );
  MUX2X1 U455 ( .B(n475), .A(n476), .S(n1181), .Y(n474) );
  MUX2X1 U456 ( .B(n478), .A(n479), .S(n1181), .Y(n477) );
  MUX2X1 U457 ( .B(n481), .A(n482), .S(n1181), .Y(n480) );
  MUX2X1 U458 ( .B(n484), .A(n485), .S(n1165), .Y(n483) );
  MUX2X1 U459 ( .B(n487), .A(n488), .S(n1181), .Y(n486) );
  MUX2X1 U460 ( .B(n490), .A(n491), .S(n1181), .Y(n489) );
  MUX2X1 U461 ( .B(n493), .A(n494), .S(n1181), .Y(n492) );
  MUX2X1 U462 ( .B(n496), .A(n497), .S(n1181), .Y(n495) );
  MUX2X1 U463 ( .B(n499), .A(n500), .S(n1165), .Y(n498) );
  MUX2X1 U464 ( .B(n502), .A(n503), .S(n1182), .Y(n501) );
  MUX2X1 U465 ( .B(n505), .A(n506), .S(n1182), .Y(n504) );
  MUX2X1 U466 ( .B(n508), .A(n509), .S(n1182), .Y(n507) );
  MUX2X1 U467 ( .B(n511), .A(n512), .S(n1182), .Y(n510) );
  MUX2X1 U468 ( .B(n514), .A(n515), .S(n1165), .Y(n513) );
  MUX2X1 U469 ( .B(n517), .A(n518), .S(n1182), .Y(n516) );
  MUX2X1 U470 ( .B(n520), .A(n521), .S(n1182), .Y(n519) );
  MUX2X1 U471 ( .B(n523), .A(n524), .S(n1182), .Y(n522) );
  MUX2X1 U472 ( .B(n526), .A(n527), .S(n1182), .Y(n525) );
  MUX2X1 U473 ( .B(n529), .A(n530), .S(n1166), .Y(n528) );
  MUX2X1 U474 ( .B(n532), .A(n533), .S(n1182), .Y(n531) );
  MUX2X1 U475 ( .B(n535), .A(n536), .S(n1182), .Y(n534) );
  MUX2X1 U476 ( .B(n538), .A(n539), .S(n1182), .Y(n537) );
  MUX2X1 U477 ( .B(n541), .A(n542), .S(n1182), .Y(n540) );
  MUX2X1 U478 ( .B(n544), .A(n545), .S(n1166), .Y(n543) );
  MUX2X1 U479 ( .B(n547), .A(n548), .S(n1183), .Y(n546) );
  MUX2X1 U480 ( .B(n550), .A(n551), .S(n1183), .Y(n549) );
  MUX2X1 U481 ( .B(n553), .A(n554), .S(n1183), .Y(n552) );
  MUX2X1 U482 ( .B(n556), .A(n557), .S(n1183), .Y(n555) );
  MUX2X1 U483 ( .B(n559), .A(n560), .S(n1165), .Y(n558) );
  MUX2X1 U484 ( .B(n562), .A(n563), .S(n1183), .Y(n561) );
  MUX2X1 U485 ( .B(n565), .A(n566), .S(n1183), .Y(n564) );
  MUX2X1 U486 ( .B(n568), .A(n569), .S(n1183), .Y(n567) );
  MUX2X1 U487 ( .B(n571), .A(n572), .S(n1183), .Y(n570) );
  MUX2X1 U488 ( .B(n574), .A(n575), .S(n1165), .Y(n573) );
  MUX2X1 U489 ( .B(n577), .A(n578), .S(n1183), .Y(n576) );
  MUX2X1 U490 ( .B(n580), .A(n581), .S(n1183), .Y(n579) );
  MUX2X1 U491 ( .B(n583), .A(n584), .S(n1183), .Y(n582) );
  MUX2X1 U492 ( .B(n586), .A(n587), .S(n1183), .Y(n585) );
  MUX2X1 U493 ( .B(n589), .A(n590), .S(n1166), .Y(n588) );
  MUX2X1 U494 ( .B(n592), .A(n593), .S(n1184), .Y(n591) );
  MUX2X1 U495 ( .B(n595), .A(n596), .S(n1184), .Y(n594) );
  MUX2X1 U496 ( .B(n598), .A(n599), .S(n1184), .Y(n597) );
  MUX2X1 U497 ( .B(n601), .A(n602), .S(n1184), .Y(n600) );
  MUX2X1 U498 ( .B(n604), .A(n605), .S(n1166), .Y(n603) );
  MUX2X1 U499 ( .B(n607), .A(n608), .S(n1184), .Y(n606) );
  MUX2X1 U500 ( .B(n610), .A(n611), .S(n1184), .Y(n609) );
  MUX2X1 U501 ( .B(n613), .A(n614), .S(n1184), .Y(n612) );
  MUX2X1 U502 ( .B(n616), .A(n617), .S(n1184), .Y(n615) );
  MUX2X1 U503 ( .B(n619), .A(n620), .S(n1165), .Y(n618) );
  MUX2X1 U504 ( .B(n622), .A(n623), .S(n1184), .Y(n621) );
  MUX2X1 U505 ( .B(n625), .A(n626), .S(n1184), .Y(n624) );
  MUX2X1 U506 ( .B(n628), .A(n629), .S(n1184), .Y(n627) );
  MUX2X1 U507 ( .B(n631), .A(n632), .S(n1184), .Y(n630) );
  MUX2X1 U508 ( .B(n634), .A(n635), .S(n1165), .Y(n633) );
  MUX2X1 U509 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1192), .Y(n157) );
  MUX2X1 U510 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1192), .Y(n156) );
  MUX2X1 U511 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1192), .Y(n160) );
  MUX2X1 U512 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1192), .Y(n159) );
  MUX2X1 U513 ( .B(n158), .A(n155), .S(n1171), .Y(n169) );
  MUX2X1 U514 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1193), .Y(n163) );
  MUX2X1 U515 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1193), .Y(n162) );
  MUX2X1 U516 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1193), .Y(n166) );
  MUX2X1 U517 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1193), .Y(n165) );
  MUX2X1 U518 ( .B(n164), .A(n161), .S(n1171), .Y(n168) );
  MUX2X1 U519 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1193), .Y(n172) );
  MUX2X1 U520 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1193), .Y(n171) );
  MUX2X1 U521 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1193), .Y(n175) );
  MUX2X1 U522 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1193), .Y(n174) );
  MUX2X1 U523 ( .B(n173), .A(n170), .S(n1171), .Y(n184) );
  MUX2X1 U524 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1193), .Y(n178) );
  MUX2X1 U525 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1193), .Y(n177) );
  MUX2X1 U526 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1193), .Y(n181) );
  MUX2X1 U527 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1193), .Y(n180) );
  MUX2X1 U528 ( .B(n179), .A(n176), .S(n1171), .Y(n183) );
  MUX2X1 U529 ( .B(n182), .A(n167), .S(n1164), .Y(n636) );
  MUX2X1 U530 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1194), .Y(n187) );
  MUX2X1 U531 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1194), .Y(n186) );
  MUX2X1 U532 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1194), .Y(n190) );
  MUX2X1 U533 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1194), .Y(n189) );
  MUX2X1 U534 ( .B(n188), .A(n185), .S(n1171), .Y(n199) );
  MUX2X1 U535 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1194), .Y(n193) );
  MUX2X1 U536 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1194), .Y(n192) );
  MUX2X1 U537 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1194), .Y(n196) );
  MUX2X1 U538 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1194), .Y(n195) );
  MUX2X1 U539 ( .B(n194), .A(n191), .S(n1171), .Y(n198) );
  MUX2X1 U540 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1194), .Y(n202) );
  MUX2X1 U541 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1194), .Y(n201) );
  MUX2X1 U542 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1194), .Y(n205) );
  MUX2X1 U543 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1194), .Y(n204) );
  MUX2X1 U544 ( .B(n203), .A(n200), .S(n1171), .Y(n215) );
  MUX2X1 U545 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1195), .Y(n208) );
  MUX2X1 U546 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1195), .Y(n207) );
  MUX2X1 U547 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1195), .Y(n211) );
  MUX2X1 U548 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1195), .Y(n210) );
  MUX2X1 U549 ( .B(n209), .A(n206), .S(n1171), .Y(n213) );
  MUX2X1 U550 ( .B(n212), .A(n197), .S(n1164), .Y(n637) );
  MUX2X1 U551 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1195), .Y(n218) );
  MUX2X1 U552 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1195), .Y(n217) );
  MUX2X1 U553 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1195), .Y(n221) );
  MUX2X1 U554 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1195), .Y(n220) );
  MUX2X1 U555 ( .B(n219), .A(n216), .S(n1171), .Y(n230) );
  MUX2X1 U556 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1195), .Y(n224) );
  MUX2X1 U557 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1195), .Y(n223) );
  MUX2X1 U558 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1195), .Y(n227) );
  MUX2X1 U559 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1195), .Y(n226) );
  MUX2X1 U560 ( .B(n225), .A(n222), .S(n1171), .Y(n229) );
  MUX2X1 U561 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1196), .Y(n233) );
  MUX2X1 U562 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1196), .Y(n232) );
  MUX2X1 U563 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1196), .Y(n236) );
  MUX2X1 U564 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1196), .Y(n235) );
  MUX2X1 U565 ( .B(n234), .A(n231), .S(n1171), .Y(n245) );
  MUX2X1 U566 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1196), .Y(n239) );
  MUX2X1 U567 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1196), .Y(n238) );
  MUX2X1 U568 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1196), .Y(n242) );
  MUX2X1 U569 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1196), .Y(n241) );
  MUX2X1 U570 ( .B(n240), .A(n237), .S(n1171), .Y(n244) );
  MUX2X1 U571 ( .B(n243), .A(n228), .S(n1164), .Y(n638) );
  MUX2X1 U572 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1196), .Y(n248) );
  MUX2X1 U573 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1196), .Y(n247) );
  MUX2X1 U574 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1196), .Y(n251) );
  MUX2X1 U575 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1196), .Y(n250) );
  MUX2X1 U576 ( .B(n249), .A(n246), .S(n1170), .Y(n260) );
  MUX2X1 U577 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1197), .Y(n254) );
  MUX2X1 U578 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1197), .Y(n253) );
  MUX2X1 U579 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1197), .Y(n257) );
  MUX2X1 U580 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1197), .Y(n256) );
  MUX2X1 U581 ( .B(n255), .A(n252), .S(n1170), .Y(n259) );
  MUX2X1 U582 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1197), .Y(n263) );
  MUX2X1 U583 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1197), .Y(n262) );
  MUX2X1 U584 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1197), .Y(n266) );
  MUX2X1 U585 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1197), .Y(n265) );
  MUX2X1 U586 ( .B(n264), .A(n261), .S(n1170), .Y(n275) );
  MUX2X1 U587 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1197), .Y(n269) );
  MUX2X1 U588 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1197), .Y(n268) );
  MUX2X1 U589 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1197), .Y(n272) );
  MUX2X1 U590 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1197), .Y(n271) );
  MUX2X1 U591 ( .B(n270), .A(n267), .S(n1170), .Y(n274) );
  MUX2X1 U592 ( .B(n273), .A(n258), .S(n1164), .Y(n639) );
  MUX2X1 U593 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1198), .Y(n278) );
  MUX2X1 U594 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1198), .Y(n277) );
  MUX2X1 U595 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1198), .Y(n281) );
  MUX2X1 U596 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1198), .Y(n280) );
  MUX2X1 U597 ( .B(n279), .A(n276), .S(n1170), .Y(n290) );
  MUX2X1 U598 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1198), .Y(n284) );
  MUX2X1 U599 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1198), .Y(n283) );
  MUX2X1 U600 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1198), .Y(n287) );
  MUX2X1 U601 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1198), .Y(n286) );
  MUX2X1 U602 ( .B(n285), .A(n282), .S(n1170), .Y(n289) );
  MUX2X1 U603 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1198), .Y(n293) );
  MUX2X1 U604 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1198), .Y(n292) );
  MUX2X1 U605 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1198), .Y(n296) );
  MUX2X1 U606 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1198), .Y(n295) );
  MUX2X1 U607 ( .B(n294), .A(n291), .S(n1170), .Y(n305) );
  MUX2X1 U608 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1199), .Y(n299) );
  MUX2X1 U609 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1199), .Y(n298) );
  MUX2X1 U610 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1199), .Y(n302) );
  MUX2X1 U611 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1199), .Y(n301) );
  MUX2X1 U612 ( .B(n300), .A(n297), .S(n1170), .Y(n304) );
  MUX2X1 U613 ( .B(n303), .A(n288), .S(n1164), .Y(n640) );
  MUX2X1 U614 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1199), .Y(n308) );
  MUX2X1 U615 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1199), .Y(n307) );
  MUX2X1 U616 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1199), .Y(n311) );
  MUX2X1 U617 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1199), .Y(n310) );
  MUX2X1 U618 ( .B(n309), .A(n306), .S(n1170), .Y(n320) );
  MUX2X1 U619 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1199), .Y(n314) );
  MUX2X1 U620 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1199), .Y(n313) );
  MUX2X1 U621 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1199), .Y(n317) );
  MUX2X1 U622 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1199), .Y(n316) );
  MUX2X1 U623 ( .B(n315), .A(n312), .S(n1170), .Y(n319) );
  MUX2X1 U624 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1200), .Y(n323) );
  MUX2X1 U625 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1200), .Y(n322) );
  MUX2X1 U626 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1200), .Y(n326) );
  MUX2X1 U627 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1200), .Y(n325) );
  MUX2X1 U628 ( .B(n324), .A(n321), .S(n1170), .Y(n335) );
  MUX2X1 U629 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1200), .Y(n329) );
  MUX2X1 U630 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1200), .Y(n328) );
  MUX2X1 U631 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1200), .Y(n332) );
  MUX2X1 U632 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1200), .Y(n331) );
  MUX2X1 U633 ( .B(n330), .A(n327), .S(n1170), .Y(n334) );
  MUX2X1 U634 ( .B(n333), .A(n318), .S(n1164), .Y(n641) );
  MUX2X1 U635 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1200), .Y(n338) );
  MUX2X1 U636 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1200), .Y(n337) );
  MUX2X1 U637 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1200), .Y(n341) );
  MUX2X1 U638 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1200), .Y(n340) );
  MUX2X1 U639 ( .B(n339), .A(n336), .S(n1169), .Y(n350) );
  MUX2X1 U640 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1201), .Y(n344) );
  MUX2X1 U641 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1201), .Y(n343) );
  MUX2X1 U642 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1201), .Y(n347) );
  MUX2X1 U643 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1201), .Y(n346) );
  MUX2X1 U644 ( .B(n345), .A(n342), .S(n1169), .Y(n349) );
  MUX2X1 U645 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1201), .Y(n353) );
  MUX2X1 U646 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1201), .Y(n352) );
  MUX2X1 U647 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1201), .Y(n356) );
  MUX2X1 U648 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1201), .Y(n355) );
  MUX2X1 U649 ( .B(n354), .A(n351), .S(n1169), .Y(n365) );
  MUX2X1 U650 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1201), .Y(n359) );
  MUX2X1 U651 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1201), .Y(n358) );
  MUX2X1 U652 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1201), .Y(n362) );
  MUX2X1 U653 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1201), .Y(n361) );
  MUX2X1 U654 ( .B(n360), .A(n357), .S(n1169), .Y(n364) );
  MUX2X1 U655 ( .B(n363), .A(n348), .S(n1164), .Y(n642) );
  MUX2X1 U656 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1202), .Y(n368) );
  MUX2X1 U657 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1202), .Y(n367) );
  MUX2X1 U658 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1202), .Y(n371) );
  MUX2X1 U659 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1202), .Y(n370) );
  MUX2X1 U660 ( .B(n369), .A(n366), .S(n1169), .Y(n380) );
  MUX2X1 U661 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1202), .Y(n374) );
  MUX2X1 U662 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1202), .Y(n373) );
  MUX2X1 U663 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1202), .Y(n377) );
  MUX2X1 U664 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1202), .Y(n376) );
  MUX2X1 U665 ( .B(n375), .A(n372), .S(n1169), .Y(n379) );
  MUX2X1 U666 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1202), .Y(n383) );
  MUX2X1 U667 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1202), .Y(n382) );
  MUX2X1 U668 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1202), .Y(n386) );
  MUX2X1 U669 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1202), .Y(n385) );
  MUX2X1 U670 ( .B(n384), .A(n381), .S(n1169), .Y(n395) );
  MUX2X1 U671 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1203), .Y(n389) );
  MUX2X1 U672 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1203), .Y(n388) );
  MUX2X1 U673 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1203), .Y(n392) );
  MUX2X1 U674 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1203), .Y(n391) );
  MUX2X1 U675 ( .B(n390), .A(n387), .S(n1169), .Y(n394) );
  MUX2X1 U676 ( .B(n393), .A(n378), .S(n1164), .Y(n643) );
  MUX2X1 U677 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1203), .Y(n398) );
  MUX2X1 U678 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1203), .Y(n397) );
  MUX2X1 U679 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1203), .Y(n401) );
  MUX2X1 U680 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1203), .Y(n400) );
  MUX2X1 U681 ( .B(n399), .A(n396), .S(n1169), .Y(n410) );
  MUX2X1 U682 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1203), .Y(n404) );
  MUX2X1 U683 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1203), .Y(n403) );
  MUX2X1 U684 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1203), .Y(n407) );
  MUX2X1 U685 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1203), .Y(n406) );
  MUX2X1 U686 ( .B(n405), .A(n402), .S(n1169), .Y(n409) );
  MUX2X1 U687 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1204), .Y(n413) );
  MUX2X1 U688 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1204), .Y(n412) );
  MUX2X1 U689 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1204), .Y(n416) );
  MUX2X1 U690 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1204), .Y(n415) );
  MUX2X1 U691 ( .B(n414), .A(n411), .S(n1169), .Y(n425) );
  MUX2X1 U692 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1204), .Y(n419) );
  MUX2X1 U693 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1204), .Y(n418) );
  MUX2X1 U694 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1204), .Y(n422) );
  MUX2X1 U695 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1204), .Y(n421) );
  MUX2X1 U696 ( .B(n420), .A(n417), .S(n1169), .Y(n424) );
  MUX2X1 U697 ( .B(n423), .A(n408), .S(n1164), .Y(n644) );
  MUX2X1 U698 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1204), .Y(n428) );
  MUX2X1 U699 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1204), .Y(n427) );
  MUX2X1 U700 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1204), .Y(n431) );
  MUX2X1 U701 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1204), .Y(n430) );
  MUX2X1 U702 ( .B(n429), .A(n426), .S(n1168), .Y(n440) );
  MUX2X1 U703 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1205), .Y(n434) );
  MUX2X1 U704 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1205), .Y(n433) );
  MUX2X1 U705 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1205), .Y(n437) );
  MUX2X1 U706 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1205), .Y(n436) );
  MUX2X1 U707 ( .B(n435), .A(n432), .S(n1168), .Y(n439) );
  MUX2X1 U708 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1205), .Y(n443) );
  MUX2X1 U709 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1205), .Y(n442) );
  MUX2X1 U710 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1205), .Y(n446) );
  MUX2X1 U711 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1205), .Y(n445) );
  MUX2X1 U712 ( .B(n444), .A(n441), .S(n1168), .Y(n455) );
  MUX2X1 U713 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1205), .Y(n449) );
  MUX2X1 U714 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1205), .Y(n448) );
  MUX2X1 U715 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1205), .Y(n452) );
  MUX2X1 U716 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1205), .Y(n451) );
  MUX2X1 U717 ( .B(n450), .A(n447), .S(n1168), .Y(n454) );
  MUX2X1 U718 ( .B(n453), .A(n438), .S(n1164), .Y(n645) );
  MUX2X1 U719 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1206), .Y(n458) );
  MUX2X1 U720 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1206), .Y(n457) );
  MUX2X1 U721 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1206), .Y(n461) );
  MUX2X1 U722 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1206), .Y(n460) );
  MUX2X1 U723 ( .B(n459), .A(n456), .S(n1168), .Y(n470) );
  MUX2X1 U724 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1206), .Y(n464) );
  MUX2X1 U725 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1206), .Y(n463) );
  MUX2X1 U726 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1206), .Y(n467) );
  MUX2X1 U727 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1206), .Y(n466) );
  MUX2X1 U728 ( .B(n465), .A(n462), .S(n1168), .Y(n469) );
  MUX2X1 U729 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1206), .Y(n473) );
  MUX2X1 U730 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1206), .Y(n472) );
  MUX2X1 U731 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1206), .Y(n476) );
  MUX2X1 U732 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1206), .Y(n475) );
  MUX2X1 U733 ( .B(n474), .A(n471), .S(n1168), .Y(n485) );
  MUX2X1 U734 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1207), .Y(n479) );
  MUX2X1 U735 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1207), .Y(n478) );
  MUX2X1 U736 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1207), .Y(n482) );
  MUX2X1 U737 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1207), .Y(n481) );
  MUX2X1 U738 ( .B(n480), .A(n477), .S(n1168), .Y(n484) );
  MUX2X1 U739 ( .B(n483), .A(n468), .S(n1164), .Y(n646) );
  MUX2X1 U740 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1207), .Y(n488) );
  MUX2X1 U741 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1207), .Y(n487) );
  MUX2X1 U742 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1207), .Y(n491) );
  MUX2X1 U743 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1207), .Y(n490) );
  MUX2X1 U744 ( .B(n489), .A(n486), .S(n1168), .Y(n500) );
  MUX2X1 U745 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1207), .Y(n494) );
  MUX2X1 U746 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1207), .Y(n493) );
  MUX2X1 U747 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1207), .Y(n497) );
  MUX2X1 U748 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1207), .Y(n496) );
  MUX2X1 U749 ( .B(n495), .A(n492), .S(n1168), .Y(n499) );
  MUX2X1 U750 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1208), .Y(n503) );
  MUX2X1 U751 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1208), .Y(n502) );
  MUX2X1 U752 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1208), .Y(n506) );
  MUX2X1 U753 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1208), .Y(n505) );
  MUX2X1 U754 ( .B(n504), .A(n501), .S(n1168), .Y(n515) );
  MUX2X1 U755 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1208), .Y(n509) );
  MUX2X1 U756 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1208), .Y(n508) );
  MUX2X1 U757 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1208), .Y(n512) );
  MUX2X1 U758 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1208), .Y(n511) );
  MUX2X1 U759 ( .B(n510), .A(n507), .S(n1168), .Y(n514) );
  MUX2X1 U760 ( .B(n513), .A(n498), .S(n1164), .Y(n647) );
  MUX2X1 U761 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1208), .Y(n518) );
  MUX2X1 U762 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1208), .Y(n517) );
  MUX2X1 U763 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1208), .Y(n521) );
  MUX2X1 U764 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1208), .Y(n520) );
  MUX2X1 U765 ( .B(n519), .A(n516), .S(n1167), .Y(n530) );
  MUX2X1 U766 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1209), .Y(n524) );
  MUX2X1 U767 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1209), .Y(n523) );
  MUX2X1 U768 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1209), .Y(n527) );
  MUX2X1 U769 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1209), .Y(n526) );
  MUX2X1 U770 ( .B(n525), .A(n522), .S(n1167), .Y(n529) );
  MUX2X1 U771 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1209), .Y(n533) );
  MUX2X1 U772 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1209), .Y(n532) );
  MUX2X1 U773 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1209), .Y(n536) );
  MUX2X1 U774 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1209), .Y(n535) );
  MUX2X1 U775 ( .B(n534), .A(n531), .S(n1167), .Y(n545) );
  MUX2X1 U776 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1209), .Y(n539) );
  MUX2X1 U777 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1209), .Y(n538) );
  MUX2X1 U778 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1209), .Y(n542) );
  MUX2X1 U779 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1209), .Y(n541) );
  MUX2X1 U780 ( .B(n540), .A(n537), .S(n1167), .Y(n544) );
  MUX2X1 U781 ( .B(n543), .A(n528), .S(n1164), .Y(n648) );
  MUX2X1 U782 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1210), .Y(n548) );
  MUX2X1 U783 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1210), .Y(n547) );
  MUX2X1 U784 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1210), .Y(n551) );
  MUX2X1 U785 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1210), .Y(n550) );
  MUX2X1 U786 ( .B(n549), .A(n546), .S(n1167), .Y(n560) );
  MUX2X1 U787 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1210), .Y(n554) );
  MUX2X1 U788 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1210), .Y(n553) );
  MUX2X1 U789 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1210), .Y(n557) );
  MUX2X1 U790 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1210), .Y(n556) );
  MUX2X1 U791 ( .B(n555), .A(n552), .S(n1167), .Y(n559) );
  MUX2X1 U792 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1210), .Y(n563) );
  MUX2X1 U793 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1210), .Y(n562) );
  MUX2X1 U794 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1210), .Y(n566) );
  MUX2X1 U795 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1210), .Y(n565) );
  MUX2X1 U796 ( .B(n564), .A(n561), .S(n1167), .Y(n575) );
  MUX2X1 U797 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1211), .Y(n569) );
  MUX2X1 U798 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1211), .Y(n568) );
  MUX2X1 U799 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1211), .Y(n572) );
  MUX2X1 U800 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1211), .Y(n571) );
  MUX2X1 U801 ( .B(n570), .A(n567), .S(n1167), .Y(n574) );
  MUX2X1 U802 ( .B(n573), .A(n558), .S(n1164), .Y(n649) );
  MUX2X1 U803 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1211), .Y(n578) );
  MUX2X1 U804 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1211), .Y(n577) );
  MUX2X1 U805 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1211), .Y(n581) );
  MUX2X1 U806 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1211), .Y(n580) );
  MUX2X1 U807 ( .B(n579), .A(n576), .S(n1167), .Y(n590) );
  MUX2X1 U808 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1211), .Y(n584) );
  MUX2X1 U809 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1211), .Y(n583) );
  MUX2X1 U810 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1211), .Y(n587) );
  MUX2X1 U811 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1211), .Y(n586) );
  MUX2X1 U812 ( .B(n585), .A(n582), .S(n1167), .Y(n589) );
  MUX2X1 U813 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1212), .Y(n593) );
  MUX2X1 U814 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1212), .Y(n592) );
  MUX2X1 U815 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1212), .Y(n596) );
  MUX2X1 U816 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1212), .Y(n595) );
  MUX2X1 U817 ( .B(n594), .A(n591), .S(n1167), .Y(n605) );
  MUX2X1 U818 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1212), .Y(n599) );
  MUX2X1 U819 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1212), .Y(n598) );
  MUX2X1 U820 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1212), .Y(n602) );
  MUX2X1 U821 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1212), .Y(n601) );
  MUX2X1 U822 ( .B(n600), .A(n597), .S(n1167), .Y(n604) );
  MUX2X1 U823 ( .B(n603), .A(n588), .S(n1164), .Y(n650) );
  MUX2X1 U824 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1212), .Y(n608) );
  MUX2X1 U825 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1212), .Y(n607) );
  MUX2X1 U826 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1212), .Y(n611) );
  MUX2X1 U827 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1212), .Y(n610) );
  MUX2X1 U828 ( .B(n609), .A(n606), .S(n1167), .Y(n620) );
  MUX2X1 U829 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1213), .Y(n614) );
  MUX2X1 U830 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1213), .Y(n613) );
  MUX2X1 U831 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1213), .Y(n617) );
  MUX2X1 U832 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1213), .Y(n616) );
  MUX2X1 U833 ( .B(n615), .A(n612), .S(n1168), .Y(n619) );
  MUX2X1 U834 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1213), .Y(n623) );
  MUX2X1 U835 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1213), .Y(n622) );
  MUX2X1 U836 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1213), .Y(n626) );
  MUX2X1 U837 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1213), .Y(n625) );
  MUX2X1 U838 ( .B(n624), .A(n621), .S(n1167), .Y(n635) );
  MUX2X1 U839 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1213), .Y(n629) );
  MUX2X1 U840 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1213), .Y(n628) );
  MUX2X1 U841 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1213), .Y(n632) );
  MUX2X1 U842 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1213), .Y(n631) );
  MUX2X1 U843 ( .B(n630), .A(n627), .S(n1168), .Y(n634) );
  MUX2X1 U844 ( .B(n633), .A(n618), .S(n1164), .Y(n1163) );
  INVX8 U845 ( .A(n1188), .Y(n1201) );
  INVX8 U846 ( .A(n1188), .Y(n1202) );
  INVX8 U847 ( .A(n1188), .Y(n1203) );
  INVX8 U848 ( .A(n1187), .Y(n1204) );
  INVX8 U849 ( .A(n1187), .Y(n1205) );
  INVX8 U850 ( .A(n1187), .Y(n1206) );
  INVX8 U851 ( .A(n1186), .Y(n1207) );
  INVX8 U852 ( .A(n1186), .Y(n1208) );
  INVX8 U853 ( .A(n1186), .Y(n1209) );
  INVX8 U854 ( .A(n1186), .Y(n1210) );
  INVX8 U855 ( .A(n1186), .Y(n1211) );
  INVX8 U856 ( .A(n1186), .Y(n1212) );
  INVX8 U857 ( .A(n1186), .Y(n1213) );
  INVX1 U858 ( .A(N11), .Y(n1375) );
  INVX1 U859 ( .A(N10), .Y(n1373) );
  INVX8 U860 ( .A(n1338), .Y(n1335) );
  INVX8 U861 ( .A(n1338), .Y(n1336) );
  INVX8 U862 ( .A(n1338), .Y(n1337) );
  INVX8 U863 ( .A(n4), .Y(n1339) );
  INVX8 U864 ( .A(n4), .Y(n1340) );
  INVX8 U865 ( .A(n7), .Y(n1341) );
  INVX8 U866 ( .A(n7), .Y(n1342) );
  INVX8 U867 ( .A(n8), .Y(n1343) );
  INVX8 U868 ( .A(n8), .Y(n1344) );
  INVX8 U869 ( .A(n9), .Y(n1345) );
  INVX8 U870 ( .A(n9), .Y(n1346) );
  INVX8 U871 ( .A(n10), .Y(n1347) );
  INVX8 U872 ( .A(n10), .Y(n1348) );
  INVX8 U873 ( .A(n11), .Y(n1349) );
  INVX8 U874 ( .A(n11), .Y(n1350) );
  INVX8 U875 ( .A(n12), .Y(n1351) );
  INVX8 U876 ( .A(n12), .Y(n1352) );
  INVX8 U877 ( .A(n13), .Y(n1353) );
  INVX8 U878 ( .A(n13), .Y(n1354) );
  INVX8 U879 ( .A(n14), .Y(n1355) );
  INVX8 U880 ( .A(n14), .Y(n1356) );
  INVX8 U881 ( .A(n15), .Y(n1357) );
  INVX8 U882 ( .A(n15), .Y(n1358) );
  INVX8 U883 ( .A(n16), .Y(n1359) );
  INVX8 U884 ( .A(n16), .Y(n1360) );
  INVX8 U885 ( .A(n17), .Y(n1361) );
  INVX8 U886 ( .A(n17), .Y(n1362) );
  INVX8 U887 ( .A(n18), .Y(n1363) );
  INVX8 U888 ( .A(n18), .Y(n1364) );
  INVX8 U889 ( .A(n19), .Y(n1365) );
  INVX8 U890 ( .A(n19), .Y(n1366) );
  INVX8 U891 ( .A(n20), .Y(n1367) );
  INVX8 U892 ( .A(n20), .Y(n1368) );
  INVX8 U893 ( .A(n21), .Y(n1369) );
  INVX8 U894 ( .A(n21), .Y(n1370) );
  AND2X2 U895 ( .A(n2), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U896 ( .A(n2), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U897 ( .A(n2), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U898 ( .A(n1), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U899 ( .A(n1), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U900 ( .A(n1), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U901 ( .A(n2), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U902 ( .A(n1), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U903 ( .A(n2), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U904 ( .A(n1), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U905 ( .A(n1), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U906 ( .A(n2), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U907 ( .A(n2), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U908 ( .A(n1), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U909 ( .A(n1), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U910 ( .A(n2), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U911 ( .A(\mem<31><0> ), .B(n1219), .Y(n1382) );
  OAI21X1 U912 ( .A(n1218), .B(n1339), .C(n1382), .Y(n2422) );
  NAND2X1 U913 ( .A(\mem<31><1> ), .B(n1219), .Y(n1383) );
  OAI21X1 U914 ( .A(n1342), .B(n1217), .C(n1383), .Y(n2421) );
  NAND2X1 U915 ( .A(\mem<31><2> ), .B(n1219), .Y(n1384) );
  OAI21X1 U916 ( .A(n1344), .B(n1217), .C(n1384), .Y(n2420) );
  NAND2X1 U917 ( .A(\mem<31><3> ), .B(n1219), .Y(n1385) );
  OAI21X1 U918 ( .A(n1346), .B(n1217), .C(n1385), .Y(n2419) );
  NAND2X1 U919 ( .A(\mem<31><4> ), .B(n1219), .Y(n1386) );
  OAI21X1 U920 ( .A(n1348), .B(n1217), .C(n1386), .Y(n2418) );
  NAND2X1 U921 ( .A(\mem<31><5> ), .B(n1219), .Y(n1387) );
  OAI21X1 U922 ( .A(n1350), .B(n1217), .C(n1387), .Y(n2417) );
  NAND2X1 U923 ( .A(\mem<31><6> ), .B(n1219), .Y(n1388) );
  OAI21X1 U924 ( .A(n1352), .B(n1217), .C(n1388), .Y(n2416) );
  NAND2X1 U925 ( .A(\mem<31><7> ), .B(n1219), .Y(n1389) );
  OAI21X1 U926 ( .A(n1354), .B(n1217), .C(n1389), .Y(n2415) );
  NAND2X1 U927 ( .A(\mem<31><8> ), .B(n1220), .Y(n1390) );
  OAI21X1 U928 ( .A(n1356), .B(n1217), .C(n1390), .Y(n2414) );
  NAND2X1 U929 ( .A(\mem<31><9> ), .B(n1220), .Y(n1391) );
  OAI21X1 U930 ( .A(n1358), .B(n1218), .C(n1391), .Y(n2413) );
  NAND2X1 U931 ( .A(\mem<31><10> ), .B(n1220), .Y(n1392) );
  OAI21X1 U932 ( .A(n1360), .B(n1218), .C(n1392), .Y(n2412) );
  NAND2X1 U933 ( .A(\mem<31><11> ), .B(n1220), .Y(n1393) );
  OAI21X1 U934 ( .A(n1362), .B(n1218), .C(n1393), .Y(n2411) );
  NAND2X1 U935 ( .A(\mem<31><12> ), .B(n1220), .Y(n1394) );
  OAI21X1 U936 ( .A(n1364), .B(n1218), .C(n1394), .Y(n2410) );
  NAND2X1 U937 ( .A(\mem<31><13> ), .B(n1220), .Y(n1395) );
  OAI21X1 U938 ( .A(n1366), .B(n1218), .C(n1395), .Y(n2409) );
  NAND2X1 U939 ( .A(\mem<31><14> ), .B(n1220), .Y(n1396) );
  OAI21X1 U940 ( .A(n1368), .B(n1218), .C(n1396), .Y(n2408) );
  NAND2X1 U941 ( .A(\mem<31><15> ), .B(n1220), .Y(n1397) );
  OAI21X1 U942 ( .A(n1370), .B(n1218), .C(n1397), .Y(n2407) );
  NAND2X1 U943 ( .A(\mem<30><0> ), .B(n1223), .Y(n1398) );
  OAI21X1 U944 ( .A(n1221), .B(n1339), .C(n1398), .Y(n2406) );
  NAND2X1 U945 ( .A(\mem<30><1> ), .B(n1223), .Y(n1399) );
  OAI21X1 U946 ( .A(n1221), .B(n1342), .C(n1399), .Y(n2405) );
  NAND2X1 U947 ( .A(\mem<30><2> ), .B(n1223), .Y(n1400) );
  OAI21X1 U948 ( .A(n1221), .B(n1344), .C(n1400), .Y(n2404) );
  NAND2X1 U949 ( .A(\mem<30><3> ), .B(n1223), .Y(n1401) );
  OAI21X1 U950 ( .A(n1221), .B(n1346), .C(n1401), .Y(n2403) );
  NAND2X1 U951 ( .A(\mem<30><4> ), .B(n1223), .Y(n1402) );
  OAI21X1 U952 ( .A(n1221), .B(n1348), .C(n1402), .Y(n2402) );
  NAND2X1 U953 ( .A(\mem<30><5> ), .B(n1223), .Y(n1403) );
  OAI21X1 U954 ( .A(n1221), .B(n1350), .C(n1403), .Y(n2401) );
  NAND2X1 U955 ( .A(\mem<30><6> ), .B(n1223), .Y(n1404) );
  OAI21X1 U956 ( .A(n1221), .B(n1352), .C(n1404), .Y(n2400) );
  NAND2X1 U957 ( .A(\mem<30><7> ), .B(n1223), .Y(n1405) );
  OAI21X1 U958 ( .A(n1221), .B(n1354), .C(n1405), .Y(n2399) );
  NAND2X1 U959 ( .A(\mem<30><8> ), .B(n1224), .Y(n1406) );
  OAI21X1 U960 ( .A(n1222), .B(n1355), .C(n1406), .Y(n2398) );
  NAND2X1 U961 ( .A(\mem<30><9> ), .B(n1224), .Y(n1407) );
  OAI21X1 U962 ( .A(n1222), .B(n1357), .C(n1407), .Y(n2397) );
  NAND2X1 U963 ( .A(\mem<30><10> ), .B(n1224), .Y(n1408) );
  OAI21X1 U964 ( .A(n1222), .B(n1359), .C(n1408), .Y(n2396) );
  NAND2X1 U965 ( .A(\mem<30><11> ), .B(n1224), .Y(n1409) );
  OAI21X1 U966 ( .A(n1222), .B(n1361), .C(n1409), .Y(n2395) );
  NAND2X1 U967 ( .A(\mem<30><12> ), .B(n1224), .Y(n1410) );
  OAI21X1 U968 ( .A(n1222), .B(n1363), .C(n1410), .Y(n2394) );
  NAND2X1 U969 ( .A(\mem<30><13> ), .B(n1224), .Y(n1411) );
  OAI21X1 U970 ( .A(n1222), .B(n1365), .C(n1411), .Y(n2393) );
  NAND2X1 U971 ( .A(\mem<30><14> ), .B(n1224), .Y(n1412) );
  OAI21X1 U972 ( .A(n1222), .B(n1367), .C(n1412), .Y(n2392) );
  NAND2X1 U973 ( .A(\mem<30><15> ), .B(n1224), .Y(n1413) );
  OAI21X1 U974 ( .A(n1222), .B(n1369), .C(n1413), .Y(n2391) );
  NAND3X1 U975 ( .A(n1372), .B(n1376), .C(n1375), .Y(n1414) );
  NAND2X1 U976 ( .A(\mem<29><0> ), .B(n1227), .Y(n1415) );
  OAI21X1 U977 ( .A(n1225), .B(n1339), .C(n1415), .Y(n2390) );
  NAND2X1 U978 ( .A(\mem<29><1> ), .B(n1227), .Y(n1416) );
  OAI21X1 U979 ( .A(n1225), .B(n1341), .C(n1416), .Y(n2389) );
  NAND2X1 U980 ( .A(\mem<29><2> ), .B(n1227), .Y(n1417) );
  OAI21X1 U981 ( .A(n1225), .B(n1343), .C(n1417), .Y(n2388) );
  NAND2X1 U982 ( .A(\mem<29><3> ), .B(n1227), .Y(n1418) );
  OAI21X1 U983 ( .A(n1225), .B(n1345), .C(n1418), .Y(n2387) );
  NAND2X1 U984 ( .A(\mem<29><4> ), .B(n1227), .Y(n1419) );
  OAI21X1 U985 ( .A(n1225), .B(n1347), .C(n1419), .Y(n2386) );
  NAND2X1 U986 ( .A(\mem<29><5> ), .B(n1227), .Y(n1420) );
  OAI21X1 U987 ( .A(n1225), .B(n1349), .C(n1420), .Y(n2385) );
  NAND2X1 U988 ( .A(\mem<29><6> ), .B(n1227), .Y(n1421) );
  OAI21X1 U989 ( .A(n1225), .B(n1351), .C(n1421), .Y(n2384) );
  NAND2X1 U990 ( .A(\mem<29><7> ), .B(n1227), .Y(n1422) );
  OAI21X1 U991 ( .A(n1225), .B(n1353), .C(n1422), .Y(n2383) );
  NAND2X1 U992 ( .A(\mem<29><8> ), .B(n1228), .Y(n1423) );
  OAI21X1 U993 ( .A(n1226), .B(n1356), .C(n1423), .Y(n2382) );
  NAND2X1 U994 ( .A(\mem<29><9> ), .B(n1228), .Y(n1424) );
  OAI21X1 U995 ( .A(n1226), .B(n1358), .C(n1424), .Y(n2381) );
  NAND2X1 U996 ( .A(\mem<29><10> ), .B(n1228), .Y(n1425) );
  OAI21X1 U997 ( .A(n1226), .B(n1360), .C(n1425), .Y(n2380) );
  NAND2X1 U998 ( .A(\mem<29><11> ), .B(n1228), .Y(n1426) );
  OAI21X1 U999 ( .A(n1226), .B(n1362), .C(n1426), .Y(n2379) );
  NAND2X1 U1000 ( .A(\mem<29><12> ), .B(n1228), .Y(n1427) );
  OAI21X1 U1001 ( .A(n1226), .B(n1364), .C(n1427), .Y(n2378) );
  NAND2X1 U1002 ( .A(\mem<29><13> ), .B(n1228), .Y(n1428) );
  OAI21X1 U1003 ( .A(n1226), .B(n1366), .C(n1428), .Y(n2377) );
  NAND2X1 U1004 ( .A(\mem<29><14> ), .B(n1228), .Y(n1429) );
  OAI21X1 U1005 ( .A(n1226), .B(n1368), .C(n1429), .Y(n2376) );
  NAND2X1 U1006 ( .A(\mem<29><15> ), .B(n1228), .Y(n1430) );
  OAI21X1 U1007 ( .A(n1226), .B(n1370), .C(n1430), .Y(n2375) );
  NAND3X1 U1008 ( .A(n1376), .B(n1375), .C(n1373), .Y(n1431) );
  NAND2X1 U1009 ( .A(\mem<28><0> ), .B(n1231), .Y(n1432) );
  OAI21X1 U1010 ( .A(n1229), .B(n1339), .C(n1432), .Y(n2374) );
  NAND2X1 U1011 ( .A(\mem<28><1> ), .B(n1231), .Y(n1433) );
  OAI21X1 U1012 ( .A(n1229), .B(n1342), .C(n1433), .Y(n2373) );
  NAND2X1 U1013 ( .A(\mem<28><2> ), .B(n1231), .Y(n1434) );
  OAI21X1 U1014 ( .A(n1229), .B(n1344), .C(n1434), .Y(n2372) );
  NAND2X1 U1015 ( .A(\mem<28><3> ), .B(n1231), .Y(n1435) );
  OAI21X1 U1016 ( .A(n1229), .B(n1346), .C(n1435), .Y(n2371) );
  NAND2X1 U1017 ( .A(\mem<28><4> ), .B(n1231), .Y(n1436) );
  OAI21X1 U1018 ( .A(n1229), .B(n1348), .C(n1436), .Y(n2370) );
  NAND2X1 U1019 ( .A(\mem<28><5> ), .B(n1231), .Y(n1437) );
  OAI21X1 U1020 ( .A(n1229), .B(n1350), .C(n1437), .Y(n2369) );
  NAND2X1 U1021 ( .A(\mem<28><6> ), .B(n1231), .Y(n1438) );
  OAI21X1 U1022 ( .A(n1229), .B(n1352), .C(n1438), .Y(n2368) );
  NAND2X1 U1023 ( .A(\mem<28><7> ), .B(n1231), .Y(n1439) );
  OAI21X1 U1024 ( .A(n1229), .B(n1354), .C(n1439), .Y(n2367) );
  NAND2X1 U1025 ( .A(\mem<28><8> ), .B(n1232), .Y(n1440) );
  OAI21X1 U1026 ( .A(n1230), .B(n1355), .C(n1440), .Y(n2366) );
  NAND2X1 U1027 ( .A(\mem<28><9> ), .B(n1232), .Y(n1441) );
  OAI21X1 U1028 ( .A(n1230), .B(n1357), .C(n1441), .Y(n2365) );
  NAND2X1 U1029 ( .A(\mem<28><10> ), .B(n1232), .Y(n1442) );
  OAI21X1 U1030 ( .A(n1230), .B(n1359), .C(n1442), .Y(n2364) );
  NAND2X1 U1031 ( .A(\mem<28><11> ), .B(n1232), .Y(n1443) );
  OAI21X1 U1032 ( .A(n1230), .B(n1361), .C(n1443), .Y(n2363) );
  NAND2X1 U1033 ( .A(\mem<28><12> ), .B(n1232), .Y(n1444) );
  OAI21X1 U1034 ( .A(n1230), .B(n1363), .C(n1444), .Y(n2362) );
  NAND2X1 U1035 ( .A(\mem<28><13> ), .B(n1232), .Y(n1445) );
  OAI21X1 U1036 ( .A(n1230), .B(n1365), .C(n1445), .Y(n2361) );
  NAND2X1 U1037 ( .A(\mem<28><14> ), .B(n1232), .Y(n1446) );
  OAI21X1 U1038 ( .A(n1230), .B(n1367), .C(n1446), .Y(n2360) );
  NAND2X1 U1039 ( .A(\mem<28><15> ), .B(n1232), .Y(n1447) );
  OAI21X1 U1040 ( .A(n1230), .B(n1369), .C(n1447), .Y(n2359) );
  NAND3X1 U1041 ( .A(n1372), .B(n1374), .C(n1377), .Y(n1448) );
  NAND2X1 U1042 ( .A(\mem<27><0> ), .B(n1235), .Y(n1449) );
  OAI21X1 U1043 ( .A(n1233), .B(n1339), .C(n1449), .Y(n2358) );
  NAND2X1 U1044 ( .A(\mem<27><1> ), .B(n1235), .Y(n1450) );
  OAI21X1 U1045 ( .A(n1233), .B(n1341), .C(n1450), .Y(n2357) );
  NAND2X1 U1046 ( .A(\mem<27><2> ), .B(n1235), .Y(n1451) );
  OAI21X1 U1047 ( .A(n1233), .B(n1343), .C(n1451), .Y(n2356) );
  NAND2X1 U1048 ( .A(\mem<27><3> ), .B(n1235), .Y(n1452) );
  OAI21X1 U1049 ( .A(n1233), .B(n1345), .C(n1452), .Y(n2355) );
  NAND2X1 U1050 ( .A(\mem<27><4> ), .B(n1235), .Y(n1453) );
  OAI21X1 U1051 ( .A(n1233), .B(n1347), .C(n1453), .Y(n2354) );
  NAND2X1 U1052 ( .A(\mem<27><5> ), .B(n1235), .Y(n1454) );
  OAI21X1 U1053 ( .A(n1233), .B(n1349), .C(n1454), .Y(n2353) );
  NAND2X1 U1054 ( .A(\mem<27><6> ), .B(n1235), .Y(n1455) );
  OAI21X1 U1055 ( .A(n1233), .B(n1351), .C(n1455), .Y(n2352) );
  NAND2X1 U1056 ( .A(\mem<27><7> ), .B(n1235), .Y(n1456) );
  OAI21X1 U1057 ( .A(n1233), .B(n1353), .C(n1456), .Y(n2351) );
  NAND2X1 U1058 ( .A(\mem<27><8> ), .B(n1236), .Y(n1457) );
  OAI21X1 U1059 ( .A(n1234), .B(n1356), .C(n1457), .Y(n2350) );
  NAND2X1 U1060 ( .A(\mem<27><9> ), .B(n1236), .Y(n1458) );
  OAI21X1 U1061 ( .A(n1234), .B(n1358), .C(n1458), .Y(n2349) );
  NAND2X1 U1062 ( .A(\mem<27><10> ), .B(n1236), .Y(n1459) );
  OAI21X1 U1063 ( .A(n1234), .B(n1360), .C(n1459), .Y(n2348) );
  NAND2X1 U1064 ( .A(\mem<27><11> ), .B(n1236), .Y(n1460) );
  OAI21X1 U1065 ( .A(n1234), .B(n1362), .C(n1460), .Y(n2347) );
  NAND2X1 U1066 ( .A(\mem<27><12> ), .B(n1236), .Y(n1461) );
  OAI21X1 U1067 ( .A(n1234), .B(n1364), .C(n1461), .Y(n2346) );
  NAND2X1 U1068 ( .A(\mem<27><13> ), .B(n1236), .Y(n1462) );
  OAI21X1 U1069 ( .A(n1234), .B(n1366), .C(n1462), .Y(n2345) );
  NAND2X1 U1070 ( .A(\mem<27><14> ), .B(n1236), .Y(n1463) );
  OAI21X1 U1071 ( .A(n1234), .B(n1368), .C(n1463), .Y(n2344) );
  NAND2X1 U1072 ( .A(\mem<27><15> ), .B(n1236), .Y(n1464) );
  OAI21X1 U1073 ( .A(n1234), .B(n1370), .C(n1464), .Y(n2343) );
  NAND3X1 U1074 ( .A(n1377), .B(n1374), .C(n1373), .Y(n1465) );
  NAND2X1 U1075 ( .A(\mem<26><0> ), .B(n1239), .Y(n1466) );
  OAI21X1 U1076 ( .A(n1237), .B(n1339), .C(n1466), .Y(n2342) );
  NAND2X1 U1077 ( .A(\mem<26><1> ), .B(n1239), .Y(n1467) );
  OAI21X1 U1078 ( .A(n1237), .B(n1342), .C(n1467), .Y(n2341) );
  NAND2X1 U1079 ( .A(\mem<26><2> ), .B(n1239), .Y(n1468) );
  OAI21X1 U1080 ( .A(n1237), .B(n1344), .C(n1468), .Y(n2340) );
  NAND2X1 U1081 ( .A(\mem<26><3> ), .B(n1239), .Y(n1469) );
  OAI21X1 U1082 ( .A(n1237), .B(n1346), .C(n1469), .Y(n2339) );
  NAND2X1 U1083 ( .A(\mem<26><4> ), .B(n1239), .Y(n1470) );
  OAI21X1 U1084 ( .A(n1237), .B(n1348), .C(n1470), .Y(n2338) );
  NAND2X1 U1085 ( .A(\mem<26><5> ), .B(n1239), .Y(n1471) );
  OAI21X1 U1086 ( .A(n1237), .B(n1350), .C(n1471), .Y(n2337) );
  NAND2X1 U1087 ( .A(\mem<26><6> ), .B(n1239), .Y(n1472) );
  OAI21X1 U1088 ( .A(n1237), .B(n1352), .C(n1472), .Y(n2336) );
  NAND2X1 U1089 ( .A(\mem<26><7> ), .B(n1239), .Y(n1473) );
  OAI21X1 U1090 ( .A(n1237), .B(n1354), .C(n1473), .Y(n2335) );
  NAND2X1 U1091 ( .A(\mem<26><8> ), .B(n1240), .Y(n1474) );
  OAI21X1 U1092 ( .A(n1238), .B(n1355), .C(n1474), .Y(n2334) );
  NAND2X1 U1093 ( .A(\mem<26><9> ), .B(n1240), .Y(n1475) );
  OAI21X1 U1094 ( .A(n1238), .B(n1357), .C(n1475), .Y(n2333) );
  NAND2X1 U1095 ( .A(\mem<26><10> ), .B(n1240), .Y(n1476) );
  OAI21X1 U1096 ( .A(n1238), .B(n1359), .C(n1476), .Y(n2332) );
  NAND2X1 U1097 ( .A(\mem<26><11> ), .B(n1240), .Y(n1477) );
  OAI21X1 U1098 ( .A(n1238), .B(n1361), .C(n1477), .Y(n2331) );
  NAND2X1 U1099 ( .A(\mem<26><12> ), .B(n1240), .Y(n1478) );
  OAI21X1 U1100 ( .A(n1238), .B(n1363), .C(n1478), .Y(n2330) );
  NAND2X1 U1101 ( .A(\mem<26><13> ), .B(n1240), .Y(n1479) );
  OAI21X1 U1102 ( .A(n1238), .B(n1365), .C(n1479), .Y(n2329) );
  NAND2X1 U1103 ( .A(\mem<26><14> ), .B(n1240), .Y(n1480) );
  OAI21X1 U1104 ( .A(n1238), .B(n1367), .C(n1480), .Y(n2328) );
  NAND2X1 U1105 ( .A(\mem<26><15> ), .B(n1240), .Y(n1481) );
  OAI21X1 U1106 ( .A(n1238), .B(n1369), .C(n1481), .Y(n2327) );
  NAND3X1 U1107 ( .A(n1372), .B(n1377), .C(n1375), .Y(n1482) );
  NAND2X1 U1108 ( .A(\mem<25><0> ), .B(n1243), .Y(n1483) );
  OAI21X1 U1109 ( .A(n1241), .B(n1339), .C(n1483), .Y(n2326) );
  NAND2X1 U1110 ( .A(\mem<25><1> ), .B(n1243), .Y(n1484) );
  OAI21X1 U1111 ( .A(n1241), .B(n1341), .C(n1484), .Y(n2325) );
  NAND2X1 U1112 ( .A(\mem<25><2> ), .B(n1243), .Y(n1485) );
  OAI21X1 U1113 ( .A(n1241), .B(n1343), .C(n1485), .Y(n2324) );
  NAND2X1 U1114 ( .A(\mem<25><3> ), .B(n1243), .Y(n1486) );
  OAI21X1 U1115 ( .A(n1241), .B(n1345), .C(n1486), .Y(n2323) );
  NAND2X1 U1116 ( .A(\mem<25><4> ), .B(n1243), .Y(n1487) );
  OAI21X1 U1117 ( .A(n1241), .B(n1347), .C(n1487), .Y(n2322) );
  NAND2X1 U1118 ( .A(\mem<25><5> ), .B(n1243), .Y(n1488) );
  OAI21X1 U1119 ( .A(n1241), .B(n1349), .C(n1488), .Y(n2321) );
  NAND2X1 U1120 ( .A(\mem<25><6> ), .B(n1243), .Y(n1489) );
  OAI21X1 U1121 ( .A(n1241), .B(n1351), .C(n1489), .Y(n2320) );
  NAND2X1 U1122 ( .A(\mem<25><7> ), .B(n1243), .Y(n1490) );
  OAI21X1 U1123 ( .A(n1241), .B(n1353), .C(n1490), .Y(n2319) );
  NAND2X1 U1124 ( .A(\mem<25><8> ), .B(n1244), .Y(n1491) );
  OAI21X1 U1125 ( .A(n1242), .B(n1356), .C(n1491), .Y(n2318) );
  NAND2X1 U1126 ( .A(\mem<25><9> ), .B(n1244), .Y(n1492) );
  OAI21X1 U1127 ( .A(n1242), .B(n1358), .C(n1492), .Y(n2317) );
  NAND2X1 U1128 ( .A(\mem<25><10> ), .B(n1244), .Y(n1493) );
  OAI21X1 U1129 ( .A(n1242), .B(n1360), .C(n1493), .Y(n2316) );
  NAND2X1 U1130 ( .A(\mem<25><11> ), .B(n1244), .Y(n1494) );
  OAI21X1 U1131 ( .A(n1242), .B(n1362), .C(n1494), .Y(n2315) );
  NAND2X1 U1132 ( .A(\mem<25><12> ), .B(n1244), .Y(n1495) );
  OAI21X1 U1133 ( .A(n1242), .B(n1364), .C(n1495), .Y(n2314) );
  NAND2X1 U1134 ( .A(\mem<25><13> ), .B(n1244), .Y(n1496) );
  OAI21X1 U1135 ( .A(n1242), .B(n1366), .C(n1496), .Y(n2313) );
  NAND2X1 U1136 ( .A(\mem<25><14> ), .B(n1244), .Y(n1497) );
  OAI21X1 U1137 ( .A(n1242), .B(n1368), .C(n1497), .Y(n2312) );
  NAND2X1 U1138 ( .A(\mem<25><15> ), .B(n1244), .Y(n1498) );
  OAI21X1 U1139 ( .A(n1242), .B(n1370), .C(n1498), .Y(n2311) );
  NOR3X1 U1140 ( .A(n1372), .B(n1374), .C(n1376), .Y(n1894) );
  NAND2X1 U1141 ( .A(\mem<24><0> ), .B(n1246), .Y(n1499) );
  OAI21X1 U1142 ( .A(n1245), .B(n1339), .C(n1499), .Y(n2310) );
  NAND2X1 U1143 ( .A(\mem<24><1> ), .B(n1246), .Y(n1500) );
  OAI21X1 U1144 ( .A(n1245), .B(n1341), .C(n1500), .Y(n2309) );
  NAND2X1 U1145 ( .A(\mem<24><2> ), .B(n1246), .Y(n1501) );
  OAI21X1 U1146 ( .A(n1245), .B(n1343), .C(n1501), .Y(n2308) );
  NAND2X1 U1147 ( .A(\mem<24><3> ), .B(n1246), .Y(n1502) );
  OAI21X1 U1148 ( .A(n1245), .B(n1345), .C(n1502), .Y(n2307) );
  NAND2X1 U1149 ( .A(\mem<24><4> ), .B(n1246), .Y(n1503) );
  OAI21X1 U1150 ( .A(n1245), .B(n1347), .C(n1503), .Y(n2306) );
  NAND2X1 U1151 ( .A(\mem<24><5> ), .B(n1246), .Y(n1504) );
  OAI21X1 U1152 ( .A(n1245), .B(n1349), .C(n1504), .Y(n2305) );
  NAND2X1 U1153 ( .A(\mem<24><6> ), .B(n1246), .Y(n1505) );
  OAI21X1 U1154 ( .A(n1245), .B(n1351), .C(n1505), .Y(n2304) );
  NAND2X1 U1155 ( .A(\mem<24><7> ), .B(n1246), .Y(n1506) );
  OAI21X1 U1156 ( .A(n1245), .B(n1353), .C(n1506), .Y(n2303) );
  NAND2X1 U1157 ( .A(\mem<24><8> ), .B(n1247), .Y(n1507) );
  OAI21X1 U1158 ( .A(n1245), .B(n1355), .C(n1507), .Y(n2302) );
  NAND2X1 U1159 ( .A(\mem<24><9> ), .B(n1247), .Y(n1508) );
  OAI21X1 U1160 ( .A(n1245), .B(n1357), .C(n1508), .Y(n2301) );
  NAND2X1 U1161 ( .A(\mem<24><10> ), .B(n1247), .Y(n1509) );
  OAI21X1 U1162 ( .A(n1245), .B(n1359), .C(n1509), .Y(n2300) );
  NAND2X1 U1163 ( .A(\mem<24><11> ), .B(n1247), .Y(n1510) );
  OAI21X1 U1164 ( .A(n1245), .B(n1361), .C(n1510), .Y(n2299) );
  NAND2X1 U1165 ( .A(\mem<24><12> ), .B(n1247), .Y(n1511) );
  OAI21X1 U1166 ( .A(n1245), .B(n1363), .C(n1511), .Y(n2298) );
  NAND2X1 U1167 ( .A(\mem<24><13> ), .B(n1247), .Y(n1512) );
  OAI21X1 U1168 ( .A(n1245), .B(n1365), .C(n1512), .Y(n2297) );
  NAND2X1 U1169 ( .A(\mem<24><14> ), .B(n1247), .Y(n1513) );
  OAI21X1 U1170 ( .A(n1245), .B(n1367), .C(n1513), .Y(n2296) );
  NAND2X1 U1171 ( .A(\mem<24><15> ), .B(n1247), .Y(n1514) );
  OAI21X1 U1172 ( .A(n1245), .B(n1369), .C(n1514), .Y(n2295) );
  NAND2X1 U1173 ( .A(\mem<23><0> ), .B(n1250), .Y(n1515) );
  OAI21X1 U1174 ( .A(n1248), .B(n1339), .C(n1515), .Y(n2294) );
  NAND2X1 U1175 ( .A(\mem<23><1> ), .B(n1250), .Y(n1516) );
  OAI21X1 U1177 ( .A(n1248), .B(n1342), .C(n1516), .Y(n2293) );
  NAND2X1 U1178 ( .A(\mem<23><2> ), .B(n1250), .Y(n1517) );
  OAI21X1 U1179 ( .A(n1248), .B(n1344), .C(n1517), .Y(n2292) );
  NAND2X1 U1180 ( .A(\mem<23><3> ), .B(n1250), .Y(n1518) );
  OAI21X1 U1181 ( .A(n1248), .B(n1346), .C(n1518), .Y(n2291) );
  NAND2X1 U1182 ( .A(\mem<23><4> ), .B(n1250), .Y(n1519) );
  OAI21X1 U1183 ( .A(n1248), .B(n1348), .C(n1519), .Y(n2290) );
  NAND2X1 U1184 ( .A(\mem<23><5> ), .B(n1250), .Y(n1520) );
  OAI21X1 U1185 ( .A(n1248), .B(n1350), .C(n1520), .Y(n2289) );
  NAND2X1 U1186 ( .A(\mem<23><6> ), .B(n1250), .Y(n1521) );
  OAI21X1 U1187 ( .A(n1248), .B(n1352), .C(n1521), .Y(n2288) );
  NAND2X1 U1188 ( .A(\mem<23><7> ), .B(n1250), .Y(n1522) );
  OAI21X1 U1189 ( .A(n1248), .B(n1354), .C(n1522), .Y(n2287) );
  NAND2X1 U1190 ( .A(\mem<23><8> ), .B(n1251), .Y(n1523) );
  OAI21X1 U1191 ( .A(n1249), .B(n1356), .C(n1523), .Y(n2286) );
  NAND2X1 U1192 ( .A(\mem<23><9> ), .B(n1251), .Y(n1524) );
  OAI21X1 U1193 ( .A(n1249), .B(n1358), .C(n1524), .Y(n2285) );
  NAND2X1 U1194 ( .A(\mem<23><10> ), .B(n1251), .Y(n1525) );
  OAI21X1 U1195 ( .A(n1249), .B(n1360), .C(n1525), .Y(n2284) );
  NAND2X1 U1196 ( .A(\mem<23><11> ), .B(n1251), .Y(n1526) );
  OAI21X1 U1197 ( .A(n1249), .B(n1362), .C(n1526), .Y(n2283) );
  NAND2X1 U1198 ( .A(\mem<23><12> ), .B(n1251), .Y(n1527) );
  OAI21X1 U1199 ( .A(n1249), .B(n1364), .C(n1527), .Y(n2282) );
  NAND2X1 U1200 ( .A(\mem<23><13> ), .B(n1251), .Y(n1528) );
  OAI21X1 U1201 ( .A(n1249), .B(n1366), .C(n1528), .Y(n2281) );
  NAND2X1 U1202 ( .A(\mem<23><14> ), .B(n1251), .Y(n1529) );
  OAI21X1 U1203 ( .A(n1249), .B(n1368), .C(n1529), .Y(n2280) );
  NAND2X1 U1204 ( .A(\mem<23><15> ), .B(n1251), .Y(n1530) );
  OAI21X1 U1205 ( .A(n1249), .B(n1370), .C(n1530), .Y(n2279) );
  NAND2X1 U1206 ( .A(\mem<22><0> ), .B(n1254), .Y(n1531) );
  OAI21X1 U1207 ( .A(n1252), .B(n1339), .C(n1531), .Y(n2278) );
  NAND2X1 U1208 ( .A(\mem<22><1> ), .B(n1254), .Y(n1532) );
  OAI21X1 U1209 ( .A(n1252), .B(n1342), .C(n1532), .Y(n2277) );
  NAND2X1 U1210 ( .A(\mem<22><2> ), .B(n1254), .Y(n1533) );
  OAI21X1 U1211 ( .A(n1252), .B(n1344), .C(n1533), .Y(n2276) );
  NAND2X1 U1212 ( .A(\mem<22><3> ), .B(n1254), .Y(n1534) );
  OAI21X1 U1213 ( .A(n1252), .B(n1346), .C(n1534), .Y(n2275) );
  NAND2X1 U1214 ( .A(\mem<22><4> ), .B(n1254), .Y(n1535) );
  OAI21X1 U1215 ( .A(n1252), .B(n1348), .C(n1535), .Y(n2274) );
  NAND2X1 U1216 ( .A(\mem<22><5> ), .B(n1254), .Y(n1536) );
  OAI21X1 U1217 ( .A(n1252), .B(n1350), .C(n1536), .Y(n2273) );
  NAND2X1 U1218 ( .A(\mem<22><6> ), .B(n1254), .Y(n1537) );
  OAI21X1 U1219 ( .A(n1252), .B(n1352), .C(n1537), .Y(n2272) );
  NAND2X1 U1220 ( .A(\mem<22><7> ), .B(n1254), .Y(n1538) );
  OAI21X1 U1221 ( .A(n1252), .B(n1354), .C(n1538), .Y(n2271) );
  NAND2X1 U1222 ( .A(\mem<22><8> ), .B(n1255), .Y(n1539) );
  OAI21X1 U1223 ( .A(n1253), .B(n1356), .C(n1539), .Y(n2270) );
  NAND2X1 U1224 ( .A(\mem<22><9> ), .B(n1255), .Y(n1540) );
  OAI21X1 U1225 ( .A(n1253), .B(n1358), .C(n1540), .Y(n2269) );
  NAND2X1 U1226 ( .A(\mem<22><10> ), .B(n1255), .Y(n1541) );
  OAI21X1 U1227 ( .A(n1253), .B(n1360), .C(n1541), .Y(n2268) );
  NAND2X1 U1228 ( .A(\mem<22><11> ), .B(n1255), .Y(n1542) );
  OAI21X1 U1229 ( .A(n1253), .B(n1362), .C(n1542), .Y(n2267) );
  NAND2X1 U1230 ( .A(\mem<22><12> ), .B(n1255), .Y(n1543) );
  OAI21X1 U1231 ( .A(n1253), .B(n1364), .C(n1543), .Y(n2266) );
  NAND2X1 U1232 ( .A(\mem<22><13> ), .B(n1255), .Y(n1544) );
  OAI21X1 U1233 ( .A(n1253), .B(n1366), .C(n1544), .Y(n2265) );
  NAND2X1 U1234 ( .A(\mem<22><14> ), .B(n1255), .Y(n1545) );
  OAI21X1 U1235 ( .A(n1253), .B(n1368), .C(n1545), .Y(n2264) );
  NAND2X1 U1236 ( .A(\mem<22><15> ), .B(n1255), .Y(n1546) );
  OAI21X1 U1237 ( .A(n1253), .B(n1370), .C(n1546), .Y(n2263) );
  NAND2X1 U1238 ( .A(\mem<21><0> ), .B(n1258), .Y(n1547) );
  OAI21X1 U1239 ( .A(n1256), .B(n1339), .C(n1547), .Y(n2262) );
  NAND2X1 U1240 ( .A(\mem<21><1> ), .B(n1258), .Y(n1548) );
  OAI21X1 U1241 ( .A(n1256), .B(n1342), .C(n1548), .Y(n2261) );
  NAND2X1 U1242 ( .A(\mem<21><2> ), .B(n1258), .Y(n1549) );
  OAI21X1 U1243 ( .A(n1256), .B(n1344), .C(n1549), .Y(n2260) );
  NAND2X1 U1244 ( .A(\mem<21><3> ), .B(n1258), .Y(n1550) );
  OAI21X1 U1245 ( .A(n1256), .B(n1346), .C(n1550), .Y(n2259) );
  NAND2X1 U1246 ( .A(\mem<21><4> ), .B(n1258), .Y(n1551) );
  OAI21X1 U1247 ( .A(n1256), .B(n1348), .C(n1551), .Y(n2258) );
  NAND2X1 U1248 ( .A(\mem<21><5> ), .B(n1258), .Y(n1552) );
  OAI21X1 U1249 ( .A(n1256), .B(n1350), .C(n1552), .Y(n2257) );
  NAND2X1 U1250 ( .A(\mem<21><6> ), .B(n1258), .Y(n1553) );
  OAI21X1 U1251 ( .A(n1256), .B(n1352), .C(n1553), .Y(n2256) );
  NAND2X1 U1252 ( .A(\mem<21><7> ), .B(n1258), .Y(n1554) );
  OAI21X1 U1253 ( .A(n1256), .B(n1354), .C(n1554), .Y(n2255) );
  NAND2X1 U1254 ( .A(\mem<21><8> ), .B(n1259), .Y(n1555) );
  OAI21X1 U1255 ( .A(n1257), .B(n1356), .C(n1555), .Y(n2254) );
  NAND2X1 U1256 ( .A(\mem<21><9> ), .B(n1259), .Y(n1556) );
  OAI21X1 U1257 ( .A(n1257), .B(n1358), .C(n1556), .Y(n2253) );
  NAND2X1 U1258 ( .A(\mem<21><10> ), .B(n1259), .Y(n1557) );
  OAI21X1 U1259 ( .A(n1257), .B(n1360), .C(n1557), .Y(n2252) );
  NAND2X1 U1260 ( .A(\mem<21><11> ), .B(n1259), .Y(n1558) );
  OAI21X1 U1261 ( .A(n1257), .B(n1362), .C(n1558), .Y(n2251) );
  NAND2X1 U1262 ( .A(\mem<21><12> ), .B(n1259), .Y(n1559) );
  OAI21X1 U1263 ( .A(n1257), .B(n1364), .C(n1559), .Y(n2250) );
  NAND2X1 U1264 ( .A(\mem<21><13> ), .B(n1259), .Y(n1560) );
  OAI21X1 U1265 ( .A(n1257), .B(n1366), .C(n1560), .Y(n2249) );
  NAND2X1 U1266 ( .A(\mem<21><14> ), .B(n1259), .Y(n1561) );
  OAI21X1 U1267 ( .A(n1257), .B(n1368), .C(n1561), .Y(n2248) );
  NAND2X1 U1268 ( .A(\mem<21><15> ), .B(n1259), .Y(n1562) );
  OAI21X1 U1269 ( .A(n1257), .B(n1370), .C(n1562), .Y(n2247) );
  NAND2X1 U1270 ( .A(\mem<20><0> ), .B(n1262), .Y(n1563) );
  OAI21X1 U1271 ( .A(n1260), .B(n1339), .C(n1563), .Y(n2246) );
  NAND2X1 U1272 ( .A(\mem<20><1> ), .B(n1262), .Y(n1564) );
  OAI21X1 U1273 ( .A(n1260), .B(n1342), .C(n1564), .Y(n2245) );
  NAND2X1 U1274 ( .A(\mem<20><2> ), .B(n1262), .Y(n1565) );
  OAI21X1 U1275 ( .A(n1260), .B(n1344), .C(n1565), .Y(n2244) );
  NAND2X1 U1276 ( .A(\mem<20><3> ), .B(n1262), .Y(n1566) );
  OAI21X1 U1277 ( .A(n1260), .B(n1346), .C(n1566), .Y(n2243) );
  NAND2X1 U1278 ( .A(\mem<20><4> ), .B(n1262), .Y(n1567) );
  OAI21X1 U1279 ( .A(n1260), .B(n1348), .C(n1567), .Y(n2242) );
  NAND2X1 U1280 ( .A(\mem<20><5> ), .B(n1262), .Y(n1568) );
  OAI21X1 U1281 ( .A(n1260), .B(n1350), .C(n1568), .Y(n2241) );
  NAND2X1 U1282 ( .A(\mem<20><6> ), .B(n1262), .Y(n1569) );
  OAI21X1 U1283 ( .A(n1260), .B(n1352), .C(n1569), .Y(n2240) );
  NAND2X1 U1284 ( .A(\mem<20><7> ), .B(n1262), .Y(n1570) );
  OAI21X1 U1285 ( .A(n1260), .B(n1354), .C(n1570), .Y(n2239) );
  NAND2X1 U1286 ( .A(\mem<20><8> ), .B(n1263), .Y(n1571) );
  OAI21X1 U1287 ( .A(n1261), .B(n1356), .C(n1571), .Y(n2238) );
  NAND2X1 U1288 ( .A(\mem<20><9> ), .B(n1263), .Y(n1572) );
  OAI21X1 U1289 ( .A(n1261), .B(n1358), .C(n1572), .Y(n2237) );
  NAND2X1 U1290 ( .A(\mem<20><10> ), .B(n1263), .Y(n1573) );
  OAI21X1 U1291 ( .A(n1261), .B(n1360), .C(n1573), .Y(n2236) );
  NAND2X1 U1292 ( .A(\mem<20><11> ), .B(n1263), .Y(n1574) );
  OAI21X1 U1293 ( .A(n1261), .B(n1362), .C(n1574), .Y(n2235) );
  NAND2X1 U1294 ( .A(\mem<20><12> ), .B(n1263), .Y(n1575) );
  OAI21X1 U1295 ( .A(n1261), .B(n1364), .C(n1575), .Y(n2234) );
  NAND2X1 U1296 ( .A(\mem<20><13> ), .B(n1263), .Y(n1576) );
  OAI21X1 U1297 ( .A(n1261), .B(n1366), .C(n1576), .Y(n2233) );
  NAND2X1 U1298 ( .A(\mem<20><14> ), .B(n1263), .Y(n1577) );
  OAI21X1 U1299 ( .A(n1261), .B(n1368), .C(n1577), .Y(n2232) );
  NAND2X1 U1300 ( .A(\mem<20><15> ), .B(n1263), .Y(n1578) );
  OAI21X1 U1301 ( .A(n1261), .B(n1370), .C(n1578), .Y(n2231) );
  NAND2X1 U1302 ( .A(\mem<19><0> ), .B(n1266), .Y(n1579) );
  OAI21X1 U1303 ( .A(n1264), .B(n1340), .C(n1579), .Y(n2230) );
  NAND2X1 U1304 ( .A(\mem<19><1> ), .B(n1266), .Y(n1580) );
  OAI21X1 U1305 ( .A(n1264), .B(n1342), .C(n1580), .Y(n2229) );
  NAND2X1 U1306 ( .A(\mem<19><2> ), .B(n1266), .Y(n1581) );
  OAI21X1 U1307 ( .A(n1264), .B(n1344), .C(n1581), .Y(n2228) );
  NAND2X1 U1308 ( .A(\mem<19><3> ), .B(n1266), .Y(n1582) );
  OAI21X1 U1309 ( .A(n1264), .B(n1346), .C(n1582), .Y(n2227) );
  NAND2X1 U1310 ( .A(\mem<19><4> ), .B(n1266), .Y(n1583) );
  OAI21X1 U1311 ( .A(n1264), .B(n1348), .C(n1583), .Y(n2226) );
  NAND2X1 U1312 ( .A(\mem<19><5> ), .B(n1266), .Y(n1584) );
  OAI21X1 U1313 ( .A(n1264), .B(n1350), .C(n1584), .Y(n2225) );
  NAND2X1 U1314 ( .A(\mem<19><6> ), .B(n1266), .Y(n1585) );
  OAI21X1 U1315 ( .A(n1264), .B(n1352), .C(n1585), .Y(n2224) );
  NAND2X1 U1316 ( .A(\mem<19><7> ), .B(n1266), .Y(n1586) );
  OAI21X1 U1317 ( .A(n1264), .B(n1354), .C(n1586), .Y(n2223) );
  NAND2X1 U1318 ( .A(\mem<19><8> ), .B(n1267), .Y(n1587) );
  OAI21X1 U1319 ( .A(n1265), .B(n1356), .C(n1587), .Y(n2222) );
  NAND2X1 U1320 ( .A(\mem<19><9> ), .B(n1267), .Y(n1588) );
  OAI21X1 U1321 ( .A(n1265), .B(n1358), .C(n1588), .Y(n2221) );
  NAND2X1 U1322 ( .A(\mem<19><10> ), .B(n1267), .Y(n1589) );
  OAI21X1 U1323 ( .A(n1265), .B(n1360), .C(n1589), .Y(n2220) );
  NAND2X1 U1324 ( .A(\mem<19><11> ), .B(n1267), .Y(n1590) );
  OAI21X1 U1325 ( .A(n1265), .B(n1362), .C(n1590), .Y(n2219) );
  NAND2X1 U1326 ( .A(\mem<19><12> ), .B(n1267), .Y(n1591) );
  OAI21X1 U1327 ( .A(n1265), .B(n1364), .C(n1591), .Y(n2218) );
  NAND2X1 U1328 ( .A(\mem<19><13> ), .B(n1267), .Y(n1592) );
  OAI21X1 U1329 ( .A(n1265), .B(n1366), .C(n1592), .Y(n2217) );
  NAND2X1 U1330 ( .A(\mem<19><14> ), .B(n1267), .Y(n1593) );
  OAI21X1 U1331 ( .A(n1265), .B(n1368), .C(n1593), .Y(n2216) );
  NAND2X1 U1332 ( .A(\mem<19><15> ), .B(n1267), .Y(n1594) );
  OAI21X1 U1333 ( .A(n1265), .B(n1370), .C(n1594), .Y(n2215) );
  NAND2X1 U1334 ( .A(\mem<18><0> ), .B(n1270), .Y(n1595) );
  OAI21X1 U1335 ( .A(n1268), .B(n1340), .C(n1595), .Y(n2214) );
  NAND2X1 U1336 ( .A(\mem<18><1> ), .B(n1270), .Y(n1596) );
  OAI21X1 U1337 ( .A(n1268), .B(n1342), .C(n1596), .Y(n2213) );
  NAND2X1 U1338 ( .A(\mem<18><2> ), .B(n1270), .Y(n1597) );
  OAI21X1 U1339 ( .A(n1268), .B(n1344), .C(n1597), .Y(n2212) );
  NAND2X1 U1340 ( .A(\mem<18><3> ), .B(n1270), .Y(n1598) );
  OAI21X1 U1341 ( .A(n1268), .B(n1346), .C(n1598), .Y(n2211) );
  NAND2X1 U1342 ( .A(\mem<18><4> ), .B(n1270), .Y(n1599) );
  OAI21X1 U1343 ( .A(n1268), .B(n1348), .C(n1599), .Y(n2210) );
  NAND2X1 U1344 ( .A(\mem<18><5> ), .B(n1270), .Y(n1600) );
  OAI21X1 U1345 ( .A(n1268), .B(n1350), .C(n1600), .Y(n2209) );
  NAND2X1 U1346 ( .A(\mem<18><6> ), .B(n1270), .Y(n1601) );
  OAI21X1 U1347 ( .A(n1268), .B(n1352), .C(n1601), .Y(n2208) );
  NAND2X1 U1348 ( .A(\mem<18><7> ), .B(n1270), .Y(n1602) );
  OAI21X1 U1349 ( .A(n1268), .B(n1354), .C(n1602), .Y(n2207) );
  NAND2X1 U1350 ( .A(\mem<18><8> ), .B(n1271), .Y(n1603) );
  OAI21X1 U1351 ( .A(n1269), .B(n1356), .C(n1603), .Y(n2206) );
  NAND2X1 U1352 ( .A(\mem<18><9> ), .B(n1271), .Y(n1604) );
  OAI21X1 U1353 ( .A(n1269), .B(n1358), .C(n1604), .Y(n2205) );
  NAND2X1 U1354 ( .A(\mem<18><10> ), .B(n1271), .Y(n1605) );
  OAI21X1 U1355 ( .A(n1269), .B(n1360), .C(n1605), .Y(n2204) );
  NAND2X1 U1356 ( .A(\mem<18><11> ), .B(n1271), .Y(n1606) );
  OAI21X1 U1357 ( .A(n1269), .B(n1362), .C(n1606), .Y(n2203) );
  NAND2X1 U1358 ( .A(\mem<18><12> ), .B(n1271), .Y(n1607) );
  OAI21X1 U1359 ( .A(n1269), .B(n1364), .C(n1607), .Y(n2202) );
  NAND2X1 U1360 ( .A(\mem<18><13> ), .B(n1271), .Y(n1608) );
  OAI21X1 U1361 ( .A(n1269), .B(n1366), .C(n1608), .Y(n2201) );
  NAND2X1 U1362 ( .A(\mem<18><14> ), .B(n1271), .Y(n1609) );
  OAI21X1 U1363 ( .A(n1269), .B(n1368), .C(n1609), .Y(n2200) );
  NAND2X1 U1364 ( .A(\mem<18><15> ), .B(n1271), .Y(n1610) );
  OAI21X1 U1365 ( .A(n1269), .B(n1370), .C(n1610), .Y(n2199) );
  NAND2X1 U1366 ( .A(\mem<17><0> ), .B(n1626), .Y(n1611) );
  OAI21X1 U1367 ( .A(n1272), .B(n1340), .C(n1611), .Y(n2198) );
  NAND2X1 U1368 ( .A(\mem<17><1> ), .B(n1626), .Y(n1612) );
  OAI21X1 U1369 ( .A(n1272), .B(n1342), .C(n1612), .Y(n2197) );
  NAND2X1 U1370 ( .A(\mem<17><2> ), .B(n1626), .Y(n1613) );
  OAI21X1 U1371 ( .A(n1272), .B(n1344), .C(n1613), .Y(n2196) );
  NAND2X1 U1372 ( .A(\mem<17><3> ), .B(n1626), .Y(n1614) );
  OAI21X1 U1373 ( .A(n1272), .B(n1346), .C(n1614), .Y(n2195) );
  NAND2X1 U1374 ( .A(\mem<17><4> ), .B(n1626), .Y(n1615) );
  OAI21X1 U1375 ( .A(n1272), .B(n1348), .C(n1615), .Y(n2194) );
  NAND2X1 U1376 ( .A(\mem<17><5> ), .B(n1626), .Y(n1616) );
  OAI21X1 U1377 ( .A(n1272), .B(n1350), .C(n1616), .Y(n2193) );
  NAND2X1 U1378 ( .A(\mem<17><6> ), .B(n1626), .Y(n1617) );
  OAI21X1 U1379 ( .A(n1272), .B(n1352), .C(n1617), .Y(n2192) );
  NAND2X1 U1380 ( .A(\mem<17><7> ), .B(n1626), .Y(n1618) );
  OAI21X1 U1381 ( .A(n1272), .B(n1354), .C(n1618), .Y(n2191) );
  NAND2X1 U1382 ( .A(\mem<17><8> ), .B(n1626), .Y(n1619) );
  OAI21X1 U1383 ( .A(n1273), .B(n1356), .C(n1619), .Y(n2190) );
  NAND2X1 U1384 ( .A(\mem<17><9> ), .B(n1626), .Y(n1620) );
  OAI21X1 U1385 ( .A(n1273), .B(n1358), .C(n1620), .Y(n2189) );
  NAND2X1 U1386 ( .A(\mem<17><10> ), .B(n1626), .Y(n1621) );
  OAI21X1 U1387 ( .A(n1273), .B(n1360), .C(n1621), .Y(n2188) );
  NAND2X1 U1388 ( .A(\mem<17><11> ), .B(n1626), .Y(n1622) );
  OAI21X1 U1389 ( .A(n1273), .B(n1362), .C(n1622), .Y(n2187) );
  NAND2X1 U1390 ( .A(\mem<17><12> ), .B(n1626), .Y(n1623) );
  OAI21X1 U1391 ( .A(n1273), .B(n1364), .C(n1623), .Y(n2186) );
  NAND2X1 U1392 ( .A(\mem<17><13> ), .B(n1626), .Y(n1624) );
  OAI21X1 U1393 ( .A(n1273), .B(n1366), .C(n1624), .Y(n2185) );
  NAND2X1 U1394 ( .A(\mem<17><14> ), .B(n1626), .Y(n1625) );
  OAI21X1 U1395 ( .A(n1273), .B(n1368), .C(n1625), .Y(n2184) );
  NAND2X1 U1396 ( .A(\mem<17><15> ), .B(n1626), .Y(n1627) );
  OAI21X1 U1397 ( .A(n1273), .B(n1370), .C(n1627), .Y(n2183) );
  NAND2X1 U1398 ( .A(\mem<16><0> ), .B(n1275), .Y(n1628) );
  OAI21X1 U1399 ( .A(n1274), .B(n1340), .C(n1628), .Y(n2182) );
  NAND2X1 U1400 ( .A(\mem<16><1> ), .B(n1275), .Y(n1629) );
  OAI21X1 U1401 ( .A(n1274), .B(n1342), .C(n1629), .Y(n2181) );
  NAND2X1 U1402 ( .A(\mem<16><2> ), .B(n1275), .Y(n1630) );
  OAI21X1 U1403 ( .A(n1274), .B(n1344), .C(n1630), .Y(n2180) );
  NAND2X1 U1404 ( .A(\mem<16><3> ), .B(n1275), .Y(n1631) );
  OAI21X1 U1405 ( .A(n1274), .B(n1346), .C(n1631), .Y(n2179) );
  NAND2X1 U1406 ( .A(\mem<16><4> ), .B(n1275), .Y(n1632) );
  OAI21X1 U1407 ( .A(n1274), .B(n1348), .C(n1632), .Y(n2178) );
  NAND2X1 U1408 ( .A(\mem<16><5> ), .B(n1275), .Y(n1633) );
  OAI21X1 U1409 ( .A(n1274), .B(n1350), .C(n1633), .Y(n2177) );
  NAND2X1 U1410 ( .A(\mem<16><6> ), .B(n1275), .Y(n1634) );
  OAI21X1 U1411 ( .A(n1274), .B(n1352), .C(n1634), .Y(n2176) );
  NAND2X1 U1412 ( .A(\mem<16><7> ), .B(n1275), .Y(n1635) );
  OAI21X1 U1413 ( .A(n1274), .B(n1354), .C(n1635), .Y(n2175) );
  NAND2X1 U1414 ( .A(\mem<16><8> ), .B(n1276), .Y(n1636) );
  OAI21X1 U1415 ( .A(n1274), .B(n1356), .C(n1636), .Y(n2174) );
  NAND2X1 U1416 ( .A(\mem<16><9> ), .B(n1276), .Y(n1637) );
  OAI21X1 U1417 ( .A(n1274), .B(n1358), .C(n1637), .Y(n2173) );
  NAND2X1 U1418 ( .A(\mem<16><10> ), .B(n1276), .Y(n1638) );
  OAI21X1 U1419 ( .A(n1274), .B(n1360), .C(n1638), .Y(n2172) );
  NAND2X1 U1420 ( .A(\mem<16><11> ), .B(n1276), .Y(n1639) );
  OAI21X1 U1421 ( .A(n1274), .B(n1362), .C(n1639), .Y(n2171) );
  NAND2X1 U1422 ( .A(\mem<16><12> ), .B(n1276), .Y(n1640) );
  OAI21X1 U1423 ( .A(n1274), .B(n1364), .C(n1640), .Y(n2170) );
  NAND2X1 U1424 ( .A(\mem<16><13> ), .B(n1276), .Y(n1641) );
  OAI21X1 U1425 ( .A(n1274), .B(n1366), .C(n1641), .Y(n2169) );
  NAND2X1 U1426 ( .A(\mem<16><14> ), .B(n1276), .Y(n1642) );
  OAI21X1 U1427 ( .A(n1274), .B(n1368), .C(n1642), .Y(n2168) );
  NAND2X1 U1428 ( .A(\mem<16><15> ), .B(n1276), .Y(n1643) );
  OAI21X1 U1429 ( .A(n1274), .B(n1370), .C(n1643), .Y(n2167) );
  NAND3X1 U1430 ( .A(n1378), .B(n2423), .C(n1381), .Y(n1644) );
  NAND2X1 U1431 ( .A(\mem<15><0> ), .B(n1279), .Y(n1645) );
  OAI21X1 U1432 ( .A(n1277), .B(n1340), .C(n1645), .Y(n2166) );
  NAND2X1 U1433 ( .A(\mem<15><1> ), .B(n1279), .Y(n1646) );
  OAI21X1 U1434 ( .A(n1277), .B(n1342), .C(n1646), .Y(n2165) );
  NAND2X1 U1435 ( .A(\mem<15><2> ), .B(n1279), .Y(n1647) );
  OAI21X1 U1436 ( .A(n1277), .B(n1344), .C(n1647), .Y(n2164) );
  NAND2X1 U1437 ( .A(\mem<15><3> ), .B(n1279), .Y(n1648) );
  OAI21X1 U1438 ( .A(n1277), .B(n1346), .C(n1648), .Y(n2163) );
  NAND2X1 U1439 ( .A(\mem<15><4> ), .B(n1279), .Y(n1649) );
  OAI21X1 U1440 ( .A(n1277), .B(n1348), .C(n1649), .Y(n2162) );
  NAND2X1 U1441 ( .A(\mem<15><5> ), .B(n1279), .Y(n1650) );
  OAI21X1 U1442 ( .A(n1277), .B(n1350), .C(n1650), .Y(n2161) );
  NAND2X1 U1443 ( .A(\mem<15><6> ), .B(n1279), .Y(n1651) );
  OAI21X1 U1444 ( .A(n1277), .B(n1352), .C(n1651), .Y(n2160) );
  NAND2X1 U1445 ( .A(\mem<15><7> ), .B(n1279), .Y(n1652) );
  OAI21X1 U1446 ( .A(n1277), .B(n1354), .C(n1652), .Y(n2159) );
  NAND2X1 U1447 ( .A(\mem<15><8> ), .B(n1280), .Y(n1653) );
  OAI21X1 U1448 ( .A(n1278), .B(n1356), .C(n1653), .Y(n2158) );
  NAND2X1 U1449 ( .A(\mem<15><9> ), .B(n1280), .Y(n1654) );
  OAI21X1 U1450 ( .A(n1278), .B(n1358), .C(n1654), .Y(n2157) );
  NAND2X1 U1451 ( .A(\mem<15><10> ), .B(n1280), .Y(n1655) );
  OAI21X1 U1452 ( .A(n1278), .B(n1360), .C(n1655), .Y(n2156) );
  NAND2X1 U1453 ( .A(\mem<15><11> ), .B(n1280), .Y(n1656) );
  OAI21X1 U1454 ( .A(n1278), .B(n1362), .C(n1656), .Y(n2155) );
  NAND2X1 U1455 ( .A(\mem<15><12> ), .B(n1280), .Y(n1657) );
  OAI21X1 U1456 ( .A(n1278), .B(n1364), .C(n1657), .Y(n2154) );
  NAND2X1 U1457 ( .A(\mem<15><13> ), .B(n1280), .Y(n1658) );
  OAI21X1 U1458 ( .A(n1278), .B(n1366), .C(n1658), .Y(n2153) );
  NAND2X1 U1459 ( .A(\mem<15><14> ), .B(n1280), .Y(n1659) );
  OAI21X1 U1460 ( .A(n1278), .B(n1368), .C(n1659), .Y(n2152) );
  NAND2X1 U1461 ( .A(\mem<15><15> ), .B(n1280), .Y(n1660) );
  OAI21X1 U1462 ( .A(n1278), .B(n1370), .C(n1660), .Y(n2151) );
  NAND2X1 U1463 ( .A(\mem<14><0> ), .B(n1283), .Y(n1661) );
  OAI21X1 U1464 ( .A(n1281), .B(n1340), .C(n1661), .Y(n2150) );
  NAND2X1 U1465 ( .A(\mem<14><1> ), .B(n1283), .Y(n1662) );
  OAI21X1 U1466 ( .A(n1281), .B(n1342), .C(n1662), .Y(n2149) );
  NAND2X1 U1467 ( .A(\mem<14><2> ), .B(n1283), .Y(n1663) );
  OAI21X1 U1468 ( .A(n1281), .B(n1344), .C(n1663), .Y(n2148) );
  NAND2X1 U1469 ( .A(\mem<14><3> ), .B(n1283), .Y(n1664) );
  OAI21X1 U1470 ( .A(n1281), .B(n1346), .C(n1664), .Y(n2147) );
  NAND2X1 U1471 ( .A(\mem<14><4> ), .B(n1283), .Y(n1665) );
  OAI21X1 U1472 ( .A(n1281), .B(n1348), .C(n1665), .Y(n2146) );
  NAND2X1 U1473 ( .A(\mem<14><5> ), .B(n1283), .Y(n1666) );
  OAI21X1 U1474 ( .A(n1281), .B(n1350), .C(n1666), .Y(n2145) );
  NAND2X1 U1475 ( .A(\mem<14><6> ), .B(n1283), .Y(n1667) );
  OAI21X1 U1476 ( .A(n1281), .B(n1352), .C(n1667), .Y(n2144) );
  NAND2X1 U1477 ( .A(\mem<14><7> ), .B(n1283), .Y(n1668) );
  OAI21X1 U1478 ( .A(n1281), .B(n1354), .C(n1668), .Y(n2143) );
  NAND2X1 U1479 ( .A(\mem<14><8> ), .B(n1284), .Y(n1669) );
  OAI21X1 U1480 ( .A(n1282), .B(n1356), .C(n1669), .Y(n2142) );
  NAND2X1 U1481 ( .A(\mem<14><9> ), .B(n1284), .Y(n1670) );
  OAI21X1 U1482 ( .A(n1282), .B(n1358), .C(n1670), .Y(n2141) );
  NAND2X1 U1483 ( .A(\mem<14><10> ), .B(n1284), .Y(n1671) );
  OAI21X1 U1484 ( .A(n1282), .B(n1360), .C(n1671), .Y(n2140) );
  NAND2X1 U1485 ( .A(\mem<14><11> ), .B(n1284), .Y(n1672) );
  OAI21X1 U1486 ( .A(n1282), .B(n1362), .C(n1672), .Y(n2139) );
  NAND2X1 U1487 ( .A(\mem<14><12> ), .B(n1284), .Y(n1673) );
  OAI21X1 U1488 ( .A(n1282), .B(n1364), .C(n1673), .Y(n2138) );
  NAND2X1 U1489 ( .A(\mem<14><13> ), .B(n1284), .Y(n1674) );
  OAI21X1 U1490 ( .A(n1282), .B(n1366), .C(n1674), .Y(n2137) );
  NAND2X1 U1491 ( .A(\mem<14><14> ), .B(n1284), .Y(n1675) );
  OAI21X1 U1492 ( .A(n1282), .B(n1368), .C(n1675), .Y(n2136) );
  NAND2X1 U1493 ( .A(\mem<14><15> ), .B(n1284), .Y(n1676) );
  OAI21X1 U1494 ( .A(n1282), .B(n1370), .C(n1676), .Y(n2135) );
  NAND2X1 U1495 ( .A(\mem<13><0> ), .B(n1287), .Y(n1677) );
  OAI21X1 U1496 ( .A(n1285), .B(n1340), .C(n1677), .Y(n2134) );
  NAND2X1 U1497 ( .A(\mem<13><1> ), .B(n1287), .Y(n1678) );
  OAI21X1 U1498 ( .A(n1285), .B(n1342), .C(n1678), .Y(n2133) );
  NAND2X1 U1499 ( .A(\mem<13><2> ), .B(n1287), .Y(n1679) );
  OAI21X1 U1500 ( .A(n1285), .B(n1344), .C(n1679), .Y(n2132) );
  NAND2X1 U1501 ( .A(\mem<13><3> ), .B(n1287), .Y(n1680) );
  OAI21X1 U1502 ( .A(n1285), .B(n1346), .C(n1680), .Y(n2131) );
  NAND2X1 U1503 ( .A(\mem<13><4> ), .B(n1287), .Y(n1681) );
  OAI21X1 U1504 ( .A(n1285), .B(n1348), .C(n1681), .Y(n2130) );
  NAND2X1 U1505 ( .A(\mem<13><5> ), .B(n1287), .Y(n1682) );
  OAI21X1 U1506 ( .A(n1285), .B(n1350), .C(n1682), .Y(n2129) );
  NAND2X1 U1507 ( .A(\mem<13><6> ), .B(n1287), .Y(n1683) );
  OAI21X1 U1508 ( .A(n1285), .B(n1352), .C(n1683), .Y(n2128) );
  NAND2X1 U1509 ( .A(\mem<13><7> ), .B(n1287), .Y(n1684) );
  OAI21X1 U1510 ( .A(n1285), .B(n1354), .C(n1684), .Y(n2127) );
  NAND2X1 U1511 ( .A(\mem<13><8> ), .B(n1288), .Y(n1685) );
  OAI21X1 U1512 ( .A(n1286), .B(n1356), .C(n1685), .Y(n2126) );
  NAND2X1 U1513 ( .A(\mem<13><9> ), .B(n1288), .Y(n1686) );
  OAI21X1 U1514 ( .A(n1286), .B(n1358), .C(n1686), .Y(n2125) );
  NAND2X1 U1515 ( .A(\mem<13><10> ), .B(n1288), .Y(n1687) );
  OAI21X1 U1516 ( .A(n1286), .B(n1360), .C(n1687), .Y(n2124) );
  NAND2X1 U1517 ( .A(\mem<13><11> ), .B(n1288), .Y(n1688) );
  OAI21X1 U1518 ( .A(n1286), .B(n1362), .C(n1688), .Y(n2123) );
  NAND2X1 U1519 ( .A(\mem<13><12> ), .B(n1288), .Y(n1689) );
  OAI21X1 U1520 ( .A(n1286), .B(n1364), .C(n1689), .Y(n2122) );
  NAND2X1 U1521 ( .A(\mem<13><13> ), .B(n1288), .Y(n1690) );
  OAI21X1 U1522 ( .A(n1286), .B(n1366), .C(n1690), .Y(n2121) );
  NAND2X1 U1523 ( .A(\mem<13><14> ), .B(n1288), .Y(n1691) );
  OAI21X1 U1524 ( .A(n1286), .B(n1368), .C(n1691), .Y(n2120) );
  NAND2X1 U1525 ( .A(\mem<13><15> ), .B(n1288), .Y(n1692) );
  OAI21X1 U1526 ( .A(n1286), .B(n1370), .C(n1692), .Y(n2119) );
  NAND2X1 U1527 ( .A(\mem<12><0> ), .B(n1708), .Y(n1693) );
  OAI21X1 U1528 ( .A(n1289), .B(n1340), .C(n1693), .Y(n2118) );
  NAND2X1 U1529 ( .A(\mem<12><1> ), .B(n1708), .Y(n1694) );
  OAI21X1 U1530 ( .A(n1289), .B(n1342), .C(n1694), .Y(n2117) );
  NAND2X1 U1531 ( .A(\mem<12><2> ), .B(n1708), .Y(n1695) );
  OAI21X1 U1532 ( .A(n1289), .B(n1344), .C(n1695), .Y(n2116) );
  NAND2X1 U1533 ( .A(\mem<12><3> ), .B(n1708), .Y(n1696) );
  OAI21X1 U1534 ( .A(n1289), .B(n1346), .C(n1696), .Y(n2115) );
  NAND2X1 U1535 ( .A(\mem<12><4> ), .B(n1708), .Y(n1697) );
  OAI21X1 U1536 ( .A(n1289), .B(n1348), .C(n1697), .Y(n2114) );
  NAND2X1 U1537 ( .A(\mem<12><5> ), .B(n1708), .Y(n1698) );
  OAI21X1 U1538 ( .A(n1289), .B(n1350), .C(n1698), .Y(n2113) );
  NAND2X1 U1539 ( .A(\mem<12><6> ), .B(n1708), .Y(n1699) );
  OAI21X1 U1540 ( .A(n1289), .B(n1352), .C(n1699), .Y(n2112) );
  NAND2X1 U1541 ( .A(\mem<12><7> ), .B(n1708), .Y(n1700) );
  OAI21X1 U1542 ( .A(n1289), .B(n1354), .C(n1700), .Y(n2111) );
  NAND2X1 U1543 ( .A(\mem<12><8> ), .B(n1708), .Y(n1701) );
  OAI21X1 U1544 ( .A(n1290), .B(n1356), .C(n1701), .Y(n2110) );
  NAND2X1 U1545 ( .A(\mem<12><9> ), .B(n1708), .Y(n1702) );
  OAI21X1 U1546 ( .A(n1290), .B(n1358), .C(n1702), .Y(n2109) );
  NAND2X1 U1547 ( .A(\mem<12><10> ), .B(n1708), .Y(n1703) );
  OAI21X1 U1548 ( .A(n1290), .B(n1360), .C(n1703), .Y(n2108) );
  NAND2X1 U1549 ( .A(\mem<12><11> ), .B(n1708), .Y(n1704) );
  OAI21X1 U1550 ( .A(n1290), .B(n1362), .C(n1704), .Y(n2107) );
  NAND2X1 U1551 ( .A(\mem<12><12> ), .B(n1708), .Y(n1705) );
  OAI21X1 U1552 ( .A(n1290), .B(n1364), .C(n1705), .Y(n2106) );
  NAND2X1 U1553 ( .A(\mem<12><13> ), .B(n1708), .Y(n1706) );
  OAI21X1 U1554 ( .A(n1290), .B(n1366), .C(n1706), .Y(n2105) );
  NAND2X1 U1555 ( .A(\mem<12><14> ), .B(n1708), .Y(n1707) );
  OAI21X1 U1556 ( .A(n1290), .B(n1368), .C(n1707), .Y(n2104) );
  NAND2X1 U1557 ( .A(\mem<12><15> ), .B(n1708), .Y(n1709) );
  OAI21X1 U1558 ( .A(n1290), .B(n1370), .C(n1709), .Y(n2103) );
  NAND2X1 U1559 ( .A(\mem<11><0> ), .B(n1293), .Y(n1710) );
  OAI21X1 U1560 ( .A(n1291), .B(n1340), .C(n1710), .Y(n2102) );
  NAND2X1 U1561 ( .A(\mem<11><1> ), .B(n1293), .Y(n1711) );
  OAI21X1 U1562 ( .A(n1291), .B(n1341), .C(n1711), .Y(n2101) );
  NAND2X1 U1563 ( .A(\mem<11><2> ), .B(n1293), .Y(n1712) );
  OAI21X1 U1564 ( .A(n1291), .B(n1343), .C(n1712), .Y(n2100) );
  NAND2X1 U1565 ( .A(\mem<11><3> ), .B(n1293), .Y(n1713) );
  OAI21X1 U1566 ( .A(n1291), .B(n1345), .C(n1713), .Y(n2099) );
  NAND2X1 U1567 ( .A(\mem<11><4> ), .B(n1293), .Y(n1714) );
  OAI21X1 U1568 ( .A(n1291), .B(n1347), .C(n1714), .Y(n2098) );
  NAND2X1 U1569 ( .A(\mem<11><5> ), .B(n1293), .Y(n1715) );
  OAI21X1 U1570 ( .A(n1291), .B(n1349), .C(n1715), .Y(n2097) );
  NAND2X1 U1571 ( .A(\mem<11><6> ), .B(n1293), .Y(n1716) );
  OAI21X1 U1572 ( .A(n1291), .B(n1351), .C(n1716), .Y(n2096) );
  NAND2X1 U1573 ( .A(\mem<11><7> ), .B(n1293), .Y(n1717) );
  OAI21X1 U1574 ( .A(n1291), .B(n1353), .C(n1717), .Y(n2095) );
  NAND2X1 U1575 ( .A(\mem<11><8> ), .B(n1294), .Y(n1718) );
  OAI21X1 U1576 ( .A(n1292), .B(n1355), .C(n1718), .Y(n2094) );
  NAND2X1 U1577 ( .A(\mem<11><9> ), .B(n1294), .Y(n1719) );
  OAI21X1 U1578 ( .A(n1292), .B(n1357), .C(n1719), .Y(n2093) );
  NAND2X1 U1579 ( .A(\mem<11><10> ), .B(n1294), .Y(n1720) );
  OAI21X1 U1580 ( .A(n1292), .B(n1359), .C(n1720), .Y(n2092) );
  NAND2X1 U1581 ( .A(\mem<11><11> ), .B(n1294), .Y(n1721) );
  OAI21X1 U1582 ( .A(n1292), .B(n1361), .C(n1721), .Y(n2091) );
  NAND2X1 U1583 ( .A(\mem<11><12> ), .B(n1294), .Y(n1722) );
  OAI21X1 U1584 ( .A(n1292), .B(n1363), .C(n1722), .Y(n2090) );
  NAND2X1 U1585 ( .A(\mem<11><13> ), .B(n1294), .Y(n1723) );
  OAI21X1 U1586 ( .A(n1292), .B(n1365), .C(n1723), .Y(n2089) );
  NAND2X1 U1587 ( .A(\mem<11><14> ), .B(n1294), .Y(n1724) );
  OAI21X1 U1588 ( .A(n1292), .B(n1367), .C(n1724), .Y(n2088) );
  NAND2X1 U1589 ( .A(\mem<11><15> ), .B(n1294), .Y(n1725) );
  OAI21X1 U1590 ( .A(n1292), .B(n1369), .C(n1725), .Y(n2087) );
  NAND2X1 U1591 ( .A(\mem<10><0> ), .B(n1297), .Y(n1726) );
  OAI21X1 U1592 ( .A(n1295), .B(n1340), .C(n1726), .Y(n2086) );
  NAND2X1 U1593 ( .A(\mem<10><1> ), .B(n1297), .Y(n1727) );
  OAI21X1 U1594 ( .A(n1295), .B(n1341), .C(n1727), .Y(n2085) );
  NAND2X1 U1595 ( .A(\mem<10><2> ), .B(n1297), .Y(n1728) );
  OAI21X1 U1596 ( .A(n1295), .B(n1343), .C(n1728), .Y(n2084) );
  NAND2X1 U1597 ( .A(\mem<10><3> ), .B(n1297), .Y(n1729) );
  OAI21X1 U1598 ( .A(n1295), .B(n1345), .C(n1729), .Y(n2083) );
  NAND2X1 U1599 ( .A(\mem<10><4> ), .B(n1297), .Y(n1730) );
  OAI21X1 U1600 ( .A(n1295), .B(n1347), .C(n1730), .Y(n2082) );
  NAND2X1 U1601 ( .A(\mem<10><5> ), .B(n1297), .Y(n1731) );
  OAI21X1 U1602 ( .A(n1295), .B(n1349), .C(n1731), .Y(n2081) );
  NAND2X1 U1603 ( .A(\mem<10><6> ), .B(n1297), .Y(n1732) );
  OAI21X1 U1604 ( .A(n1295), .B(n1351), .C(n1732), .Y(n2080) );
  NAND2X1 U1605 ( .A(\mem<10><7> ), .B(n1297), .Y(n1733) );
  OAI21X1 U1606 ( .A(n1295), .B(n1353), .C(n1733), .Y(n2079) );
  NAND2X1 U1607 ( .A(\mem<10><8> ), .B(n1298), .Y(n1734) );
  OAI21X1 U1608 ( .A(n1296), .B(n1355), .C(n1734), .Y(n2078) );
  NAND2X1 U1609 ( .A(\mem<10><9> ), .B(n1298), .Y(n1735) );
  OAI21X1 U1610 ( .A(n1296), .B(n1357), .C(n1735), .Y(n2077) );
  NAND2X1 U1611 ( .A(\mem<10><10> ), .B(n1298), .Y(n1736) );
  OAI21X1 U1612 ( .A(n1296), .B(n1359), .C(n1736), .Y(n2076) );
  NAND2X1 U1613 ( .A(\mem<10><11> ), .B(n1298), .Y(n1737) );
  OAI21X1 U1614 ( .A(n1296), .B(n1361), .C(n1737), .Y(n2075) );
  NAND2X1 U1615 ( .A(\mem<10><12> ), .B(n1298), .Y(n1738) );
  OAI21X1 U1616 ( .A(n1296), .B(n1363), .C(n1738), .Y(n2074) );
  NAND2X1 U1617 ( .A(\mem<10><13> ), .B(n1298), .Y(n1739) );
  OAI21X1 U1618 ( .A(n1296), .B(n1365), .C(n1739), .Y(n2073) );
  NAND2X1 U1619 ( .A(\mem<10><14> ), .B(n1298), .Y(n1740) );
  OAI21X1 U1620 ( .A(n1296), .B(n1367), .C(n1740), .Y(n2072) );
  NAND2X1 U1621 ( .A(\mem<10><15> ), .B(n1298), .Y(n1741) );
  OAI21X1 U1622 ( .A(n1296), .B(n1369), .C(n1741), .Y(n2071) );
  NAND2X1 U1623 ( .A(\mem<9><0> ), .B(n1301), .Y(n1742) );
  OAI21X1 U1624 ( .A(n1299), .B(n1340), .C(n1742), .Y(n2070) );
  NAND2X1 U1625 ( .A(\mem<9><1> ), .B(n1301), .Y(n1743) );
  OAI21X1 U1626 ( .A(n1299), .B(n1341), .C(n1743), .Y(n2069) );
  NAND2X1 U1627 ( .A(\mem<9><2> ), .B(n1301), .Y(n1744) );
  OAI21X1 U1628 ( .A(n1299), .B(n1343), .C(n1744), .Y(n2068) );
  NAND2X1 U1629 ( .A(\mem<9><3> ), .B(n1301), .Y(n1745) );
  OAI21X1 U1630 ( .A(n1299), .B(n1345), .C(n1745), .Y(n2067) );
  NAND2X1 U1631 ( .A(\mem<9><4> ), .B(n1301), .Y(n1746) );
  OAI21X1 U1632 ( .A(n1299), .B(n1347), .C(n1746), .Y(n2066) );
  NAND2X1 U1633 ( .A(\mem<9><5> ), .B(n1301), .Y(n1747) );
  OAI21X1 U1634 ( .A(n1299), .B(n1349), .C(n1747), .Y(n2065) );
  NAND2X1 U1635 ( .A(\mem<9><6> ), .B(n1301), .Y(n1748) );
  OAI21X1 U1636 ( .A(n1299), .B(n1351), .C(n1748), .Y(n2064) );
  NAND2X1 U1637 ( .A(\mem<9><7> ), .B(n1301), .Y(n1749) );
  OAI21X1 U1638 ( .A(n1299), .B(n1353), .C(n1749), .Y(n2063) );
  NAND2X1 U1639 ( .A(\mem<9><8> ), .B(n1302), .Y(n1750) );
  OAI21X1 U1640 ( .A(n1300), .B(n1355), .C(n1750), .Y(n2062) );
  NAND2X1 U1641 ( .A(\mem<9><9> ), .B(n1302), .Y(n1751) );
  OAI21X1 U1642 ( .A(n1300), .B(n1357), .C(n1751), .Y(n2061) );
  NAND2X1 U1643 ( .A(\mem<9><10> ), .B(n1302), .Y(n1752) );
  OAI21X1 U1644 ( .A(n1300), .B(n1359), .C(n1752), .Y(n2060) );
  NAND2X1 U1645 ( .A(\mem<9><11> ), .B(n1302), .Y(n1753) );
  OAI21X1 U1646 ( .A(n1300), .B(n1361), .C(n1753), .Y(n2059) );
  NAND2X1 U1647 ( .A(\mem<9><12> ), .B(n1302), .Y(n1754) );
  OAI21X1 U1648 ( .A(n1300), .B(n1363), .C(n1754), .Y(n2058) );
  NAND2X1 U1649 ( .A(\mem<9><13> ), .B(n1302), .Y(n1755) );
  OAI21X1 U1650 ( .A(n1300), .B(n1365), .C(n1755), .Y(n2057) );
  NAND2X1 U1651 ( .A(\mem<9><14> ), .B(n1302), .Y(n1756) );
  OAI21X1 U1652 ( .A(n1300), .B(n1367), .C(n1756), .Y(n2056) );
  NAND2X1 U1653 ( .A(\mem<9><15> ), .B(n1302), .Y(n1757) );
  OAI21X1 U1654 ( .A(n1300), .B(n1369), .C(n1757), .Y(n2055) );
  NAND2X1 U1655 ( .A(\mem<8><0> ), .B(n1304), .Y(n1759) );
  OAI21X1 U1656 ( .A(n1303), .B(n1340), .C(n1759), .Y(n2054) );
  NAND2X1 U1657 ( .A(\mem<8><1> ), .B(n1304), .Y(n1760) );
  OAI21X1 U1658 ( .A(n1303), .B(n1341), .C(n1760), .Y(n2053) );
  NAND2X1 U1659 ( .A(\mem<8><2> ), .B(n1304), .Y(n1761) );
  OAI21X1 U1660 ( .A(n1303), .B(n1343), .C(n1761), .Y(n2052) );
  NAND2X1 U1661 ( .A(\mem<8><3> ), .B(n1304), .Y(n1762) );
  OAI21X1 U1662 ( .A(n1303), .B(n1345), .C(n1762), .Y(n2051) );
  NAND2X1 U1663 ( .A(\mem<8><4> ), .B(n1304), .Y(n1763) );
  OAI21X1 U1664 ( .A(n1303), .B(n1347), .C(n1763), .Y(n2050) );
  NAND2X1 U1665 ( .A(\mem<8><5> ), .B(n1304), .Y(n1764) );
  OAI21X1 U1666 ( .A(n1303), .B(n1349), .C(n1764), .Y(n2049) );
  NAND2X1 U1667 ( .A(\mem<8><6> ), .B(n1304), .Y(n1765) );
  OAI21X1 U1668 ( .A(n1303), .B(n1351), .C(n1765), .Y(n2048) );
  NAND2X1 U1669 ( .A(\mem<8><7> ), .B(n1304), .Y(n1766) );
  OAI21X1 U1670 ( .A(n1303), .B(n1353), .C(n1766), .Y(n2047) );
  NAND2X1 U1671 ( .A(\mem<8><8> ), .B(n1305), .Y(n1767) );
  OAI21X1 U1672 ( .A(n1303), .B(n1355), .C(n1767), .Y(n2046) );
  NAND2X1 U1673 ( .A(\mem<8><9> ), .B(n1305), .Y(n1768) );
  OAI21X1 U1674 ( .A(n1303), .B(n1357), .C(n1768), .Y(n2045) );
  NAND2X1 U1675 ( .A(\mem<8><10> ), .B(n1305), .Y(n1769) );
  OAI21X1 U1676 ( .A(n1303), .B(n1359), .C(n1769), .Y(n2044) );
  NAND2X1 U1677 ( .A(\mem<8><11> ), .B(n1305), .Y(n1770) );
  OAI21X1 U1678 ( .A(n1303), .B(n1361), .C(n1770), .Y(n2043) );
  NAND2X1 U1679 ( .A(\mem<8><12> ), .B(n1305), .Y(n1771) );
  OAI21X1 U1680 ( .A(n1303), .B(n1363), .C(n1771), .Y(n2042) );
  NAND2X1 U1681 ( .A(\mem<8><13> ), .B(n1305), .Y(n1772) );
  OAI21X1 U1682 ( .A(n1303), .B(n1365), .C(n1772), .Y(n2041) );
  NAND2X1 U1683 ( .A(\mem<8><14> ), .B(n1305), .Y(n1773) );
  OAI21X1 U1684 ( .A(n1303), .B(n1367), .C(n1773), .Y(n2040) );
  NAND2X1 U1685 ( .A(\mem<8><15> ), .B(n1305), .Y(n1774) );
  OAI21X1 U1686 ( .A(n1303), .B(n1369), .C(n1774), .Y(n2039) );
  NAND3X1 U1687 ( .A(n1379), .B(n2423), .C(n1381), .Y(n1775) );
  NAND2X1 U1688 ( .A(\mem<7><0> ), .B(n1308), .Y(n1776) );
  OAI21X1 U1689 ( .A(n1306), .B(n1339), .C(n1776), .Y(n2038) );
  NAND2X1 U1690 ( .A(\mem<7><1> ), .B(n1308), .Y(n1777) );
  OAI21X1 U1691 ( .A(n1306), .B(n1341), .C(n1777), .Y(n2037) );
  NAND2X1 U1692 ( .A(\mem<7><2> ), .B(n1308), .Y(n1778) );
  OAI21X1 U1693 ( .A(n1306), .B(n1343), .C(n1778), .Y(n2036) );
  NAND2X1 U1694 ( .A(\mem<7><3> ), .B(n1308), .Y(n1779) );
  OAI21X1 U1695 ( .A(n1306), .B(n1345), .C(n1779), .Y(n2035) );
  NAND2X1 U1696 ( .A(\mem<7><4> ), .B(n1308), .Y(n1780) );
  OAI21X1 U1697 ( .A(n1306), .B(n1347), .C(n1780), .Y(n2034) );
  NAND2X1 U1698 ( .A(\mem<7><5> ), .B(n1308), .Y(n1781) );
  OAI21X1 U1699 ( .A(n1306), .B(n1349), .C(n1781), .Y(n2033) );
  NAND2X1 U1700 ( .A(\mem<7><6> ), .B(n1308), .Y(n1782) );
  OAI21X1 U1701 ( .A(n1306), .B(n1351), .C(n1782), .Y(n2032) );
  NAND2X1 U1702 ( .A(\mem<7><7> ), .B(n1308), .Y(n1783) );
  OAI21X1 U1703 ( .A(n1306), .B(n1353), .C(n1783), .Y(n2031) );
  NAND2X1 U1704 ( .A(\mem<7><8> ), .B(n1309), .Y(n1784) );
  OAI21X1 U1705 ( .A(n1307), .B(n1355), .C(n1784), .Y(n2030) );
  NAND2X1 U1706 ( .A(\mem<7><9> ), .B(n1309), .Y(n1785) );
  OAI21X1 U1707 ( .A(n1307), .B(n1357), .C(n1785), .Y(n2029) );
  NAND2X1 U1708 ( .A(\mem<7><10> ), .B(n1309), .Y(n1786) );
  OAI21X1 U1709 ( .A(n1307), .B(n1359), .C(n1786), .Y(n2028) );
  NAND2X1 U1710 ( .A(\mem<7><11> ), .B(n1309), .Y(n1787) );
  OAI21X1 U1711 ( .A(n1307), .B(n1361), .C(n1787), .Y(n2027) );
  NAND2X1 U1712 ( .A(\mem<7><12> ), .B(n1309), .Y(n1788) );
  OAI21X1 U1713 ( .A(n1307), .B(n1363), .C(n1788), .Y(n2026) );
  NAND2X1 U1714 ( .A(\mem<7><13> ), .B(n1309), .Y(n1789) );
  OAI21X1 U1715 ( .A(n1307), .B(n1365), .C(n1789), .Y(n2025) );
  NAND2X1 U1716 ( .A(\mem<7><14> ), .B(n1309), .Y(n1790) );
  OAI21X1 U1717 ( .A(n1307), .B(n1367), .C(n1790), .Y(n2024) );
  NAND2X1 U1718 ( .A(\mem<7><15> ), .B(n1309), .Y(n1791) );
  OAI21X1 U1719 ( .A(n1307), .B(n1369), .C(n1791), .Y(n2023) );
  NAND2X1 U1720 ( .A(\mem<6><0> ), .B(n1312), .Y(n1792) );
  OAI21X1 U1721 ( .A(n1310), .B(n1340), .C(n1792), .Y(n2022) );
  NAND2X1 U1722 ( .A(\mem<6><1> ), .B(n1312), .Y(n1793) );
  OAI21X1 U1723 ( .A(n1310), .B(n1341), .C(n1793), .Y(n2021) );
  NAND2X1 U1724 ( .A(\mem<6><2> ), .B(n1312), .Y(n1794) );
  OAI21X1 U1725 ( .A(n1310), .B(n1343), .C(n1794), .Y(n2020) );
  NAND2X1 U1726 ( .A(\mem<6><3> ), .B(n1312), .Y(n1795) );
  OAI21X1 U1727 ( .A(n1310), .B(n1345), .C(n1795), .Y(n2019) );
  NAND2X1 U1728 ( .A(\mem<6><4> ), .B(n1312), .Y(n1796) );
  OAI21X1 U1729 ( .A(n1310), .B(n1347), .C(n1796), .Y(n2018) );
  NAND2X1 U1730 ( .A(\mem<6><5> ), .B(n1312), .Y(n1797) );
  OAI21X1 U1731 ( .A(n1310), .B(n1349), .C(n1797), .Y(n2017) );
  NAND2X1 U1732 ( .A(\mem<6><6> ), .B(n1312), .Y(n1798) );
  OAI21X1 U1733 ( .A(n1310), .B(n1351), .C(n1798), .Y(n2016) );
  NAND2X1 U1734 ( .A(\mem<6><7> ), .B(n1312), .Y(n1799) );
  OAI21X1 U1735 ( .A(n1310), .B(n1353), .C(n1799), .Y(n2015) );
  NAND2X1 U1736 ( .A(\mem<6><8> ), .B(n1313), .Y(n1800) );
  OAI21X1 U1737 ( .A(n1311), .B(n1355), .C(n1800), .Y(n2014) );
  NAND2X1 U1738 ( .A(\mem<6><9> ), .B(n1313), .Y(n1801) );
  OAI21X1 U1739 ( .A(n1311), .B(n1357), .C(n1801), .Y(n2013) );
  NAND2X1 U1740 ( .A(\mem<6><10> ), .B(n1313), .Y(n1802) );
  OAI21X1 U1741 ( .A(n1311), .B(n1359), .C(n1802), .Y(n2012) );
  NAND2X1 U1742 ( .A(\mem<6><11> ), .B(n1313), .Y(n1803) );
  OAI21X1 U1743 ( .A(n1311), .B(n1361), .C(n1803), .Y(n2011) );
  NAND2X1 U1744 ( .A(\mem<6><12> ), .B(n1313), .Y(n1804) );
  OAI21X1 U1745 ( .A(n1311), .B(n1363), .C(n1804), .Y(n2010) );
  NAND2X1 U1746 ( .A(\mem<6><13> ), .B(n1313), .Y(n1805) );
  OAI21X1 U1747 ( .A(n1311), .B(n1365), .C(n1805), .Y(n2009) );
  NAND2X1 U1748 ( .A(\mem<6><14> ), .B(n1313), .Y(n1806) );
  OAI21X1 U1749 ( .A(n1311), .B(n1367), .C(n1806), .Y(n2008) );
  NAND2X1 U1750 ( .A(\mem<6><15> ), .B(n1313), .Y(n1807) );
  OAI21X1 U1751 ( .A(n1311), .B(n1369), .C(n1807), .Y(n2007) );
  NAND2X1 U1752 ( .A(\mem<5><0> ), .B(n1316), .Y(n1809) );
  OAI21X1 U1753 ( .A(n1314), .B(n1339), .C(n1809), .Y(n2006) );
  NAND2X1 U1754 ( .A(\mem<5><1> ), .B(n1316), .Y(n1810) );
  OAI21X1 U1755 ( .A(n1314), .B(n1341), .C(n1810), .Y(n2005) );
  NAND2X1 U1756 ( .A(\mem<5><2> ), .B(n1316), .Y(n1811) );
  OAI21X1 U1757 ( .A(n1314), .B(n1343), .C(n1811), .Y(n2004) );
  NAND2X1 U1758 ( .A(\mem<5><3> ), .B(n1316), .Y(n1812) );
  OAI21X1 U1759 ( .A(n1314), .B(n1345), .C(n1812), .Y(n2003) );
  NAND2X1 U1760 ( .A(\mem<5><4> ), .B(n1316), .Y(n1813) );
  OAI21X1 U1761 ( .A(n1314), .B(n1347), .C(n1813), .Y(n2002) );
  NAND2X1 U1762 ( .A(\mem<5><5> ), .B(n1316), .Y(n1814) );
  OAI21X1 U1763 ( .A(n1314), .B(n1349), .C(n1814), .Y(n2001) );
  NAND2X1 U1764 ( .A(\mem<5><6> ), .B(n1316), .Y(n1815) );
  OAI21X1 U1765 ( .A(n1314), .B(n1351), .C(n1815), .Y(n2000) );
  NAND2X1 U1766 ( .A(\mem<5><7> ), .B(n1316), .Y(n1816) );
  OAI21X1 U1767 ( .A(n1314), .B(n1353), .C(n1816), .Y(n1999) );
  NAND2X1 U1768 ( .A(\mem<5><8> ), .B(n1317), .Y(n1817) );
  OAI21X1 U1769 ( .A(n1315), .B(n1355), .C(n1817), .Y(n1998) );
  NAND2X1 U1770 ( .A(\mem<5><9> ), .B(n1317), .Y(n1818) );
  OAI21X1 U1771 ( .A(n1315), .B(n1357), .C(n1818), .Y(n1997) );
  NAND2X1 U1772 ( .A(\mem<5><10> ), .B(n1317), .Y(n1819) );
  OAI21X1 U1773 ( .A(n1315), .B(n1359), .C(n1819), .Y(n1996) );
  NAND2X1 U1774 ( .A(\mem<5><11> ), .B(n1317), .Y(n1820) );
  OAI21X1 U1775 ( .A(n1315), .B(n1361), .C(n1820), .Y(n1995) );
  NAND2X1 U1776 ( .A(\mem<5><12> ), .B(n1317), .Y(n1821) );
  OAI21X1 U1777 ( .A(n1315), .B(n1363), .C(n1821), .Y(n1994) );
  NAND2X1 U1778 ( .A(\mem<5><13> ), .B(n1317), .Y(n1822) );
  OAI21X1 U1779 ( .A(n1315), .B(n1365), .C(n1822), .Y(n1993) );
  NAND2X1 U1780 ( .A(\mem<5><14> ), .B(n1317), .Y(n1823) );
  OAI21X1 U1781 ( .A(n1315), .B(n1367), .C(n1823), .Y(n1992) );
  NAND2X1 U1782 ( .A(\mem<5><15> ), .B(n1317), .Y(n1824) );
  OAI21X1 U1783 ( .A(n1315), .B(n1369), .C(n1824), .Y(n1991) );
  NAND2X1 U1784 ( .A(\mem<4><0> ), .B(n92), .Y(n1826) );
  OAI21X1 U1785 ( .A(n1318), .B(n1340), .C(n1826), .Y(n1990) );
  NAND2X1 U1786 ( .A(\mem<4><1> ), .B(n92), .Y(n1827) );
  OAI21X1 U1787 ( .A(n1318), .B(n1341), .C(n1827), .Y(n1989) );
  NAND2X1 U1788 ( .A(\mem<4><2> ), .B(n92), .Y(n1828) );
  OAI21X1 U1789 ( .A(n1318), .B(n1343), .C(n1828), .Y(n1988) );
  NAND2X1 U1790 ( .A(\mem<4><3> ), .B(n92), .Y(n1829) );
  OAI21X1 U1791 ( .A(n1318), .B(n1345), .C(n1829), .Y(n1987) );
  NAND2X1 U1792 ( .A(\mem<4><4> ), .B(n92), .Y(n1830) );
  OAI21X1 U1793 ( .A(n1318), .B(n1347), .C(n1830), .Y(n1986) );
  NAND2X1 U1794 ( .A(\mem<4><5> ), .B(n92), .Y(n1831) );
  OAI21X1 U1795 ( .A(n1318), .B(n1349), .C(n1831), .Y(n1985) );
  NAND2X1 U1796 ( .A(\mem<4><6> ), .B(n92), .Y(n1832) );
  OAI21X1 U1797 ( .A(n1318), .B(n1351), .C(n1832), .Y(n1984) );
  NAND2X1 U1798 ( .A(\mem<4><7> ), .B(n92), .Y(n1833) );
  OAI21X1 U1799 ( .A(n1318), .B(n1353), .C(n1833), .Y(n1983) );
  NAND2X1 U1800 ( .A(\mem<4><8> ), .B(n92), .Y(n1834) );
  OAI21X1 U1801 ( .A(n1319), .B(n1355), .C(n1834), .Y(n1982) );
  NAND2X1 U1802 ( .A(\mem<4><9> ), .B(n92), .Y(n1835) );
  OAI21X1 U1803 ( .A(n1319), .B(n1357), .C(n1835), .Y(n1981) );
  NAND2X1 U1804 ( .A(\mem<4><10> ), .B(n92), .Y(n1836) );
  OAI21X1 U1805 ( .A(n1319), .B(n1359), .C(n1836), .Y(n1980) );
  NAND2X1 U1806 ( .A(\mem<4><11> ), .B(n92), .Y(n1837) );
  OAI21X1 U1807 ( .A(n1319), .B(n1361), .C(n1837), .Y(n1979) );
  NAND2X1 U1808 ( .A(\mem<4><12> ), .B(n92), .Y(n1838) );
  OAI21X1 U1809 ( .A(n1319), .B(n1363), .C(n1838), .Y(n1978) );
  NAND2X1 U1810 ( .A(\mem<4><13> ), .B(n92), .Y(n1839) );
  OAI21X1 U1811 ( .A(n1319), .B(n1365), .C(n1839), .Y(n1977) );
  NAND2X1 U1812 ( .A(\mem<4><14> ), .B(n92), .Y(n1840) );
  OAI21X1 U1813 ( .A(n1319), .B(n1367), .C(n1840), .Y(n1976) );
  NAND2X1 U1814 ( .A(\mem<4><15> ), .B(n92), .Y(n1841) );
  OAI21X1 U1815 ( .A(n1319), .B(n1369), .C(n1841), .Y(n1975) );
  NAND2X1 U1816 ( .A(\mem<3><0> ), .B(n1322), .Y(n1843) );
  OAI21X1 U1817 ( .A(n1320), .B(n1339), .C(n1843), .Y(n1974) );
  NAND2X1 U1818 ( .A(\mem<3><1> ), .B(n1322), .Y(n1844) );
  OAI21X1 U1819 ( .A(n1320), .B(n1341), .C(n1844), .Y(n1973) );
  NAND2X1 U1820 ( .A(\mem<3><2> ), .B(n1322), .Y(n1845) );
  OAI21X1 U1821 ( .A(n1320), .B(n1343), .C(n1845), .Y(n1972) );
  NAND2X1 U1822 ( .A(\mem<3><3> ), .B(n1322), .Y(n1846) );
  OAI21X1 U1823 ( .A(n1320), .B(n1345), .C(n1846), .Y(n1971) );
  NAND2X1 U1824 ( .A(\mem<3><4> ), .B(n1322), .Y(n1847) );
  OAI21X1 U1825 ( .A(n1320), .B(n1347), .C(n1847), .Y(n1970) );
  NAND2X1 U1826 ( .A(\mem<3><5> ), .B(n1322), .Y(n1848) );
  OAI21X1 U1827 ( .A(n1320), .B(n1349), .C(n1848), .Y(n1969) );
  NAND2X1 U1828 ( .A(\mem<3><6> ), .B(n1322), .Y(n1849) );
  OAI21X1 U1829 ( .A(n1320), .B(n1351), .C(n1849), .Y(n1968) );
  NAND2X1 U1830 ( .A(\mem<3><7> ), .B(n1322), .Y(n1850) );
  OAI21X1 U1831 ( .A(n1320), .B(n1353), .C(n1850), .Y(n1967) );
  NAND2X1 U1832 ( .A(\mem<3><8> ), .B(n1323), .Y(n1851) );
  OAI21X1 U1833 ( .A(n1321), .B(n1355), .C(n1851), .Y(n1966) );
  NAND2X1 U1834 ( .A(\mem<3><9> ), .B(n1323), .Y(n1852) );
  OAI21X1 U1835 ( .A(n1321), .B(n1357), .C(n1852), .Y(n1965) );
  NAND2X1 U1836 ( .A(\mem<3><10> ), .B(n1323), .Y(n1853) );
  OAI21X1 U1837 ( .A(n1321), .B(n1359), .C(n1853), .Y(n1964) );
  NAND2X1 U1838 ( .A(\mem<3><11> ), .B(n1323), .Y(n1854) );
  OAI21X1 U1839 ( .A(n1321), .B(n1361), .C(n1854), .Y(n1963) );
  NAND2X1 U1840 ( .A(\mem<3><12> ), .B(n1323), .Y(n1855) );
  OAI21X1 U1841 ( .A(n1321), .B(n1363), .C(n1855), .Y(n1962) );
  NAND2X1 U1842 ( .A(\mem<3><13> ), .B(n1323), .Y(n1856) );
  OAI21X1 U1843 ( .A(n1321), .B(n1365), .C(n1856), .Y(n1961) );
  NAND2X1 U1844 ( .A(\mem<3><14> ), .B(n1323), .Y(n1857) );
  OAI21X1 U1845 ( .A(n1321), .B(n1367), .C(n1857), .Y(n1960) );
  NAND2X1 U1846 ( .A(\mem<3><15> ), .B(n1323), .Y(n1858) );
  OAI21X1 U1847 ( .A(n1321), .B(n1369), .C(n1858), .Y(n1959) );
  NAND2X1 U1848 ( .A(\mem<2><0> ), .B(n1326), .Y(n1860) );
  OAI21X1 U1849 ( .A(n1324), .B(n1340), .C(n1860), .Y(n1958) );
  NAND2X1 U1850 ( .A(\mem<2><1> ), .B(n1326), .Y(n1861) );
  OAI21X1 U1851 ( .A(n1324), .B(n1341), .C(n1861), .Y(n1957) );
  NAND2X1 U1852 ( .A(\mem<2><2> ), .B(n1326), .Y(n1862) );
  OAI21X1 U1853 ( .A(n1324), .B(n1343), .C(n1862), .Y(n1956) );
  NAND2X1 U1854 ( .A(\mem<2><3> ), .B(n1326), .Y(n1863) );
  OAI21X1 U1855 ( .A(n1324), .B(n1345), .C(n1863), .Y(n1955) );
  NAND2X1 U1856 ( .A(\mem<2><4> ), .B(n1326), .Y(n1864) );
  OAI21X1 U1857 ( .A(n1324), .B(n1347), .C(n1864), .Y(n1954) );
  NAND2X1 U1858 ( .A(\mem<2><5> ), .B(n1326), .Y(n1865) );
  OAI21X1 U1859 ( .A(n1324), .B(n1349), .C(n1865), .Y(n1953) );
  NAND2X1 U1860 ( .A(\mem<2><6> ), .B(n1326), .Y(n1866) );
  OAI21X1 U1861 ( .A(n1324), .B(n1351), .C(n1866), .Y(n1952) );
  NAND2X1 U1862 ( .A(\mem<2><7> ), .B(n1326), .Y(n1867) );
  OAI21X1 U1863 ( .A(n1324), .B(n1353), .C(n1867), .Y(n1951) );
  NAND2X1 U1864 ( .A(\mem<2><8> ), .B(n1327), .Y(n1868) );
  OAI21X1 U1865 ( .A(n1325), .B(n1355), .C(n1868), .Y(n1950) );
  NAND2X1 U1866 ( .A(\mem<2><9> ), .B(n1327), .Y(n1869) );
  OAI21X1 U1867 ( .A(n1325), .B(n1357), .C(n1869), .Y(n1949) );
  NAND2X1 U1868 ( .A(\mem<2><10> ), .B(n1327), .Y(n1870) );
  OAI21X1 U1869 ( .A(n1325), .B(n1359), .C(n1870), .Y(n1948) );
  NAND2X1 U1870 ( .A(\mem<2><11> ), .B(n1327), .Y(n1871) );
  OAI21X1 U1871 ( .A(n1325), .B(n1361), .C(n1871), .Y(n1947) );
  NAND2X1 U1872 ( .A(\mem<2><12> ), .B(n1327), .Y(n1872) );
  OAI21X1 U1873 ( .A(n1325), .B(n1363), .C(n1872), .Y(n1946) );
  NAND2X1 U1874 ( .A(\mem<2><13> ), .B(n1327), .Y(n1873) );
  OAI21X1 U1875 ( .A(n1325), .B(n1365), .C(n1873), .Y(n1945) );
  NAND2X1 U1876 ( .A(\mem<2><14> ), .B(n1327), .Y(n1874) );
  OAI21X1 U1877 ( .A(n1325), .B(n1367), .C(n1874), .Y(n1944) );
  NAND2X1 U1878 ( .A(\mem<2><15> ), .B(n1327), .Y(n1875) );
  OAI21X1 U1879 ( .A(n1325), .B(n1369), .C(n1875), .Y(n1943) );
  NAND2X1 U1880 ( .A(\mem<1><0> ), .B(n1330), .Y(n1877) );
  OAI21X1 U1881 ( .A(n1328), .B(n1339), .C(n1877), .Y(n1942) );
  NAND2X1 U1882 ( .A(\mem<1><1> ), .B(n1330), .Y(n1878) );
  OAI21X1 U1883 ( .A(n1328), .B(n1341), .C(n1878), .Y(n1941) );
  NAND2X1 U1884 ( .A(\mem<1><2> ), .B(n1330), .Y(n1879) );
  OAI21X1 U1885 ( .A(n1328), .B(n1343), .C(n1879), .Y(n1940) );
  NAND2X1 U1886 ( .A(\mem<1><3> ), .B(n1330), .Y(n1880) );
  OAI21X1 U1887 ( .A(n1328), .B(n1345), .C(n1880), .Y(n1939) );
  NAND2X1 U1888 ( .A(\mem<1><4> ), .B(n1330), .Y(n1881) );
  OAI21X1 U1889 ( .A(n1328), .B(n1347), .C(n1881), .Y(n1938) );
  NAND2X1 U1890 ( .A(\mem<1><5> ), .B(n1330), .Y(n1882) );
  OAI21X1 U1891 ( .A(n1328), .B(n1349), .C(n1882), .Y(n1937) );
  NAND2X1 U1892 ( .A(\mem<1><6> ), .B(n1330), .Y(n1883) );
  OAI21X1 U1893 ( .A(n1328), .B(n1351), .C(n1883), .Y(n1936) );
  NAND2X1 U1894 ( .A(\mem<1><7> ), .B(n1330), .Y(n1884) );
  OAI21X1 U1895 ( .A(n1328), .B(n1353), .C(n1884), .Y(n1935) );
  NAND2X1 U1896 ( .A(\mem<1><8> ), .B(n1331), .Y(n1885) );
  OAI21X1 U1897 ( .A(n1329), .B(n1355), .C(n1885), .Y(n1934) );
  NAND2X1 U1898 ( .A(\mem<1><9> ), .B(n1331), .Y(n1886) );
  OAI21X1 U1899 ( .A(n1329), .B(n1357), .C(n1886), .Y(n1933) );
  NAND2X1 U1900 ( .A(\mem<1><10> ), .B(n1331), .Y(n1887) );
  OAI21X1 U1901 ( .A(n1329), .B(n1359), .C(n1887), .Y(n1932) );
  NAND2X1 U1902 ( .A(\mem<1><11> ), .B(n1331), .Y(n1888) );
  OAI21X1 U1903 ( .A(n1329), .B(n1361), .C(n1888), .Y(n1931) );
  NAND2X1 U1904 ( .A(\mem<1><12> ), .B(n1331), .Y(n1889) );
  OAI21X1 U1905 ( .A(n1329), .B(n1363), .C(n1889), .Y(n1930) );
  NAND2X1 U1906 ( .A(\mem<1><13> ), .B(n1331), .Y(n1890) );
  OAI21X1 U1907 ( .A(n1329), .B(n1365), .C(n1890), .Y(n1929) );
  NAND2X1 U1908 ( .A(\mem<1><14> ), .B(n1331), .Y(n1891) );
  OAI21X1 U1909 ( .A(n1329), .B(n1367), .C(n1891), .Y(n1928) );
  NAND2X1 U1910 ( .A(\mem<1><15> ), .B(n1331), .Y(n1892) );
  OAI21X1 U1911 ( .A(n1329), .B(n1369), .C(n1892), .Y(n1927) );
  NAND2X1 U1912 ( .A(\mem<0><0> ), .B(n1333), .Y(n1895) );
  OAI21X1 U1913 ( .A(n1332), .B(n1340), .C(n1895), .Y(n1926) );
  NAND2X1 U1914 ( .A(\mem<0><1> ), .B(n1333), .Y(n1896) );
  OAI21X1 U1915 ( .A(n1332), .B(n1341), .C(n1896), .Y(n1925) );
  NAND2X1 U1916 ( .A(\mem<0><2> ), .B(n1333), .Y(n1897) );
  OAI21X1 U1917 ( .A(n1332), .B(n1343), .C(n1897), .Y(n1924) );
  NAND2X1 U1918 ( .A(\mem<0><3> ), .B(n1333), .Y(n1898) );
  OAI21X1 U1919 ( .A(n1332), .B(n1345), .C(n1898), .Y(n1923) );
  NAND2X1 U1920 ( .A(\mem<0><4> ), .B(n1333), .Y(n1899) );
  OAI21X1 U1921 ( .A(n1332), .B(n1347), .C(n1899), .Y(n1922) );
  NAND2X1 U1922 ( .A(\mem<0><5> ), .B(n1333), .Y(n1900) );
  OAI21X1 U1923 ( .A(n1332), .B(n1349), .C(n1900), .Y(n1921) );
  NAND2X1 U1924 ( .A(\mem<0><6> ), .B(n1333), .Y(n1901) );
  OAI21X1 U1925 ( .A(n1332), .B(n1351), .C(n1901), .Y(n1920) );
  NAND2X1 U1926 ( .A(\mem<0><7> ), .B(n1333), .Y(n1902) );
  OAI21X1 U1927 ( .A(n1332), .B(n1353), .C(n1902), .Y(n1919) );
  NAND2X1 U1928 ( .A(\mem<0><8> ), .B(n1334), .Y(n1903) );
  OAI21X1 U1929 ( .A(n1332), .B(n1355), .C(n1903), .Y(n1918) );
  NAND2X1 U1930 ( .A(\mem<0><9> ), .B(n1334), .Y(n1904) );
  OAI21X1 U1931 ( .A(n1332), .B(n1357), .C(n1904), .Y(n1917) );
  NAND2X1 U1932 ( .A(\mem<0><10> ), .B(n1334), .Y(n1905) );
  OAI21X1 U1933 ( .A(n1332), .B(n1359), .C(n1905), .Y(n1916) );
  NAND2X1 U1934 ( .A(\mem<0><11> ), .B(n1334), .Y(n1906) );
  OAI21X1 U1935 ( .A(n1332), .B(n1361), .C(n1906), .Y(n1915) );
  NAND2X1 U1936 ( .A(\mem<0><12> ), .B(n1334), .Y(n1907) );
  OAI21X1 U1937 ( .A(n1332), .B(n1363), .C(n1907), .Y(n1914) );
  NAND2X1 U1938 ( .A(\mem<0><13> ), .B(n1334), .Y(n1908) );
  OAI21X1 U1939 ( .A(n1332), .B(n1365), .C(n1908), .Y(n1913) );
  NAND2X1 U1940 ( .A(\mem<0><14> ), .B(n1334), .Y(n1909) );
  OAI21X1 U1941 ( .A(n1332), .B(n1367), .C(n1909), .Y(n1912) );
  NAND2X1 U1942 ( .A(\mem<0><15> ), .B(n1334), .Y(n1910) );
  OAI21X1 U1943 ( .A(n1332), .B(n1369), .C(n1910), .Y(n1911) );
endmodule


module memc_Size5_1 ( .data_out({\data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        write, clk, rst, createdump, .file_id({\file_id<4> , \file_id<3> , 
        \file_id<2> , \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<4> , \data_in<3> , \data_in<2> ,
         \data_in<1> , \data_in<0> , write, clk, rst, createdump, \file_id<4> ,
         \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> ,
         \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><4> , \mem<0><3> , \mem<0><2> ,
         \mem<0><1> , \mem<0><0> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><4> , \mem<3><3> , \mem<3><2> ,
         \mem<3><1> , \mem<3><0> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><4> , \mem<5><3> , \mem<5><2> ,
         \mem<5><1> , \mem<5><0> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><4> , \mem<8><3> , \mem<8><2> ,
         \mem<8><1> , \mem<8><0> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><4> , \mem<10><3> , \mem<10><2> ,
         \mem<10><1> , \mem<10><0> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><4> , \mem<13><3> , \mem<13><2> ,
         \mem<13><1> , \mem<13><0> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><4> , \mem<15><3> , \mem<15><2> ,
         \mem<15><1> , \mem<15><0> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><4> , \mem<18><3> , \mem<18><2> ,
         \mem<18><1> , \mem<18><0> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><4> , \mem<20><3> , \mem<20><2> ,
         \mem<20><1> , \mem<20><0> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><4> , \mem<23><3> , \mem<23><2> ,
         \mem<23><1> , \mem<23><0> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><4> , \mem<25><3> , \mem<25><2> ,
         \mem<25><1> , \mem<25><0> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><4> , \mem<28><3> , \mem<28><2> ,
         \mem<28><1> , \mem<28><0> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><4> , \mem<30><3> , \mem<30><2> ,
         \mem<30><1> , \mem<30><0> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , N17, N18, N19, N20, N21, n56, n57, n65,
         n73, n81, n89, n97, n105, n113, n114, n115, n172, n229, n286, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n58, n59, n60, n61, n62, n63, n64, n66, n67, n68, n69,
         n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85,
         n86, n87, n88, n90, n91, n92, n93, n94, n95, n96, n98, n99, n100,
         n101, n102, n103, n104, n106, n107, n108, n109, n110, n111, n112,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n287, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><4>  ( .D(n447), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n446), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n445), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n444), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n443), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n442), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n441), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n440), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n439), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n438), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n437), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n436), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n435), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n434), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n433), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n432), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n431), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n430), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n429), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n428), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n427), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n426), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n425), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n424), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n423), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n422), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n421), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n420), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n419), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n418), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n417), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n416), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n415), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n414), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n413), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n412), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n411), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n410), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n409), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n408), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n407), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n406), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n405), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n404), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n403), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n402), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n401), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n400), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n399), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n398), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n397), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n396), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n395), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n394), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n393), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n392), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n391), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n390), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n389), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n388), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n387), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n386), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n385), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n384), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n383), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n382), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n381), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n380), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n379), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n378), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n377), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n376), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n375), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n374), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n373), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n372), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n371), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n370), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n369), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n368), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n367), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n366), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n365), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n364), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n363), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n362), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n361), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n360), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n359), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n358), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n357), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n356), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n355), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n354), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n353), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n352), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n351), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n350), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n349), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n348), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n347), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n346), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n345), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n344), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n343), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n342), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n341), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n340), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n339), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n338), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n337), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n336), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n335), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n334), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n333), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n332), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n331), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n330), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n329), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n328), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n327), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n326), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n325), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n324), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n323), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n322), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n321), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n320), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n319), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n318), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n317), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n316), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n315), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n314), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n313), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n312), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n311), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n310), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n309), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n308), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n307), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n306), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n305), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n304), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n303), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n302), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n301), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n300), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n299), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n298), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n297), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n296), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n295), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n294), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n292), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n291), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n290), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n289), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n288), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(n648), .B(n824), .Y(n56) );
  OAI21X1 U50 ( .A(n579), .B(n823), .C(n497), .Y(n288) );
  OAI21X1 U52 ( .A(n579), .B(n822), .C(n495), .Y(n289) );
  OAI21X1 U54 ( .A(n579), .B(n821), .C(n493), .Y(n290) );
  OAI21X1 U56 ( .A(n579), .B(n820), .C(n491), .Y(n291) );
  OAI21X1 U58 ( .A(n579), .B(n819), .C(n489), .Y(n292) );
  OAI21X1 U62 ( .A(n823), .B(n642), .C(n487), .Y(n293) );
  OAI21X1 U64 ( .A(n822), .B(n642), .C(n485), .Y(n294) );
  OAI21X1 U66 ( .A(n821), .B(n642), .C(n483), .Y(n295) );
  OAI21X1 U68 ( .A(n820), .B(n642), .C(n481), .Y(n296) );
  OAI21X1 U70 ( .A(n819), .B(n642), .C(n479), .Y(n297) );
  OAI21X1 U74 ( .A(n823), .B(n640), .C(n477), .Y(n298) );
  OAI21X1 U76 ( .A(n822), .B(n640), .C(n475), .Y(n299) );
  OAI21X1 U78 ( .A(n821), .B(n640), .C(n473), .Y(n300) );
  OAI21X1 U80 ( .A(n820), .B(n640), .C(n471), .Y(n301) );
  OAI21X1 U82 ( .A(n819), .B(n640), .C(n469), .Y(n302) );
  OAI21X1 U86 ( .A(n823), .B(n638), .C(n467), .Y(n303) );
  OAI21X1 U88 ( .A(n822), .B(n638), .C(n465), .Y(n304) );
  OAI21X1 U90 ( .A(n821), .B(n638), .C(n463), .Y(n305) );
  OAI21X1 U92 ( .A(n820), .B(n638), .C(n461), .Y(n306) );
  OAI21X1 U94 ( .A(n819), .B(n638), .C(n459), .Y(n307) );
  OAI21X1 U98 ( .A(n823), .B(n636), .C(n457), .Y(n308) );
  OAI21X1 U100 ( .A(n822), .B(n636), .C(n455), .Y(n309) );
  OAI21X1 U102 ( .A(n821), .B(n636), .C(n453), .Y(n310) );
  OAI21X1 U104 ( .A(n820), .B(n636), .C(n451), .Y(n311) );
  OAI21X1 U106 ( .A(n819), .B(n636), .C(n449), .Y(n312) );
  OAI21X1 U110 ( .A(n823), .B(n634), .C(n287), .Y(n313) );
  OAI21X1 U112 ( .A(n822), .B(n634), .C(n284), .Y(n314) );
  OAI21X1 U114 ( .A(n821), .B(n634), .C(n282), .Y(n315) );
  OAI21X1 U116 ( .A(n820), .B(n634), .C(n280), .Y(n316) );
  OAI21X1 U118 ( .A(n819), .B(n634), .C(n278), .Y(n317) );
  OAI21X1 U122 ( .A(n823), .B(n632), .C(n276), .Y(n318) );
  OAI21X1 U124 ( .A(n822), .B(n632), .C(n274), .Y(n319) );
  OAI21X1 U126 ( .A(n821), .B(n632), .C(n272), .Y(n320) );
  OAI21X1 U128 ( .A(n820), .B(n632), .C(n270), .Y(n321) );
  OAI21X1 U130 ( .A(n819), .B(n632), .C(n268), .Y(n322) );
  OAI21X1 U134 ( .A(n823), .B(n630), .C(n266), .Y(n323) );
  OAI21X1 U136 ( .A(n822), .B(n630), .C(n264), .Y(n324) );
  OAI21X1 U138 ( .A(n821), .B(n630), .C(n262), .Y(n325) );
  OAI21X1 U140 ( .A(n820), .B(n630), .C(n260), .Y(n326) );
  OAI21X1 U142 ( .A(n819), .B(n630), .C(n258), .Y(n327) );
  NAND3X1 U146 ( .A(N13), .B(n115), .C(N14), .Y(n114) );
  OAI21X1 U147 ( .A(n823), .B(n628), .C(n256), .Y(n328) );
  OAI21X1 U149 ( .A(n822), .B(n628), .C(n254), .Y(n329) );
  OAI21X1 U151 ( .A(n821), .B(n628), .C(n252), .Y(n330) );
  OAI21X1 U153 ( .A(n820), .B(n628), .C(n250), .Y(n331) );
  OAI21X1 U155 ( .A(n819), .B(n628), .C(n248), .Y(n332) );
  OAI21X1 U159 ( .A(n823), .B(n626), .C(n246), .Y(n333) );
  OAI21X1 U161 ( .A(n822), .B(n626), .C(n244), .Y(n334) );
  OAI21X1 U163 ( .A(n821), .B(n626), .C(n242), .Y(n335) );
  OAI21X1 U165 ( .A(n820), .B(n626), .C(n240), .Y(n336) );
  OAI21X1 U167 ( .A(n819), .B(n626), .C(n238), .Y(n337) );
  OAI21X1 U171 ( .A(n823), .B(n623), .C(n236), .Y(n338) );
  OAI21X1 U173 ( .A(n822), .B(n623), .C(n234), .Y(n339) );
  OAI21X1 U175 ( .A(n821), .B(n623), .C(n232), .Y(n340) );
  OAI21X1 U177 ( .A(n820), .B(n623), .C(n230), .Y(n341) );
  OAI21X1 U179 ( .A(n819), .B(n623), .C(n227), .Y(n342) );
  OAI21X1 U183 ( .A(n823), .B(n622), .C(n225), .Y(n343) );
  OAI21X1 U185 ( .A(n822), .B(n622), .C(n223), .Y(n344) );
  OAI21X1 U187 ( .A(n821), .B(n622), .C(n221), .Y(n345) );
  OAI21X1 U189 ( .A(n820), .B(n622), .C(n219), .Y(n346) );
  OAI21X1 U191 ( .A(n819), .B(n622), .C(n217), .Y(n347) );
  OAI21X1 U195 ( .A(n823), .B(n619), .C(n215), .Y(n348) );
  OAI21X1 U197 ( .A(n822), .B(n619), .C(n213), .Y(n349) );
  OAI21X1 U199 ( .A(n821), .B(n619), .C(n211), .Y(n350) );
  OAI21X1 U201 ( .A(n820), .B(n619), .C(n209), .Y(n351) );
  OAI21X1 U203 ( .A(n819), .B(n619), .C(n207), .Y(n352) );
  OAI21X1 U207 ( .A(n823), .B(n618), .C(n205), .Y(n353) );
  OAI21X1 U209 ( .A(n822), .B(n618), .C(n203), .Y(n354) );
  OAI21X1 U211 ( .A(n821), .B(n618), .C(n201), .Y(n355) );
  OAI21X1 U213 ( .A(n820), .B(n618), .C(n199), .Y(n356) );
  OAI21X1 U215 ( .A(n819), .B(n618), .C(n197), .Y(n357) );
  OAI21X1 U219 ( .A(n823), .B(n616), .C(n195), .Y(n358) );
  OAI21X1 U221 ( .A(n822), .B(n616), .C(n193), .Y(n359) );
  OAI21X1 U223 ( .A(n821), .B(n616), .C(n191), .Y(n360) );
  OAI21X1 U225 ( .A(n820), .B(n616), .C(n189), .Y(n361) );
  OAI21X1 U227 ( .A(n819), .B(n616), .C(n187), .Y(n362) );
  OAI21X1 U231 ( .A(n823), .B(n614), .C(n185), .Y(n363) );
  OAI21X1 U233 ( .A(n822), .B(n614), .C(n183), .Y(n364) );
  OAI21X1 U235 ( .A(n821), .B(n614), .C(n181), .Y(n365) );
  OAI21X1 U237 ( .A(n820), .B(n614), .C(n179), .Y(n366) );
  OAI21X1 U239 ( .A(n819), .B(n614), .C(n177), .Y(n367) );
  NAND3X1 U243 ( .A(n115), .B(n830), .C(N14), .Y(n172) );
  OAI21X1 U244 ( .A(n823), .B(n611), .C(n175), .Y(n368) );
  OAI21X1 U246 ( .A(n822), .B(n611), .C(n173), .Y(n369) );
  OAI21X1 U248 ( .A(n821), .B(n611), .C(n170), .Y(n370) );
  OAI21X1 U250 ( .A(n820), .B(n611), .C(n168), .Y(n371) );
  OAI21X1 U252 ( .A(n819), .B(n611), .C(n166), .Y(n372) );
  OAI21X1 U256 ( .A(n823), .B(n609), .C(n164), .Y(n373) );
  OAI21X1 U258 ( .A(n822), .B(n609), .C(n162), .Y(n374) );
  OAI21X1 U260 ( .A(n821), .B(n609), .C(n160), .Y(n375) );
  OAI21X1 U262 ( .A(n820), .B(n609), .C(n158), .Y(n376) );
  OAI21X1 U264 ( .A(n819), .B(n609), .C(n156), .Y(n377) );
  OAI21X1 U268 ( .A(n823), .B(n608), .C(n154), .Y(n378) );
  OAI21X1 U270 ( .A(n822), .B(n608), .C(n152), .Y(n379) );
  OAI21X1 U272 ( .A(n821), .B(n608), .C(n150), .Y(n380) );
  OAI21X1 U274 ( .A(n820), .B(n608), .C(n148), .Y(n381) );
  OAI21X1 U276 ( .A(n819), .B(n608), .C(n146), .Y(n382) );
  OAI21X1 U280 ( .A(n823), .B(n606), .C(n144), .Y(n383) );
  OAI21X1 U282 ( .A(n822), .B(n606), .C(n142), .Y(n384) );
  OAI21X1 U284 ( .A(n821), .B(n606), .C(n140), .Y(n385) );
  OAI21X1 U286 ( .A(n820), .B(n606), .C(n138), .Y(n386) );
  OAI21X1 U288 ( .A(n819), .B(n606), .C(n136), .Y(n387) );
  OAI21X1 U292 ( .A(n823), .B(n604), .C(n134), .Y(n388) );
  OAI21X1 U294 ( .A(n822), .B(n604), .C(n132), .Y(n389) );
  OAI21X1 U296 ( .A(n821), .B(n604), .C(n130), .Y(n390) );
  OAI21X1 U298 ( .A(n820), .B(n604), .C(n128), .Y(n391) );
  OAI21X1 U300 ( .A(n819), .B(n604), .C(n126), .Y(n392) );
  OAI21X1 U304 ( .A(n823), .B(n601), .C(n124), .Y(n393) );
  OAI21X1 U306 ( .A(n822), .B(n601), .C(n122), .Y(n394) );
  OAI21X1 U308 ( .A(n821), .B(n601), .C(n120), .Y(n395) );
  OAI21X1 U310 ( .A(n820), .B(n601), .C(n118), .Y(n396) );
  OAI21X1 U312 ( .A(n819), .B(n601), .C(n116), .Y(n397) );
  OAI21X1 U316 ( .A(n823), .B(n599), .C(n111), .Y(n398) );
  OAI21X1 U318 ( .A(n822), .B(n599), .C(n109), .Y(n399) );
  OAI21X1 U320 ( .A(n821), .B(n599), .C(n107), .Y(n400) );
  OAI21X1 U322 ( .A(n820), .B(n599), .C(n104), .Y(n401) );
  OAI21X1 U324 ( .A(n819), .B(n599), .C(n102), .Y(n402) );
  OAI21X1 U328 ( .A(n823), .B(n597), .C(n100), .Y(n403) );
  OAI21X1 U330 ( .A(n822), .B(n597), .C(n98), .Y(n404) );
  OAI21X1 U332 ( .A(n821), .B(n597), .C(n95), .Y(n405) );
  OAI21X1 U334 ( .A(n820), .B(n597), .C(n93), .Y(n406) );
  OAI21X1 U336 ( .A(n819), .B(n597), .C(n91), .Y(n407) );
  NAND3X1 U340 ( .A(n115), .B(n831), .C(N13), .Y(n229) );
  OAI21X1 U341 ( .A(n823), .B(n595), .C(n88), .Y(n408) );
  OAI21X1 U343 ( .A(n822), .B(n595), .C(n86), .Y(n409) );
  OAI21X1 U345 ( .A(n821), .B(n595), .C(n84), .Y(n410) );
  OAI21X1 U347 ( .A(n820), .B(n595), .C(n82), .Y(n411) );
  OAI21X1 U349 ( .A(n819), .B(n595), .C(n79), .Y(n412) );
  NOR3X1 U353 ( .A(n827), .B(n818), .C(n829), .Y(n57) );
  OAI21X1 U354 ( .A(n823), .B(n593), .C(n77), .Y(n413) );
  OAI21X1 U356 ( .A(n822), .B(n593), .C(n75), .Y(n414) );
  OAI21X1 U358 ( .A(n821), .B(n593), .C(n72), .Y(n415) );
  OAI21X1 U360 ( .A(n820), .B(n593), .C(n70), .Y(n416) );
  OAI21X1 U362 ( .A(n819), .B(n593), .C(n68), .Y(n417) );
  NOR3X1 U366 ( .A(n827), .B(n816), .C(n829), .Y(n65) );
  OAI21X1 U367 ( .A(n823), .B(n592), .C(n66), .Y(n418) );
  OAI21X1 U369 ( .A(n822), .B(n592), .C(n63), .Y(n419) );
  OAI21X1 U371 ( .A(n821), .B(n592), .C(n61), .Y(n420) );
  OAI21X1 U373 ( .A(n820), .B(n592), .C(n59), .Y(n421) );
  OAI21X1 U375 ( .A(n819), .B(n592), .C(n55), .Y(n422) );
  NOR3X1 U379 ( .A(n818), .B(N11), .C(n829), .Y(n73) );
  OAI21X1 U380 ( .A(n823), .B(n590), .C(n53), .Y(n423) );
  OAI21X1 U382 ( .A(n822), .B(n590), .C(n51), .Y(n424) );
  OAI21X1 U384 ( .A(n821), .B(n590), .C(n49), .Y(n425) );
  OAI21X1 U386 ( .A(n820), .B(n590), .C(n47), .Y(n426) );
  OAI21X1 U388 ( .A(n819), .B(n590), .C(n45), .Y(n427) );
  NOR3X1 U392 ( .A(n825), .B(N11), .C(n829), .Y(n81) );
  OAI21X1 U393 ( .A(n823), .B(n588), .C(n43), .Y(n428) );
  OAI21X1 U395 ( .A(n822), .B(n588), .C(n41), .Y(n429) );
  OAI21X1 U397 ( .A(n821), .B(n588), .C(n39), .Y(n430) );
  OAI21X1 U399 ( .A(n820), .B(n588), .C(n37), .Y(n431) );
  OAI21X1 U401 ( .A(n819), .B(n588), .C(n35), .Y(n432) );
  NOR3X1 U405 ( .A(n818), .B(n828), .C(n827), .Y(n89) );
  OAI21X1 U406 ( .A(n823), .B(n586), .C(n33), .Y(n433) );
  OAI21X1 U408 ( .A(n822), .B(n586), .C(n31), .Y(n434) );
  OAI21X1 U410 ( .A(n821), .B(n586), .C(n29), .Y(n435) );
  OAI21X1 U412 ( .A(n820), .B(n586), .C(n27), .Y(n436) );
  OAI21X1 U414 ( .A(n819), .B(n586), .C(n25), .Y(n437) );
  NOR3X1 U418 ( .A(n816), .B(n828), .C(n827), .Y(n97) );
  OAI21X1 U419 ( .A(n823), .B(n584), .C(n23), .Y(n438) );
  OAI21X1 U421 ( .A(n822), .B(n584), .C(n21), .Y(n439) );
  OAI21X1 U423 ( .A(n821), .B(n584), .C(n19), .Y(n440) );
  OAI21X1 U425 ( .A(n820), .B(n584), .C(n17), .Y(n441) );
  OAI21X1 U427 ( .A(n819), .B(n584), .C(n15), .Y(n442) );
  NOR3X1 U431 ( .A(N11), .B(n828), .C(n818), .Y(n105) );
  OAI21X1 U432 ( .A(n823), .B(n582), .C(n13), .Y(n443) );
  OAI21X1 U435 ( .A(n822), .B(n582), .C(n11), .Y(n444) );
  OAI21X1 U438 ( .A(n821), .B(n582), .C(n9), .Y(n445) );
  OAI21X1 U441 ( .A(n820), .B(n582), .C(n7), .Y(n446) );
  OAI21X1 U444 ( .A(n819), .B(n582), .C(n5), .Y(n447) );
  NOR3X1 U448 ( .A(N11), .B(n828), .C(n816), .Y(n113) );
  NAND3X1 U449 ( .A(n830), .B(n831), .C(n115), .Y(n286) );
  NOR3X1 U450 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n115) );
  INVX2 U3 ( .A(n514), .Y(n823) );
  INVX2 U4 ( .A(n513), .Y(n822) );
  INVX2 U5 ( .A(n512), .Y(n821) );
  INVX2 U6 ( .A(n511), .Y(n820) );
  INVX2 U7 ( .A(n510), .Y(n819) );
  AND2X1 U8 ( .A(\mem<31><4> ), .B(n578), .Y(n488) );
  AND2X1 U9 ( .A(\mem<30><4> ), .B(n576), .Y(n478) );
  AND2X1 U10 ( .A(\mem<29><4> ), .B(n574), .Y(n468) );
  AND2X1 U11 ( .A(\mem<28><4> ), .B(n572), .Y(n458) );
  AND2X1 U12 ( .A(\mem<27><4> ), .B(n570), .Y(n448) );
  AND2X1 U13 ( .A(\mem<26><4> ), .B(n568), .Y(n277) );
  AND2X1 U14 ( .A(\mem<25><4> ), .B(n566), .Y(n267) );
  AND2X1 U15 ( .A(\mem<24><4> ), .B(n564), .Y(n257) );
  AND2X1 U16 ( .A(\mem<23><4> ), .B(n562), .Y(n247) );
  AND2X1 U17 ( .A(\mem<22><4> ), .B(n560), .Y(n237) );
  AND2X1 U18 ( .A(\mem<21><4> ), .B(n558), .Y(n226) );
  AND2X1 U19 ( .A(\mem<20><4> ), .B(n556), .Y(n216) );
  AND2X1 U20 ( .A(\mem<19><4> ), .B(n554), .Y(n206) );
  AND2X1 U21 ( .A(\mem<18><4> ), .B(n552), .Y(n196) );
  AND2X1 U22 ( .A(\mem<17><4> ), .B(n550), .Y(n186) );
  AND2X1 U23 ( .A(\mem<16><4> ), .B(n548), .Y(n176) );
  AND2X1 U24 ( .A(\mem<15><4> ), .B(n546), .Y(n165) );
  AND2X1 U25 ( .A(\mem<14><4> ), .B(n544), .Y(n155) );
  AND2X1 U26 ( .A(\mem<13><4> ), .B(n542), .Y(n145) );
  AND2X1 U27 ( .A(\mem<12><4> ), .B(n540), .Y(n135) );
  AND2X1 U28 ( .A(\mem<10><4> ), .B(n536), .Y(n112) );
  AND2X1 U29 ( .A(\mem<9><4> ), .B(n534), .Y(n101) );
  AND2X1 U30 ( .A(\mem<8><4> ), .B(n532), .Y(n90) );
  AND2X1 U31 ( .A(\mem<7><4> ), .B(n530), .Y(n78) );
  AND2X1 U32 ( .A(\mem<6><4> ), .B(n528), .Y(n67) );
  AND2X1 U33 ( .A(\mem<5><4> ), .B(n526), .Y(n54) );
  AND2X1 U34 ( .A(\mem<4><4> ), .B(n524), .Y(n44) );
  AND2X1 U35 ( .A(\mem<3><4> ), .B(n522), .Y(n34) );
  AND2X1 U36 ( .A(\mem<2><4> ), .B(n520), .Y(n24) );
  AND2X1 U37 ( .A(\mem<1><4> ), .B(n518), .Y(n14) );
  AND2X1 U38 ( .A(\mem<0><4> ), .B(n516), .Y(n4) );
  INVX1 U39 ( .A(N14), .Y(n831) );
  INVX1 U40 ( .A(N11), .Y(n827) );
  INVX1 U41 ( .A(rst), .Y(n824) );
  INVX4 U42 ( .A(n644), .Y(n810) );
  INVX1 U43 ( .A(n829), .Y(n828) );
  INVX1 U44 ( .A(N13), .Y(n830) );
  OR2X2 U45 ( .A(write), .B(rst), .Y(n1) );
  AND2X2 U46 ( .A(n501), .B(n499), .Y(n2) );
  AND2X2 U47 ( .A(n646), .B(n647), .Y(n3) );
  INVX1 U48 ( .A(n4), .Y(n5) );
  AND2X2 U49 ( .A(\mem<0><3> ), .B(n516), .Y(n6) );
  INVX1 U51 ( .A(n6), .Y(n7) );
  AND2X2 U53 ( .A(\mem<0><2> ), .B(n516), .Y(n8) );
  INVX1 U55 ( .A(n8), .Y(n9) );
  AND2X2 U57 ( .A(\mem<0><1> ), .B(n516), .Y(n10) );
  INVX1 U59 ( .A(n10), .Y(n11) );
  AND2X2 U60 ( .A(\mem<0><0> ), .B(n516), .Y(n12) );
  INVX1 U61 ( .A(n12), .Y(n13) );
  INVX1 U63 ( .A(n14), .Y(n15) );
  AND2X2 U65 ( .A(\mem<1><3> ), .B(n518), .Y(n16) );
  INVX1 U67 ( .A(n16), .Y(n17) );
  AND2X2 U69 ( .A(\mem<1><2> ), .B(n518), .Y(n18) );
  INVX1 U71 ( .A(n18), .Y(n19) );
  AND2X2 U72 ( .A(\mem<1><1> ), .B(n518), .Y(n20) );
  INVX1 U73 ( .A(n20), .Y(n21) );
  AND2X2 U75 ( .A(\mem<1><0> ), .B(n518), .Y(n22) );
  INVX1 U77 ( .A(n22), .Y(n23) );
  INVX1 U79 ( .A(n24), .Y(n25) );
  AND2X2 U81 ( .A(\mem<2><3> ), .B(n520), .Y(n26) );
  INVX1 U83 ( .A(n26), .Y(n27) );
  AND2X2 U84 ( .A(\mem<2><2> ), .B(n520), .Y(n28) );
  INVX1 U85 ( .A(n28), .Y(n29) );
  AND2X2 U87 ( .A(\mem<2><1> ), .B(n520), .Y(n30) );
  INVX1 U89 ( .A(n30), .Y(n31) );
  AND2X2 U91 ( .A(\mem<2><0> ), .B(n520), .Y(n32) );
  INVX1 U93 ( .A(n32), .Y(n33) );
  INVX1 U95 ( .A(n34), .Y(n35) );
  AND2X2 U96 ( .A(\mem<3><3> ), .B(n522), .Y(n36) );
  INVX1 U97 ( .A(n36), .Y(n37) );
  AND2X2 U99 ( .A(\mem<3><2> ), .B(n522), .Y(n38) );
  INVX1 U101 ( .A(n38), .Y(n39) );
  AND2X2 U103 ( .A(\mem<3><1> ), .B(n522), .Y(n40) );
  INVX1 U105 ( .A(n40), .Y(n41) );
  AND2X2 U107 ( .A(\mem<3><0> ), .B(n522), .Y(n42) );
  INVX1 U108 ( .A(n42), .Y(n43) );
  INVX1 U109 ( .A(n44), .Y(n45) );
  AND2X2 U111 ( .A(\mem<4><3> ), .B(n524), .Y(n46) );
  INVX1 U113 ( .A(n46), .Y(n47) );
  AND2X2 U115 ( .A(\mem<4><2> ), .B(n524), .Y(n48) );
  INVX1 U117 ( .A(n48), .Y(n49) );
  AND2X2 U119 ( .A(\mem<4><1> ), .B(n524), .Y(n50) );
  INVX1 U120 ( .A(n50), .Y(n51) );
  AND2X2 U121 ( .A(\mem<4><0> ), .B(n524), .Y(n52) );
  INVX1 U123 ( .A(n52), .Y(n53) );
  INVX1 U125 ( .A(n54), .Y(n55) );
  AND2X2 U127 ( .A(\mem<5><3> ), .B(n526), .Y(n58) );
  INVX1 U129 ( .A(n58), .Y(n59) );
  AND2X2 U131 ( .A(\mem<5><2> ), .B(n526), .Y(n60) );
  INVX1 U132 ( .A(n60), .Y(n61) );
  AND2X2 U133 ( .A(\mem<5><1> ), .B(n526), .Y(n62) );
  INVX1 U135 ( .A(n62), .Y(n63) );
  AND2X2 U137 ( .A(\mem<5><0> ), .B(n526), .Y(n64) );
  INVX1 U139 ( .A(n64), .Y(n66) );
  INVX1 U141 ( .A(n67), .Y(n68) );
  AND2X2 U143 ( .A(\mem<6><3> ), .B(n528), .Y(n69) );
  INVX1 U144 ( .A(n69), .Y(n70) );
  AND2X2 U145 ( .A(\mem<6><2> ), .B(n528), .Y(n71) );
  INVX1 U148 ( .A(n71), .Y(n72) );
  AND2X2 U150 ( .A(\mem<6><1> ), .B(n528), .Y(n74) );
  INVX1 U152 ( .A(n74), .Y(n75) );
  AND2X2 U154 ( .A(\mem<6><0> ), .B(n528), .Y(n76) );
  INVX1 U156 ( .A(n76), .Y(n77) );
  INVX1 U157 ( .A(n78), .Y(n79) );
  AND2X2 U158 ( .A(\mem<7><3> ), .B(n530), .Y(n80) );
  INVX1 U160 ( .A(n80), .Y(n82) );
  AND2X2 U162 ( .A(\mem<7><2> ), .B(n530), .Y(n83) );
  INVX1 U164 ( .A(n83), .Y(n84) );
  AND2X2 U166 ( .A(\mem<7><1> ), .B(n530), .Y(n85) );
  INVX1 U168 ( .A(n85), .Y(n86) );
  AND2X2 U169 ( .A(\mem<7><0> ), .B(n530), .Y(n87) );
  INVX1 U170 ( .A(n87), .Y(n88) );
  INVX1 U172 ( .A(n90), .Y(n91) );
  AND2X2 U174 ( .A(\mem<8><3> ), .B(n532), .Y(n92) );
  INVX1 U176 ( .A(n92), .Y(n93) );
  AND2X2 U178 ( .A(\mem<8><2> ), .B(n532), .Y(n94) );
  INVX1 U180 ( .A(n94), .Y(n95) );
  AND2X2 U181 ( .A(\mem<8><1> ), .B(n532), .Y(n96) );
  INVX1 U182 ( .A(n96), .Y(n98) );
  AND2X2 U184 ( .A(\mem<8><0> ), .B(n532), .Y(n99) );
  INVX1 U186 ( .A(n99), .Y(n100) );
  INVX1 U188 ( .A(n101), .Y(n102) );
  AND2X2 U190 ( .A(\mem<9><3> ), .B(n534), .Y(n103) );
  INVX1 U192 ( .A(n103), .Y(n104) );
  AND2X2 U193 ( .A(\mem<9><2> ), .B(n534), .Y(n106) );
  INVX1 U194 ( .A(n106), .Y(n107) );
  AND2X2 U196 ( .A(\mem<9><1> ), .B(n534), .Y(n108) );
  INVX1 U198 ( .A(n108), .Y(n109) );
  AND2X2 U200 ( .A(\mem<9><0> ), .B(n534), .Y(n110) );
  INVX1 U202 ( .A(n110), .Y(n111) );
  INVX1 U204 ( .A(n112), .Y(n116) );
  AND2X2 U205 ( .A(\mem<10><3> ), .B(n536), .Y(n117) );
  INVX1 U206 ( .A(n117), .Y(n118) );
  AND2X2 U208 ( .A(\mem<10><2> ), .B(n536), .Y(n119) );
  INVX1 U210 ( .A(n119), .Y(n120) );
  AND2X2 U212 ( .A(\mem<10><1> ), .B(n536), .Y(n121) );
  INVX1 U214 ( .A(n121), .Y(n122) );
  AND2X2 U216 ( .A(\mem<10><0> ), .B(n536), .Y(n123) );
  INVX1 U217 ( .A(n123), .Y(n124) );
  AND2X2 U218 ( .A(\mem<11><4> ), .B(n538), .Y(n125) );
  INVX1 U220 ( .A(n125), .Y(n126) );
  AND2X2 U222 ( .A(\mem<11><3> ), .B(n538), .Y(n127) );
  INVX1 U224 ( .A(n127), .Y(n128) );
  AND2X2 U226 ( .A(\mem<11><2> ), .B(n538), .Y(n129) );
  INVX1 U228 ( .A(n129), .Y(n130) );
  AND2X2 U229 ( .A(\mem<11><1> ), .B(n538), .Y(n131) );
  INVX1 U230 ( .A(n131), .Y(n132) );
  AND2X2 U232 ( .A(\mem<11><0> ), .B(n538), .Y(n133) );
  INVX1 U234 ( .A(n133), .Y(n134) );
  INVX1 U236 ( .A(n135), .Y(n136) );
  AND2X2 U238 ( .A(\mem<12><3> ), .B(n540), .Y(n137) );
  INVX1 U240 ( .A(n137), .Y(n138) );
  AND2X2 U241 ( .A(\mem<12><2> ), .B(n540), .Y(n139) );
  INVX1 U242 ( .A(n139), .Y(n140) );
  AND2X2 U245 ( .A(\mem<12><1> ), .B(n540), .Y(n141) );
  INVX1 U247 ( .A(n141), .Y(n142) );
  AND2X2 U249 ( .A(\mem<12><0> ), .B(n540), .Y(n143) );
  INVX1 U251 ( .A(n143), .Y(n144) );
  INVX1 U253 ( .A(n145), .Y(n146) );
  AND2X2 U254 ( .A(\mem<13><3> ), .B(n542), .Y(n147) );
  INVX1 U255 ( .A(n147), .Y(n148) );
  AND2X2 U257 ( .A(\mem<13><2> ), .B(n542), .Y(n149) );
  INVX1 U259 ( .A(n149), .Y(n150) );
  AND2X2 U261 ( .A(\mem<13><1> ), .B(n542), .Y(n151) );
  INVX1 U263 ( .A(n151), .Y(n152) );
  AND2X2 U265 ( .A(\mem<13><0> ), .B(n542), .Y(n153) );
  INVX1 U266 ( .A(n153), .Y(n154) );
  INVX1 U267 ( .A(n155), .Y(n156) );
  AND2X2 U269 ( .A(\mem<14><3> ), .B(n544), .Y(n157) );
  INVX1 U271 ( .A(n157), .Y(n158) );
  AND2X2 U273 ( .A(\mem<14><2> ), .B(n544), .Y(n159) );
  INVX1 U275 ( .A(n159), .Y(n160) );
  AND2X2 U277 ( .A(\mem<14><1> ), .B(n544), .Y(n161) );
  INVX1 U278 ( .A(n161), .Y(n162) );
  AND2X2 U279 ( .A(\mem<14><0> ), .B(n544), .Y(n163) );
  INVX1 U281 ( .A(n163), .Y(n164) );
  INVX1 U283 ( .A(n165), .Y(n166) );
  AND2X2 U285 ( .A(\mem<15><3> ), .B(n546), .Y(n167) );
  INVX1 U287 ( .A(n167), .Y(n168) );
  AND2X2 U289 ( .A(\mem<15><2> ), .B(n546), .Y(n169) );
  INVX1 U290 ( .A(n169), .Y(n170) );
  AND2X2 U291 ( .A(\mem<15><1> ), .B(n546), .Y(n171) );
  INVX1 U293 ( .A(n171), .Y(n173) );
  AND2X2 U295 ( .A(\mem<15><0> ), .B(n546), .Y(n174) );
  INVX1 U297 ( .A(n174), .Y(n175) );
  INVX1 U299 ( .A(n176), .Y(n177) );
  AND2X2 U301 ( .A(\mem<16><3> ), .B(n548), .Y(n178) );
  INVX1 U302 ( .A(n178), .Y(n179) );
  AND2X2 U303 ( .A(\mem<16><2> ), .B(n548), .Y(n180) );
  INVX1 U305 ( .A(n180), .Y(n181) );
  AND2X2 U307 ( .A(\mem<16><1> ), .B(n548), .Y(n182) );
  INVX1 U309 ( .A(n182), .Y(n183) );
  AND2X2 U311 ( .A(\mem<16><0> ), .B(n548), .Y(n184) );
  INVX1 U313 ( .A(n184), .Y(n185) );
  INVX1 U314 ( .A(n186), .Y(n187) );
  AND2X2 U315 ( .A(\mem<17><3> ), .B(n550), .Y(n188) );
  INVX1 U317 ( .A(n188), .Y(n189) );
  AND2X2 U319 ( .A(\mem<17><2> ), .B(n550), .Y(n190) );
  INVX1 U321 ( .A(n190), .Y(n191) );
  AND2X2 U323 ( .A(\mem<17><1> ), .B(n550), .Y(n192) );
  INVX1 U325 ( .A(n192), .Y(n193) );
  AND2X2 U326 ( .A(\mem<17><0> ), .B(n550), .Y(n194) );
  INVX1 U327 ( .A(n194), .Y(n195) );
  INVX1 U329 ( .A(n196), .Y(n197) );
  AND2X2 U331 ( .A(\mem<18><3> ), .B(n552), .Y(n198) );
  INVX1 U333 ( .A(n198), .Y(n199) );
  AND2X2 U335 ( .A(\mem<18><2> ), .B(n552), .Y(n200) );
  INVX1 U337 ( .A(n200), .Y(n201) );
  AND2X2 U338 ( .A(\mem<18><1> ), .B(n552), .Y(n202) );
  INVX1 U339 ( .A(n202), .Y(n203) );
  AND2X2 U342 ( .A(\mem<18><0> ), .B(n552), .Y(n204) );
  INVX1 U344 ( .A(n204), .Y(n205) );
  INVX1 U346 ( .A(n206), .Y(n207) );
  AND2X2 U348 ( .A(\mem<19><3> ), .B(n554), .Y(n208) );
  INVX1 U350 ( .A(n208), .Y(n209) );
  AND2X2 U351 ( .A(\mem<19><2> ), .B(n554), .Y(n210) );
  INVX1 U352 ( .A(n210), .Y(n211) );
  AND2X2 U355 ( .A(\mem<19><1> ), .B(n554), .Y(n212) );
  INVX1 U357 ( .A(n212), .Y(n213) );
  AND2X2 U359 ( .A(\mem<19><0> ), .B(n554), .Y(n214) );
  INVX1 U361 ( .A(n214), .Y(n215) );
  INVX1 U363 ( .A(n216), .Y(n217) );
  AND2X2 U364 ( .A(\mem<20><3> ), .B(n556), .Y(n218) );
  INVX1 U365 ( .A(n218), .Y(n219) );
  AND2X2 U368 ( .A(\mem<20><2> ), .B(n556), .Y(n220) );
  INVX1 U370 ( .A(n220), .Y(n221) );
  AND2X2 U372 ( .A(\mem<20><1> ), .B(n556), .Y(n222) );
  INVX1 U374 ( .A(n222), .Y(n223) );
  AND2X2 U376 ( .A(\mem<20><0> ), .B(n556), .Y(n224) );
  INVX1 U377 ( .A(n224), .Y(n225) );
  INVX1 U378 ( .A(n226), .Y(n227) );
  AND2X2 U381 ( .A(\mem<21><3> ), .B(n558), .Y(n228) );
  INVX1 U383 ( .A(n228), .Y(n230) );
  AND2X2 U385 ( .A(\mem<21><2> ), .B(n558), .Y(n231) );
  INVX1 U387 ( .A(n231), .Y(n232) );
  AND2X2 U389 ( .A(\mem<21><1> ), .B(n558), .Y(n233) );
  INVX1 U390 ( .A(n233), .Y(n234) );
  AND2X2 U391 ( .A(\mem<21><0> ), .B(n558), .Y(n235) );
  INVX1 U394 ( .A(n235), .Y(n236) );
  INVX1 U396 ( .A(n237), .Y(n238) );
  AND2X2 U398 ( .A(\mem<22><3> ), .B(n560), .Y(n239) );
  INVX1 U400 ( .A(n239), .Y(n240) );
  AND2X2 U402 ( .A(\mem<22><2> ), .B(n560), .Y(n241) );
  INVX1 U403 ( .A(n241), .Y(n242) );
  AND2X2 U404 ( .A(\mem<22><1> ), .B(n560), .Y(n243) );
  INVX1 U407 ( .A(n243), .Y(n244) );
  AND2X2 U409 ( .A(\mem<22><0> ), .B(n560), .Y(n245) );
  INVX1 U411 ( .A(n245), .Y(n246) );
  INVX1 U413 ( .A(n247), .Y(n248) );
  AND2X2 U415 ( .A(\mem<23><3> ), .B(n562), .Y(n249) );
  INVX1 U416 ( .A(n249), .Y(n250) );
  AND2X2 U417 ( .A(\mem<23><2> ), .B(n562), .Y(n251) );
  INVX1 U420 ( .A(n251), .Y(n252) );
  AND2X2 U422 ( .A(\mem<23><1> ), .B(n562), .Y(n253) );
  INVX1 U424 ( .A(n253), .Y(n254) );
  AND2X2 U426 ( .A(\mem<23><0> ), .B(n562), .Y(n255) );
  INVX1 U428 ( .A(n255), .Y(n256) );
  INVX1 U429 ( .A(n257), .Y(n258) );
  AND2X2 U430 ( .A(\mem<24><3> ), .B(n564), .Y(n259) );
  INVX1 U433 ( .A(n259), .Y(n260) );
  AND2X2 U434 ( .A(\mem<24><2> ), .B(n564), .Y(n261) );
  INVX1 U436 ( .A(n261), .Y(n262) );
  AND2X2 U437 ( .A(\mem<24><1> ), .B(n564), .Y(n263) );
  INVX1 U439 ( .A(n263), .Y(n264) );
  AND2X2 U440 ( .A(\mem<24><0> ), .B(n564), .Y(n265) );
  INVX1 U442 ( .A(n265), .Y(n266) );
  INVX1 U443 ( .A(n267), .Y(n268) );
  AND2X2 U445 ( .A(\mem<25><3> ), .B(n566), .Y(n269) );
  INVX1 U446 ( .A(n269), .Y(n270) );
  AND2X2 U447 ( .A(\mem<25><2> ), .B(n566), .Y(n271) );
  INVX1 U451 ( .A(n271), .Y(n272) );
  AND2X2 U452 ( .A(\mem<25><1> ), .B(n566), .Y(n273) );
  INVX1 U453 ( .A(n273), .Y(n274) );
  AND2X2 U454 ( .A(\mem<25><0> ), .B(n566), .Y(n275) );
  INVX1 U455 ( .A(n275), .Y(n276) );
  INVX1 U456 ( .A(n277), .Y(n278) );
  AND2X2 U457 ( .A(\mem<26><3> ), .B(n568), .Y(n279) );
  INVX1 U458 ( .A(n279), .Y(n280) );
  AND2X2 U459 ( .A(\mem<26><2> ), .B(n568), .Y(n281) );
  INVX1 U460 ( .A(n281), .Y(n282) );
  AND2X2 U461 ( .A(\mem<26><1> ), .B(n568), .Y(n283) );
  INVX1 U462 ( .A(n283), .Y(n284) );
  AND2X2 U463 ( .A(\mem<26><0> ), .B(n568), .Y(n285) );
  INVX1 U464 ( .A(n285), .Y(n287) );
  INVX1 U465 ( .A(n448), .Y(n449) );
  AND2X2 U466 ( .A(\mem<27><3> ), .B(n570), .Y(n450) );
  INVX1 U467 ( .A(n450), .Y(n451) );
  AND2X2 U468 ( .A(\mem<27><2> ), .B(n570), .Y(n452) );
  INVX1 U469 ( .A(n452), .Y(n453) );
  AND2X2 U470 ( .A(\mem<27><1> ), .B(n570), .Y(n454) );
  INVX1 U471 ( .A(n454), .Y(n455) );
  AND2X2 U472 ( .A(\mem<27><0> ), .B(n570), .Y(n456) );
  INVX1 U473 ( .A(n456), .Y(n457) );
  INVX1 U474 ( .A(n458), .Y(n459) );
  AND2X2 U475 ( .A(\mem<28><3> ), .B(n572), .Y(n460) );
  INVX1 U476 ( .A(n460), .Y(n461) );
  AND2X2 U477 ( .A(\mem<28><2> ), .B(n572), .Y(n462) );
  INVX1 U478 ( .A(n462), .Y(n463) );
  AND2X2 U479 ( .A(\mem<28><1> ), .B(n572), .Y(n464) );
  INVX1 U480 ( .A(n464), .Y(n465) );
  AND2X2 U481 ( .A(\mem<28><0> ), .B(n572), .Y(n466) );
  INVX1 U482 ( .A(n466), .Y(n467) );
  INVX1 U483 ( .A(n468), .Y(n469) );
  AND2X2 U484 ( .A(\mem<29><3> ), .B(n574), .Y(n470) );
  INVX1 U485 ( .A(n470), .Y(n471) );
  AND2X2 U486 ( .A(\mem<29><2> ), .B(n574), .Y(n472) );
  INVX1 U487 ( .A(n472), .Y(n473) );
  AND2X2 U488 ( .A(\mem<29><1> ), .B(n574), .Y(n474) );
  INVX1 U489 ( .A(n474), .Y(n475) );
  AND2X2 U490 ( .A(\mem<29><0> ), .B(n574), .Y(n476) );
  INVX1 U491 ( .A(n476), .Y(n477) );
  INVX1 U492 ( .A(n478), .Y(n479) );
  AND2X2 U493 ( .A(\mem<30><3> ), .B(n576), .Y(n480) );
  INVX1 U494 ( .A(n480), .Y(n481) );
  AND2X2 U495 ( .A(\mem<30><2> ), .B(n576), .Y(n482) );
  INVX1 U496 ( .A(n482), .Y(n483) );
  AND2X2 U497 ( .A(\mem<30><1> ), .B(n576), .Y(n484) );
  INVX1 U498 ( .A(n484), .Y(n485) );
  AND2X2 U499 ( .A(\mem<30><0> ), .B(n576), .Y(n486) );
  INVX1 U500 ( .A(n486), .Y(n487) );
  INVX1 U501 ( .A(n488), .Y(n489) );
  AND2X2 U502 ( .A(\mem<31><3> ), .B(n578), .Y(n490) );
  INVX1 U503 ( .A(n490), .Y(n491) );
  AND2X2 U504 ( .A(\mem<31><2> ), .B(n578), .Y(n492) );
  INVX1 U505 ( .A(n492), .Y(n493) );
  AND2X2 U506 ( .A(\mem<31><1> ), .B(n578), .Y(n494) );
  INVX1 U507 ( .A(n494), .Y(n495) );
  AND2X2 U508 ( .A(\mem<31><0> ), .B(n578), .Y(n496) );
  INVX1 U509 ( .A(n496), .Y(n497) );
  AND2X2 U510 ( .A(n724), .B(n804), .Y(n498) );
  INVX1 U511 ( .A(n498), .Y(n499) );
  AND2X2 U512 ( .A(n727), .B(n643), .Y(n500) );
  INVX1 U513 ( .A(n500), .Y(n501) );
  INVX1 U514 ( .A(n1), .Y(n502) );
  INVX1 U515 ( .A(n1), .Y(n503) );
  OR2X2 U516 ( .A(write), .B(rst), .Y(n504) );
  INVX1 U517 ( .A(n504), .Y(n505) );
  BUFX2 U518 ( .A(n286), .Y(n506) );
  INVX1 U519 ( .A(n506), .Y(n832) );
  BUFX2 U520 ( .A(n229), .Y(n507) );
  INVX1 U521 ( .A(n507), .Y(n833) );
  BUFX2 U522 ( .A(n172), .Y(n508) );
  INVX1 U523 ( .A(n508), .Y(n834) );
  BUFX2 U524 ( .A(n114), .Y(n509) );
  INVX1 U525 ( .A(n509), .Y(n835) );
  AND2X1 U526 ( .A(\data_in<4> ), .B(n56), .Y(n510) );
  AND2X1 U527 ( .A(\data_in<3> ), .B(n56), .Y(n511) );
  AND2X1 U528 ( .A(\data_in<2> ), .B(n56), .Y(n512) );
  AND2X1 U529 ( .A(\data_in<1> ), .B(n56), .Y(n513) );
  AND2X1 U530 ( .A(\data_in<0> ), .B(n56), .Y(n514) );
  AND2X1 U531 ( .A(n581), .B(n56), .Y(n515) );
  INVX1 U532 ( .A(n515), .Y(n516) );
  AND2X1 U533 ( .A(n583), .B(n56), .Y(n517) );
  INVX1 U534 ( .A(n517), .Y(n518) );
  AND2X1 U535 ( .A(n585), .B(n56), .Y(n519) );
  INVX1 U536 ( .A(n519), .Y(n520) );
  AND2X1 U537 ( .A(n587), .B(n56), .Y(n521) );
  INVX1 U538 ( .A(n521), .Y(n522) );
  AND2X1 U539 ( .A(n589), .B(n56), .Y(n523) );
  INVX1 U540 ( .A(n523), .Y(n524) );
  AND2X1 U541 ( .A(n591), .B(n56), .Y(n525) );
  INVX1 U542 ( .A(n525), .Y(n526) );
  AND2X1 U543 ( .A(n594), .B(n56), .Y(n527) );
  INVX1 U544 ( .A(n527), .Y(n528) );
  AND2X1 U545 ( .A(n596), .B(n56), .Y(n529) );
  INVX1 U546 ( .A(n529), .Y(n530) );
  AND2X1 U547 ( .A(n598), .B(n56), .Y(n531) );
  INVX1 U548 ( .A(n531), .Y(n532) );
  AND2X1 U549 ( .A(n600), .B(n56), .Y(n533) );
  INVX1 U550 ( .A(n533), .Y(n534) );
  AND2X1 U551 ( .A(n602), .B(n56), .Y(n535) );
  INVX1 U552 ( .A(n535), .Y(n536) );
  AND2X1 U553 ( .A(n603), .B(n56), .Y(n537) );
  INVX1 U554 ( .A(n537), .Y(n538) );
  AND2X1 U555 ( .A(n605), .B(n56), .Y(n539) );
  INVX1 U556 ( .A(n539), .Y(n540) );
  AND2X1 U557 ( .A(n607), .B(n56), .Y(n541) );
  INVX1 U558 ( .A(n541), .Y(n542) );
  AND2X1 U559 ( .A(n610), .B(n56), .Y(n543) );
  INVX1 U560 ( .A(n543), .Y(n544) );
  AND2X1 U561 ( .A(n612), .B(n56), .Y(n545) );
  INVX1 U562 ( .A(n545), .Y(n546) );
  AND2X1 U563 ( .A(n613), .B(n56), .Y(n547) );
  INVX1 U564 ( .A(n547), .Y(n548) );
  AND2X1 U565 ( .A(n615), .B(n56), .Y(n549) );
  INVX1 U566 ( .A(n549), .Y(n550) );
  AND2X1 U567 ( .A(n617), .B(n56), .Y(n551) );
  INVX1 U568 ( .A(n551), .Y(n552) );
  AND2X1 U569 ( .A(n620), .B(n56), .Y(n553) );
  INVX1 U570 ( .A(n553), .Y(n554) );
  AND2X1 U571 ( .A(n621), .B(n56), .Y(n555) );
  INVX1 U572 ( .A(n555), .Y(n556) );
  AND2X1 U573 ( .A(n624), .B(n56), .Y(n557) );
  INVX1 U574 ( .A(n557), .Y(n558) );
  AND2X1 U575 ( .A(n625), .B(n56), .Y(n559) );
  INVX1 U576 ( .A(n559), .Y(n560) );
  AND2X1 U577 ( .A(n627), .B(n56), .Y(n561) );
  INVX1 U578 ( .A(n561), .Y(n562) );
  AND2X1 U579 ( .A(n629), .B(n56), .Y(n563) );
  INVX1 U580 ( .A(n563), .Y(n564) );
  AND2X1 U581 ( .A(n631), .B(n56), .Y(n565) );
  INVX1 U582 ( .A(n565), .Y(n566) );
  AND2X1 U583 ( .A(n633), .B(n56), .Y(n567) );
  INVX1 U584 ( .A(n567), .Y(n568) );
  AND2X1 U585 ( .A(n635), .B(n56), .Y(n569) );
  INVX1 U586 ( .A(n569), .Y(n570) );
  AND2X1 U587 ( .A(n637), .B(n56), .Y(n571) );
  INVX1 U588 ( .A(n571), .Y(n572) );
  AND2X1 U589 ( .A(n639), .B(n56), .Y(n573) );
  INVX1 U590 ( .A(n573), .Y(n574) );
  AND2X1 U591 ( .A(n641), .B(n56), .Y(n575) );
  INVX1 U592 ( .A(n575), .Y(n576) );
  AND2X1 U593 ( .A(n580), .B(n56), .Y(n577) );
  INVX1 U594 ( .A(n577), .Y(n578) );
  INVX1 U595 ( .A(n580), .Y(n579) );
  AND2X1 U596 ( .A(n57), .B(n835), .Y(n580) );
  AND2X1 U597 ( .A(n832), .B(n113), .Y(n581) );
  INVX1 U598 ( .A(n581), .Y(n582) );
  AND2X1 U599 ( .A(n832), .B(n105), .Y(n583) );
  INVX1 U600 ( .A(n583), .Y(n584) );
  AND2X1 U601 ( .A(n832), .B(n97), .Y(n585) );
  INVX1 U602 ( .A(n585), .Y(n586) );
  AND2X1 U603 ( .A(n832), .B(n89), .Y(n587) );
  INVX1 U604 ( .A(n587), .Y(n588) );
  AND2X1 U605 ( .A(n832), .B(n81), .Y(n589) );
  INVX1 U606 ( .A(n589), .Y(n590) );
  AND2X1 U607 ( .A(n832), .B(n73), .Y(n591) );
  INVX1 U608 ( .A(n591), .Y(n592) );
  INVX1 U609 ( .A(n594), .Y(n593) );
  AND2X1 U610 ( .A(n832), .B(n65), .Y(n594) );
  INVX1 U611 ( .A(n596), .Y(n595) );
  AND2X1 U612 ( .A(n832), .B(n57), .Y(n596) );
  INVX1 U613 ( .A(n598), .Y(n597) );
  AND2X1 U614 ( .A(n833), .B(n113), .Y(n598) );
  INVX1 U615 ( .A(n600), .Y(n599) );
  AND2X1 U616 ( .A(n833), .B(n105), .Y(n600) );
  INVX1 U617 ( .A(n602), .Y(n601) );
  AND2X1 U618 ( .A(n833), .B(n97), .Y(n602) );
  AND2X1 U619 ( .A(n833), .B(n89), .Y(n603) );
  INVX1 U620 ( .A(n603), .Y(n604) );
  AND2X1 U621 ( .A(n833), .B(n81), .Y(n605) );
  INVX1 U622 ( .A(n605), .Y(n606) );
  AND2X1 U623 ( .A(n833), .B(n73), .Y(n607) );
  INVX1 U624 ( .A(n607), .Y(n608) );
  INVX1 U625 ( .A(n610), .Y(n609) );
  AND2X1 U626 ( .A(n833), .B(n65), .Y(n610) );
  INVX1 U627 ( .A(n612), .Y(n611) );
  AND2X1 U628 ( .A(n833), .B(n57), .Y(n612) );
  AND2X1 U629 ( .A(n834), .B(n113), .Y(n613) );
  INVX1 U630 ( .A(n613), .Y(n614) );
  AND2X1 U631 ( .A(n834), .B(n105), .Y(n615) );
  INVX1 U632 ( .A(n615), .Y(n616) );
  AND2X1 U633 ( .A(n834), .B(n97), .Y(n617) );
  INVX1 U634 ( .A(n617), .Y(n618) );
  INVX1 U635 ( .A(n620), .Y(n619) );
  AND2X1 U636 ( .A(n834), .B(n89), .Y(n620) );
  AND2X1 U637 ( .A(n834), .B(n81), .Y(n621) );
  INVX1 U638 ( .A(n621), .Y(n622) );
  INVX1 U639 ( .A(n624), .Y(n623) );
  AND2X1 U640 ( .A(n834), .B(n73), .Y(n624) );
  AND2X1 U641 ( .A(n834), .B(n65), .Y(n625) );
  INVX1 U642 ( .A(n625), .Y(n626) );
  AND2X1 U643 ( .A(n834), .B(n57), .Y(n627) );
  INVX1 U644 ( .A(n627), .Y(n628) );
  AND2X1 U645 ( .A(n113), .B(n835), .Y(n629) );
  INVX1 U646 ( .A(n629), .Y(n630) );
  AND2X1 U647 ( .A(n105), .B(n835), .Y(n631) );
  INVX1 U648 ( .A(n631), .Y(n632) );
  AND2X1 U649 ( .A(n97), .B(n835), .Y(n633) );
  INVX1 U650 ( .A(n633), .Y(n634) );
  AND2X1 U651 ( .A(n89), .B(n835), .Y(n635) );
  INVX1 U652 ( .A(n635), .Y(n636) );
  AND2X1 U653 ( .A(n81), .B(n835), .Y(n637) );
  INVX1 U654 ( .A(n637), .Y(n638) );
  AND2X1 U655 ( .A(n73), .B(n835), .Y(n639) );
  INVX1 U656 ( .A(n639), .Y(n640) );
  AND2X1 U657 ( .A(n65), .B(n835), .Y(n641) );
  INVX1 U658 ( .A(n641), .Y(n642) );
  MUX2X1 U659 ( .B(n729), .A(n728), .S(n827), .Y(n727) );
  INVX1 U660 ( .A(n804), .Y(n643) );
  INVX1 U661 ( .A(N10), .Y(n644) );
  MUX2X1 U662 ( .B(\mem<11><4> ), .A(\mem<10><4> ), .S(n811), .Y(n788) );
  INVX1 U663 ( .A(N10), .Y(n826) );
  INVX1 U664 ( .A(n826), .Y(n825) );
  INVX2 U665 ( .A(n825), .Y(n645) );
  INVX8 U666 ( .A(n810), .Y(n811) );
  INVX1 U667 ( .A(n811), .Y(n814) );
  INVX8 U668 ( .A(n645), .Y(n815) );
  INVX1 U669 ( .A(n802), .Y(N17) );
  MUX2X1 U670 ( .B(n732), .A(n731), .S(n805), .Y(n730) );
  NAND2X1 U671 ( .A(\mem<30><2> ), .B(n811), .Y(n646) );
  NAND2X1 U672 ( .A(\mem<31><2> ), .B(n812), .Y(n647) );
  MUX2X1 U673 ( .B(\mem<9><0> ), .A(\mem<8><0> ), .S(n811), .Y(n669) );
  BUFX2 U674 ( .A(write), .Y(n648) );
  INVX1 U675 ( .A(n798), .Y(N21) );
  MUX2X1 U676 ( .B(n710), .A(n712), .S(n829), .Y(n723) );
  MUX2X1 U677 ( .B(\mem<1><3> ), .A(\mem<0><3> ), .S(n818), .Y(n763) );
  MUX2X1 U678 ( .B(\mem<9><3> ), .A(\mem<8><3> ), .S(n811), .Y(n757) );
  INVX1 U679 ( .A(n825), .Y(n649) );
  MUX2X1 U680 ( .B(\mem<11><0> ), .A(\mem<10><0> ), .S(n811), .Y(n670) );
  MUX2X1 U681 ( .B(\mem<11><1> ), .A(\mem<10><1> ), .S(n645), .Y(n700) );
  MUX2X1 U682 ( .B(\mem<3><0> ), .A(\mem<2><0> ), .S(n818), .Y(n676) );
  MUX2X1 U683 ( .B(\mem<3><3> ), .A(\mem<2><3> ), .S(n811), .Y(n764) );
  MUX2X1 U684 ( .B(\mem<11><2> ), .A(\mem<10><2> ), .S(n818), .Y(n729) );
  MUX2X1 U685 ( .B(\mem<11><3> ), .A(\mem<10><3> ), .S(n811), .Y(n758) );
  MUX2X1 U686 ( .B(n651), .A(n652), .S(n809), .Y(n650) );
  MUX2X1 U687 ( .B(n654), .A(n655), .S(n809), .Y(n653) );
  MUX2X1 U688 ( .B(n657), .A(n658), .S(n809), .Y(n656) );
  MUX2X1 U689 ( .B(n660), .A(n661), .S(n809), .Y(n659) );
  MUX2X1 U690 ( .B(n663), .A(n664), .S(N13), .Y(n662) );
  MUX2X1 U691 ( .B(n666), .A(n667), .S(n809), .Y(n665) );
  MUX2X1 U692 ( .B(n669), .A(n670), .S(n809), .Y(n668) );
  MUX2X1 U693 ( .B(n672), .A(n673), .S(n809), .Y(n671) );
  MUX2X1 U694 ( .B(n675), .A(n676), .S(n809), .Y(n674) );
  MUX2X1 U695 ( .B(n678), .A(n679), .S(N13), .Y(n677) );
  MUX2X1 U696 ( .B(n681), .A(n682), .S(n809), .Y(n680) );
  MUX2X1 U697 ( .B(n684), .A(n685), .S(n809), .Y(n683) );
  MUX2X1 U698 ( .B(n687), .A(n688), .S(n809), .Y(n686) );
  MUX2X1 U699 ( .B(n690), .A(n691), .S(n809), .Y(n689) );
  MUX2X1 U700 ( .B(n693), .A(n694), .S(N13), .Y(n692) );
  MUX2X1 U701 ( .B(n696), .A(n697), .S(n806), .Y(n695) );
  MUX2X1 U702 ( .B(n699), .A(n700), .S(n808), .Y(n698) );
  MUX2X1 U703 ( .B(n702), .A(n703), .S(n807), .Y(n701) );
  MUX2X1 U704 ( .B(n705), .A(n706), .S(n808), .Y(n704) );
  MUX2X1 U705 ( .B(n708), .A(n709), .S(N13), .Y(n707) );
  MUX2X1 U706 ( .B(n711), .A(n3), .S(n806), .Y(n710) );
  MUX2X1 U707 ( .B(n713), .A(n714), .S(n806), .Y(n712) );
  MUX2X1 U708 ( .B(n716), .A(n717), .S(n806), .Y(n715) );
  MUX2X1 U709 ( .B(n719), .A(n720), .S(n807), .Y(n718) );
  MUX2X1 U710 ( .B(n722), .A(n723), .S(N13), .Y(n721) );
  MUX2X1 U711 ( .B(n725), .A(n726), .S(n806), .Y(n724) );
  MUX2X1 U712 ( .B(n734), .A(n735), .S(n808), .Y(n733) );
  MUX2X1 U713 ( .B(n737), .A(n2), .S(N13), .Y(n736) );
  MUX2X1 U714 ( .B(n739), .A(n740), .S(n807), .Y(n738) );
  MUX2X1 U715 ( .B(n742), .A(n743), .S(n807), .Y(n741) );
  MUX2X1 U716 ( .B(n745), .A(n746), .S(n807), .Y(n744) );
  MUX2X1 U717 ( .B(n748), .A(n749), .S(n807), .Y(n747) );
  MUX2X1 U718 ( .B(n751), .A(n752), .S(N13), .Y(n750) );
  MUX2X1 U719 ( .B(n754), .A(n755), .S(n807), .Y(n753) );
  MUX2X1 U720 ( .B(n757), .A(n758), .S(n808), .Y(n756) );
  MUX2X1 U721 ( .B(n760), .A(n761), .S(n806), .Y(n759) );
  MUX2X1 U722 ( .B(n763), .A(n764), .S(n808), .Y(n762) );
  MUX2X1 U723 ( .B(n766), .A(n767), .S(N13), .Y(n765) );
  MUX2X1 U724 ( .B(n769), .A(n770), .S(n806), .Y(n768) );
  MUX2X1 U725 ( .B(n772), .A(n773), .S(n806), .Y(n771) );
  MUX2X1 U726 ( .B(n775), .A(n776), .S(n807), .Y(n774) );
  MUX2X1 U727 ( .B(n778), .A(n779), .S(n806), .Y(n777) );
  MUX2X1 U728 ( .B(n781), .A(n782), .S(N13), .Y(n780) );
  MUX2X1 U729 ( .B(n784), .A(n785), .S(n807), .Y(n783) );
  MUX2X1 U730 ( .B(n787), .A(n788), .S(n807), .Y(n786) );
  MUX2X1 U731 ( .B(n790), .A(n791), .S(n806), .Y(n789) );
  MUX2X1 U732 ( .B(n793), .A(n794), .S(n807), .Y(n792) );
  MUX2X1 U733 ( .B(n796), .A(n797), .S(N13), .Y(n795) );
  MUX2X1 U734 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n817), .Y(n652) );
  MUX2X1 U735 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n817), .Y(n651) );
  MUX2X1 U736 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n817), .Y(n655) );
  MUX2X1 U737 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n817), .Y(n654) );
  MUX2X1 U738 ( .B(n653), .A(n650), .S(n804), .Y(n664) );
  MUX2X1 U739 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n817), .Y(n658) );
  MUX2X1 U740 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n817), .Y(n657) );
  MUX2X1 U741 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n817), .Y(n661) );
  MUX2X1 U742 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n817), .Y(n660) );
  MUX2X1 U743 ( .B(n659), .A(n656), .S(n804), .Y(n663) );
  MUX2X1 U744 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n817), .Y(n667) );
  MUX2X1 U745 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n817), .Y(n666) );
  MUX2X1 U746 ( .B(n668), .A(n665), .S(n804), .Y(n679) );
  MUX2X1 U747 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n815), .Y(n673) );
  MUX2X1 U748 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n816), .Y(n672) );
  MUX2X1 U749 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n814), .Y(n675) );
  MUX2X1 U750 ( .B(n674), .A(n671), .S(n804), .Y(n678) );
  MUX2X1 U751 ( .B(n677), .A(n662), .S(N14), .Y(n798) );
  MUX2X1 U752 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n816), .Y(n682) );
  MUX2X1 U753 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n816), .Y(n681) );
  MUX2X1 U754 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n815), .Y(n685) );
  MUX2X1 U755 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n816), .Y(n684) );
  MUX2X1 U756 ( .B(n683), .A(n680), .S(n804), .Y(n694) );
  MUX2X1 U757 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n816), .Y(n688) );
  MUX2X1 U758 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n816), .Y(n687) );
  MUX2X1 U759 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n816), .Y(n691) );
  MUX2X1 U760 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n816), .Y(n690) );
  MUX2X1 U761 ( .B(n689), .A(n686), .S(n804), .Y(n693) );
  MUX2X1 U762 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n815), .Y(n697) );
  MUX2X1 U763 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n816), .Y(n696) );
  MUX2X1 U764 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n813), .Y(n699) );
  MUX2X1 U765 ( .B(n698), .A(n695), .S(n804), .Y(n709) );
  MUX2X1 U766 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n816), .Y(n703) );
  MUX2X1 U767 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n816), .Y(n702) );
  MUX2X1 U768 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n816), .Y(n706) );
  MUX2X1 U769 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n816), .Y(n705) );
  MUX2X1 U770 ( .B(n704), .A(n701), .S(n804), .Y(n708) );
  MUX2X1 U771 ( .B(n707), .A(n692), .S(N14), .Y(n799) );
  MUX2X1 U772 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n815), .Y(n711) );
  MUX2X1 U773 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n816), .Y(n714) );
  MUX2X1 U774 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n816), .Y(n713) );
  MUX2X1 U775 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n816), .Y(n717) );
  MUX2X1 U776 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n816), .Y(n716) );
  MUX2X1 U777 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n815), .Y(n720) );
  MUX2X1 U778 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n816), .Y(n719) );
  MUX2X1 U779 ( .B(n718), .A(n715), .S(n804), .Y(n722) );
  MUX2X1 U780 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n810), .Y(n726) );
  MUX2X1 U781 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n815), .Y(n725) );
  MUX2X1 U782 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n810), .Y(n728) );
  MUX2X1 U783 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n812), .Y(n732) );
  MUX2X1 U784 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n815), .Y(n731) );
  MUX2X1 U785 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n817), .Y(n735) );
  MUX2X1 U786 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n816), .Y(n734) );
  MUX2X1 U787 ( .B(n733), .A(n730), .S(n804), .Y(n737) );
  MUX2X1 U788 ( .B(n736), .A(n721), .S(N14), .Y(n800) );
  MUX2X1 U789 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n813), .Y(n740) );
  MUX2X1 U790 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n812), .Y(n739) );
  MUX2X1 U791 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n815), .Y(n743) );
  MUX2X1 U792 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n814), .Y(n742) );
  MUX2X1 U793 ( .B(n741), .A(n738), .S(n803), .Y(n752) );
  MUX2X1 U794 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n813), .Y(n746) );
  MUX2X1 U795 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n813), .Y(n745) );
  MUX2X1 U796 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n815), .Y(n749) );
  MUX2X1 U797 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n812), .Y(n748) );
  MUX2X1 U798 ( .B(n747), .A(n744), .S(n803), .Y(n751) );
  MUX2X1 U799 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n815), .Y(n755) );
  MUX2X1 U800 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n815), .Y(n754) );
  MUX2X1 U801 ( .B(n756), .A(n753), .S(n803), .Y(n767) );
  MUX2X1 U802 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n815), .Y(n761) );
  MUX2X1 U803 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n813), .Y(n760) );
  MUX2X1 U804 ( .B(n762), .A(n759), .S(n803), .Y(n766) );
  MUX2X1 U805 ( .B(n765), .A(n750), .S(N14), .Y(n801) );
  MUX2X1 U806 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n812), .Y(n770) );
  MUX2X1 U807 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n812), .Y(n769) );
  MUX2X1 U808 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n813), .Y(n773) );
  MUX2X1 U809 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n813), .Y(n772) );
  MUX2X1 U810 ( .B(n771), .A(n768), .S(n803), .Y(n782) );
  MUX2X1 U811 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n813), .Y(n776) );
  MUX2X1 U812 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n813), .Y(n775) );
  MUX2X1 U813 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n812), .Y(n779) );
  MUX2X1 U814 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n813), .Y(n778) );
  MUX2X1 U815 ( .B(n777), .A(n774), .S(n803), .Y(n781) );
  MUX2X1 U816 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n812), .Y(n785) );
  MUX2X1 U817 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n813), .Y(n784) );
  MUX2X1 U818 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n812), .Y(n787) );
  MUX2X1 U819 ( .B(n786), .A(n783), .S(n803), .Y(n797) );
  MUX2X1 U820 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n812), .Y(n791) );
  MUX2X1 U821 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n812), .Y(n790) );
  MUX2X1 U822 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n813), .Y(n794) );
  MUX2X1 U823 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n812), .Y(n793) );
  MUX2X1 U824 ( .B(n792), .A(n789), .S(n803), .Y(n796) );
  MUX2X1 U825 ( .B(n795), .A(n780), .S(N14), .Y(n802) );
  INVX8 U826 ( .A(n829), .Y(n803) );
  INVX8 U827 ( .A(n829), .Y(n804) );
  INVX8 U828 ( .A(N11), .Y(n805) );
  INVX8 U829 ( .A(n805), .Y(n806) );
  INVX8 U830 ( .A(n805), .Y(n807) );
  INVX8 U831 ( .A(n805), .Y(n808) );
  INVX8 U832 ( .A(n805), .Y(n809) );
  INVX8 U833 ( .A(n811), .Y(n812) );
  INVX8 U834 ( .A(n811), .Y(n813) );
  INVX8 U835 ( .A(n645), .Y(n816) );
  INVX8 U836 ( .A(n811), .Y(n817) );
  INVX1 U837 ( .A(n800), .Y(N19) );
  INVX1 U838 ( .A(n801), .Y(N18) );
  INVX1 U839 ( .A(n799), .Y(N20) );
  BUFX2 U840 ( .A(n649), .Y(n818) );
  INVX8 U841 ( .A(N12), .Y(n829) );
  AND2X2 U842 ( .A(n502), .B(N21), .Y(\data_out<0> ) );
  AND2X2 U843 ( .A(N20), .B(n503), .Y(\data_out<1> ) );
  AND2X2 U844 ( .A(n502), .B(N19), .Y(\data_out<2> ) );
  AND2X2 U845 ( .A(n505), .B(N18), .Y(\data_out<3> ) );
  AND2X2 U846 ( .A(N17), .B(n503), .Y(\data_out<4> ) );
endmodule


module memc_Size1_1 ( .data_out(\data_out<0> ), .addr({\addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
    .data_in(\data_in<0> ), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<0> , write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><0> , \mem<1><0> , \mem<2><0> ,
         \mem<3><0> , \mem<4><0> , \mem<5><0> , \mem<6><0> , \mem<7><0> ,
         \mem<8><0> , \mem<9><0> , \mem<10><0> , \mem<11><0> , \mem<12><0> ,
         \mem<13><0> , \mem<14><0> , \mem<15><0> , \mem<16><0> , \mem<17><0> ,
         \mem<18><0> , \mem<19><0> , \mem<20><0> , \mem<21><0> , \mem<22><0> ,
         \mem<23><0> , \mem<24><0> , \mem<25><0> , \mem<26><0> , \mem<27><0> ,
         \mem<28><0> , \mem<29><0> , \mem<30><0> , \mem<31><0> , N17, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><0>  ( .D(n92), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n91), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n90), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n89), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n88), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n87), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n86), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n85), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n84), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n83), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n82), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n81), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n80), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n79), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n78), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n77), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n76), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n75), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n74), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n73), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n72), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n71), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n70), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n69), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n68), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n67), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n66), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n65), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n64), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n63), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n62), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n61), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X1 U2 ( .A(n56), .B(n154), .Y(n59) );
  INVX1 U3 ( .A(n158), .Y(n149) );
  INVX1 U4 ( .A(n148), .Y(N17) );
  OR2X1 U5 ( .A(n60), .B(\addr<5> ), .Y(n96) );
  INVX1 U6 ( .A(N12), .Y(n160) );
  INVX1 U7 ( .A(n98), .Y(n195) );
  INVX1 U8 ( .A(n99), .Y(n198) );
  INVX1 U9 ( .A(n100), .Y(n201) );
  INVX1 U10 ( .A(n101), .Y(n204) );
  INVX1 U11 ( .A(n155), .Y(n150) );
  INVX2 U12 ( .A(n112), .Y(n113) );
  INVX2 U13 ( .A(n114), .Y(n115) );
  INVX1 U14 ( .A(n192), .Y(n153) );
  BUFX2 U15 ( .A(write), .Y(n1) );
  OR2X2 U16 ( .A(write), .B(n94), .Y(n2) );
  INVX1 U17 ( .A(n2), .Y(\data_out<0> ) );
  AND2X2 U18 ( .A(\data_in<0> ), .B(n112), .Y(n4) );
  AND2X2 U19 ( .A(\data_in<0> ), .B(n114), .Y(n5) );
  AND2X2 U20 ( .A(n108), .B(n54), .Y(n6) );
  INVX1 U21 ( .A(n6), .Y(n7) );
  AND2X2 U22 ( .A(n105), .B(n54), .Y(n8) );
  INVX1 U23 ( .A(n8), .Y(n9) );
  AND2X2 U24 ( .A(n195), .B(n54), .Y(n10) );
  INVX1 U25 ( .A(n10), .Y(n11) );
  AND2X2 U26 ( .A(n198), .B(n54), .Y(n12) );
  INVX1 U27 ( .A(n12), .Y(n13) );
  AND2X2 U28 ( .A(n201), .B(n54), .Y(n14) );
  INVX1 U29 ( .A(n14), .Y(n15) );
  AND2X2 U30 ( .A(n204), .B(n54), .Y(n16) );
  INVX1 U31 ( .A(n16), .Y(n17) );
  AND2X2 U32 ( .A(n102), .B(n54), .Y(n18) );
  INVX1 U33 ( .A(n18), .Y(n19) );
  AND2X2 U34 ( .A(n107), .B(n54), .Y(n20) );
  INVX1 U35 ( .A(n20), .Y(n21) );
  AND2X2 U36 ( .A(n108), .B(n4), .Y(n22) );
  INVX1 U37 ( .A(n22), .Y(n23) );
  AND2X2 U38 ( .A(n105), .B(n4), .Y(n24) );
  INVX1 U39 ( .A(n24), .Y(n25) );
  AND2X2 U40 ( .A(n195), .B(n4), .Y(n26) );
  INVX1 U41 ( .A(n26), .Y(n27) );
  AND2X2 U42 ( .A(n198), .B(n4), .Y(n28) );
  INVX1 U43 ( .A(n28), .Y(n29) );
  AND2X2 U44 ( .A(n201), .B(n4), .Y(n30) );
  INVX1 U45 ( .A(n30), .Y(n31) );
  AND2X2 U46 ( .A(n204), .B(n4), .Y(n32) );
  INVX1 U47 ( .A(n32), .Y(n33) );
  AND2X2 U48 ( .A(n102), .B(n4), .Y(n34) );
  INVX1 U49 ( .A(n34), .Y(n35) );
  AND2X2 U50 ( .A(n107), .B(n4), .Y(n36) );
  INVX1 U51 ( .A(n36), .Y(n37) );
  AND2X2 U52 ( .A(n108), .B(n5), .Y(n38) );
  INVX1 U53 ( .A(n38), .Y(n39) );
  AND2X2 U54 ( .A(n105), .B(n5), .Y(n40) );
  INVX1 U55 ( .A(n40), .Y(n41) );
  AND2X2 U56 ( .A(n195), .B(n5), .Y(n42) );
  INVX1 U57 ( .A(n42), .Y(n43) );
  AND2X2 U58 ( .A(n198), .B(n5), .Y(n44) );
  INVX1 U59 ( .A(n44), .Y(n45) );
  AND2X2 U60 ( .A(n201), .B(n5), .Y(n46) );
  INVX1 U61 ( .A(n46), .Y(n47) );
  AND2X2 U62 ( .A(n204), .B(n5), .Y(n48) );
  INVX1 U63 ( .A(n48), .Y(n49) );
  AND2X2 U64 ( .A(n102), .B(n5), .Y(n50) );
  INVX1 U65 ( .A(n50), .Y(n51) );
  AND2X2 U66 ( .A(n107), .B(n5), .Y(n52) );
  INVX1 U67 ( .A(n52), .Y(n53) );
  INVX1 U68 ( .A(n160), .Y(n159) );
  INVX1 U69 ( .A(n158), .Y(n157) );
  INVX1 U70 ( .A(n156), .Y(n155) );
  AND2X2 U71 ( .A(\data_in<0> ), .B(n116), .Y(n54) );
  OR2X1 U72 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n55) );
  INVX1 U73 ( .A(n55), .Y(n56) );
  OR2X1 U74 ( .A(n157), .B(n159), .Y(n57) );
  INVX1 U75 ( .A(n57), .Y(n58) );
  INVX1 U76 ( .A(n59), .Y(n60) );
  AND2X1 U77 ( .A(N17), .B(n154), .Y(n93) );
  INVX1 U78 ( .A(n93), .Y(n94) );
  AND2X1 U79 ( .A(n159), .B(n157), .Y(n95) );
  INVX1 U80 ( .A(n96), .Y(n97) );
  BUFX2 U81 ( .A(n196), .Y(n98) );
  BUFX2 U82 ( .A(n199), .Y(n99) );
  BUFX2 U83 ( .A(n202), .Y(n100) );
  BUFX2 U84 ( .A(n205), .Y(n101) );
  INVX1 U85 ( .A(n103), .Y(n102) );
  BUFX2 U86 ( .A(n207), .Y(n103) );
  INVX1 U87 ( .A(n105), .Y(n104) );
  AND2X1 U88 ( .A(n156), .B(n95), .Y(n105) );
  INVX1 U89 ( .A(n107), .Y(n106) );
  AND2X2 U90 ( .A(n156), .B(n58), .Y(n107) );
  AND2X1 U91 ( .A(n155), .B(n95), .Y(n108) );
  INVX1 U92 ( .A(n108), .Y(n109) );
  AND2X2 U93 ( .A(\data_in<0> ), .B(n152), .Y(n110) );
  INVX1 U94 ( .A(n110), .Y(n111) );
  INVX1 U95 ( .A(n190), .Y(n112) );
  INVX1 U96 ( .A(n209), .Y(n114) );
  INVX1 U97 ( .A(n181), .Y(n116) );
  INVX1 U98 ( .A(n116), .Y(n117) );
  MUX2X1 U99 ( .B(n119), .A(n120), .S(n149), .Y(n118) );
  MUX2X1 U100 ( .B(n122), .A(n123), .S(n149), .Y(n121) );
  MUX2X1 U101 ( .B(n125), .A(n126), .S(n149), .Y(n124) );
  MUX2X1 U102 ( .B(n128), .A(n129), .S(n149), .Y(n127) );
  MUX2X1 U103 ( .B(n131), .A(n132), .S(n161), .Y(n130) );
  MUX2X1 U104 ( .B(n134), .A(n135), .S(n149), .Y(n133) );
  MUX2X1 U105 ( .B(n137), .A(n138), .S(n149), .Y(n136) );
  MUX2X1 U106 ( .B(n140), .A(n141), .S(n149), .Y(n139) );
  MUX2X1 U107 ( .B(n143), .A(n144), .S(n149), .Y(n142) );
  MUX2X1 U108 ( .B(n146), .A(n147), .S(n161), .Y(n145) );
  MUX2X1 U109 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n151), .Y(n120) );
  MUX2X1 U110 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n151), .Y(n119) );
  MUX2X1 U111 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n151), .Y(n123) );
  MUX2X1 U112 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n151), .Y(n122) );
  MUX2X1 U113 ( .B(n121), .A(n118), .S(n159), .Y(n132) );
  MUX2X1 U114 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n151), .Y(n126) );
  MUX2X1 U115 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n151), .Y(n125) );
  MUX2X1 U116 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n151), .Y(n129) );
  MUX2X1 U117 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n151), .Y(n128) );
  MUX2X1 U118 ( .B(n127), .A(n124), .S(n159), .Y(n131) );
  MUX2X1 U119 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n151), .Y(n135) );
  MUX2X1 U120 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n151), .Y(n134) );
  MUX2X1 U121 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n151), .Y(n138) );
  MUX2X1 U122 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n151), .Y(n137) );
  MUX2X1 U123 ( .B(n136), .A(n133), .S(n159), .Y(n147) );
  MUX2X1 U124 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n151), .Y(n141) );
  MUX2X1 U125 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n151), .Y(n140) );
  MUX2X1 U126 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n151), .Y(n144) );
  MUX2X1 U127 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n151), .Y(n143) );
  MUX2X1 U128 ( .B(n142), .A(n139), .S(n159), .Y(n146) );
  MUX2X1 U129 ( .B(n145), .A(n130), .S(n163), .Y(n148) );
  INVX8 U130 ( .A(n150), .Y(n151) );
  NOR3X1 U131 ( .A(n164), .B(n162), .C(n153), .Y(n152) );
  INVX4 U132 ( .A(n152), .Y(n172) );
  INVX1 U133 ( .A(n164), .Y(n163) );
  INVX1 U134 ( .A(N14), .Y(n164) );
  INVX1 U135 ( .A(n162), .Y(n161) );
  INVX1 U136 ( .A(N13), .Y(n162) );
  INVX1 U137 ( .A(N11), .Y(n158) );
  AND2X2 U138 ( .A(n1), .B(n97), .Y(n192) );
  INVX1 U139 ( .A(rst), .Y(n154) );
  INVX1 U140 ( .A(N10), .Y(n156) );
  OAI21X1 U141 ( .A(n172), .B(n109), .C(\mem<31><0> ), .Y(n165) );
  OAI21X1 U142 ( .A(n111), .B(n109), .C(n165), .Y(n61) );
  OAI21X1 U143 ( .A(n104), .B(n172), .C(\mem<30><0> ), .Y(n166) );
  OAI21X1 U144 ( .A(n104), .B(n111), .C(n166), .Y(n62) );
  NAND3X1 U145 ( .A(n155), .B(n159), .C(n158), .Y(n196) );
  OAI21X1 U146 ( .A(n98), .B(n172), .C(\mem<29><0> ), .Y(n167) );
  OAI21X1 U147 ( .A(n98), .B(n111), .C(n167), .Y(n63) );
  NAND3X1 U148 ( .A(n159), .B(n158), .C(n156), .Y(n199) );
  OAI21X1 U149 ( .A(n99), .B(n172), .C(\mem<28><0> ), .Y(n168) );
  OAI21X1 U150 ( .A(n99), .B(n111), .C(n168), .Y(n64) );
  NAND3X1 U151 ( .A(n155), .B(n157), .C(n160), .Y(n202) );
  OAI21X1 U152 ( .A(n100), .B(n172), .C(\mem<27><0> ), .Y(n169) );
  OAI21X1 U153 ( .A(n100), .B(n111), .C(n169), .Y(n65) );
  NAND3X1 U154 ( .A(n160), .B(n157), .C(n156), .Y(n205) );
  OAI21X1 U155 ( .A(n101), .B(n172), .C(\mem<26><0> ), .Y(n170) );
  OAI21X1 U156 ( .A(n101), .B(n111), .C(n170), .Y(n66) );
  NAND3X1 U157 ( .A(n155), .B(n160), .C(n158), .Y(n207) );
  OAI21X1 U158 ( .A(n103), .B(n172), .C(\mem<25><0> ), .Y(n171) );
  OAI21X1 U159 ( .A(n103), .B(n111), .C(n171), .Y(n67) );
  OAI21X1 U160 ( .A(n106), .B(n172), .C(\mem<24><0> ), .Y(n173) );
  OAI21X1 U161 ( .A(n106), .B(n111), .C(n173), .Y(n68) );
  NAND3X1 U162 ( .A(n163), .B(n192), .C(n162), .Y(n181) );
  OAI21X1 U163 ( .A(n117), .B(n109), .C(\mem<23><0> ), .Y(n174) );
  NAND2X1 U164 ( .A(n7), .B(n174), .Y(n69) );
  OAI21X1 U165 ( .A(n117), .B(n104), .C(\mem<22><0> ), .Y(n175) );
  NAND2X1 U166 ( .A(n9), .B(n175), .Y(n70) );
  OAI21X1 U167 ( .A(n117), .B(n98), .C(\mem<21><0> ), .Y(n176) );
  NAND2X1 U168 ( .A(n11), .B(n176), .Y(n71) );
  OAI21X1 U169 ( .A(n117), .B(n99), .C(\mem<20><0> ), .Y(n177) );
  NAND2X1 U170 ( .A(n13), .B(n177), .Y(n72) );
  OAI21X1 U171 ( .A(n117), .B(n100), .C(\mem<19><0> ), .Y(n178) );
  NAND2X1 U172 ( .A(n15), .B(n178), .Y(n73) );
  OAI21X1 U173 ( .A(n117), .B(n101), .C(\mem<18><0> ), .Y(n179) );
  NAND2X1 U174 ( .A(n17), .B(n179), .Y(n74) );
  OAI21X1 U175 ( .A(n117), .B(n103), .C(\mem<17><0> ), .Y(n180) );
  NAND2X1 U176 ( .A(n19), .B(n180), .Y(n75) );
  OAI21X1 U177 ( .A(n117), .B(n106), .C(\mem<16><0> ), .Y(n182) );
  NAND2X1 U178 ( .A(n21), .B(n182), .Y(n76) );
  NAND3X1 U179 ( .A(n161), .B(n192), .C(n164), .Y(n190) );
  OAI21X1 U180 ( .A(n113), .B(n109), .C(\mem<15><0> ), .Y(n183) );
  NAND2X1 U181 ( .A(n23), .B(n183), .Y(n77) );
  OAI21X1 U182 ( .A(n113), .B(n104), .C(\mem<14><0> ), .Y(n184) );
  NAND2X1 U183 ( .A(n25), .B(n184), .Y(n78) );
  OAI21X1 U184 ( .A(n113), .B(n98), .C(\mem<13><0> ), .Y(n185) );
  NAND2X1 U185 ( .A(n27), .B(n185), .Y(n79) );
  OAI21X1 U186 ( .A(n113), .B(n99), .C(\mem<12><0> ), .Y(n186) );
  NAND2X1 U187 ( .A(n29), .B(n186), .Y(n80) );
  OAI21X1 U188 ( .A(n113), .B(n100), .C(\mem<11><0> ), .Y(n187) );
  NAND2X1 U189 ( .A(n31), .B(n187), .Y(n81) );
  OAI21X1 U190 ( .A(n113), .B(n101), .C(\mem<10><0> ), .Y(n188) );
  NAND2X1 U191 ( .A(n33), .B(n188), .Y(n82) );
  OAI21X1 U192 ( .A(n113), .B(n103), .C(\mem<9><0> ), .Y(n189) );
  NAND2X1 U193 ( .A(n35), .B(n189), .Y(n83) );
  OAI21X1 U194 ( .A(n113), .B(n106), .C(\mem<8><0> ), .Y(n191) );
  NAND2X1 U195 ( .A(n37), .B(n191), .Y(n84) );
  NAND3X1 U196 ( .A(n162), .B(n192), .C(n164), .Y(n209) );
  OAI21X1 U197 ( .A(n115), .B(n109), .C(\mem<7><0> ), .Y(n193) );
  NAND2X1 U198 ( .A(n39), .B(n193), .Y(n85) );
  OAI21X1 U199 ( .A(n115), .B(n104), .C(\mem<6><0> ), .Y(n194) );
  NAND2X1 U200 ( .A(n41), .B(n194), .Y(n86) );
  OAI21X1 U201 ( .A(n115), .B(n98), .C(\mem<5><0> ), .Y(n197) );
  NAND2X1 U202 ( .A(n43), .B(n197), .Y(n87) );
  OAI21X1 U203 ( .A(n115), .B(n99), .C(\mem<4><0> ), .Y(n200) );
  NAND2X1 U204 ( .A(n45), .B(n200), .Y(n88) );
  OAI21X1 U205 ( .A(n115), .B(n100), .C(\mem<3><0> ), .Y(n203) );
  NAND2X1 U206 ( .A(n47), .B(n203), .Y(n89) );
  OAI21X1 U207 ( .A(n115), .B(n101), .C(\mem<2><0> ), .Y(n206) );
  NAND2X1 U208 ( .A(n49), .B(n206), .Y(n90) );
  OAI21X1 U209 ( .A(n115), .B(n103), .C(\mem<1><0> ), .Y(n208) );
  NAND2X1 U210 ( .A(n51), .B(n208), .Y(n91) );
  OAI21X1 U211 ( .A(n115), .B(n106), .C(\mem<0><0> ), .Y(n210) );
  NAND2X1 U212 ( .A(n53), .B(n210), .Y(n92) );
endmodule


module memv_1 ( data_out, .addr({\addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), data_in, write, clk, rst, 
        createdump, .file_id({\file_id<4> , \file_id<3> , \file_id<2> , 
        \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , data_in, write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output data_out;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \mem<0> , \mem<1> , \mem<2> ,
         \mem<3> , \mem<4> , \mem<5> , \mem<6> , \mem<7> , \mem<8> , \mem<9> ,
         \mem<10> , \mem<11> , \mem<12> , \mem<13> , \mem<14> , \mem<15> ,
         \mem<16> , \mem<17> , \mem<18> , \mem<19> , \mem<20> , \mem<21> ,
         \mem<22> , \mem<23> , \mem<24> , \mem<25> , \mem<26> , \mem<27> ,
         \mem<28> , \mem<29> , \mem<30> , \mem<31> , \mem<32> , \mem<33> ,
         \mem<34> , \mem<35> , \mem<36> , \mem<37> , \mem<38> , \mem<39> ,
         \mem<40> , \mem<41> , \mem<42> , \mem<43> , \mem<44> , \mem<45> ,
         \mem<46> , \mem<47> , \mem<48> , \mem<49> , \mem<50> , \mem<51> ,
         \mem<52> , \mem<53> , \mem<54> , \mem<55> , \mem<56> , \mem<57> ,
         \mem<58> , \mem<59> , \mem<60> , \mem<61> , \mem<62> , \mem<63> ,
         \mem<64> , \mem<65> , \mem<66> , \mem<67> , \mem<68> , \mem<69> ,
         \mem<70> , \mem<71> , \mem<72> , \mem<73> , \mem<74> , \mem<75> ,
         \mem<76> , \mem<77> , \mem<78> , \mem<79> , \mem<80> , \mem<81> ,
         \mem<82> , \mem<83> , \mem<84> , \mem<85> , \mem<86> , \mem<87> ,
         \mem<88> , \mem<89> , \mem<90> , \mem<91> , \mem<92> , \mem<93> ,
         \mem<94> , \mem<95> , \mem<96> , \mem<97> , \mem<98> , \mem<99> ,
         \mem<100> , \mem<101> , \mem<102> , \mem<103> , \mem<104> ,
         \mem<105> , \mem<106> , \mem<107> , \mem<108> , \mem<109> ,
         \mem<110> , \mem<111> , \mem<112> , \mem<113> , \mem<114> ,
         \mem<115> , \mem<116> , \mem<117> , \mem<118> , \mem<119> ,
         \mem<120> , \mem<121> , \mem<122> , \mem<123> , \mem<124> ,
         \mem<125> , \mem<126> , \mem<127> , \mem<128> , \mem<129> ,
         \mem<130> , \mem<131> , \mem<132> , \mem<133> , \mem<134> ,
         \mem<135> , \mem<136> , \mem<137> , \mem<138> , \mem<139> ,
         \mem<140> , \mem<141> , \mem<142> , \mem<143> , \mem<144> ,
         \mem<145> , \mem<146> , \mem<147> , \mem<148> , \mem<149> ,
         \mem<150> , \mem<151> , \mem<152> , \mem<153> , \mem<154> ,
         \mem<155> , \mem<156> , \mem<157> , \mem<158> , \mem<159> ,
         \mem<160> , \mem<161> , \mem<162> , \mem<163> , \mem<164> ,
         \mem<165> , \mem<166> , \mem<167> , \mem<168> , \mem<169> ,
         \mem<170> , \mem<171> , \mem<172> , \mem<173> , \mem<174> ,
         \mem<175> , \mem<176> , \mem<177> , \mem<178> , \mem<179> ,
         \mem<180> , \mem<181> , \mem<182> , \mem<183> , \mem<184> ,
         \mem<185> , \mem<186> , \mem<187> , \mem<188> , \mem<189> ,
         \mem<190> , \mem<191> , \mem<192> , \mem<193> , \mem<194> ,
         \mem<195> , \mem<196> , \mem<197> , \mem<198> , \mem<199> ,
         \mem<200> , \mem<201> , \mem<202> , \mem<203> , \mem<204> ,
         \mem<205> , \mem<206> , \mem<207> , \mem<208> , \mem<209> ,
         \mem<210> , \mem<211> , \mem<212> , \mem<213> , \mem<214> ,
         \mem<215> , \mem<216> , \mem<217> , \mem<218> , \mem<219> ,
         \mem<220> , \mem<221> , \mem<222> , \mem<223> , \mem<224> ,
         \mem<225> , \mem<226> , \mem<227> , \mem<228> , \mem<229> ,
         \mem<230> , \mem<231> , \mem<232> , \mem<233> , \mem<234> ,
         \mem<235> , \mem<236> , \mem<237> , \mem<238> , \mem<239> ,
         \mem<240> , \mem<241> , \mem<242> , \mem<243> , \mem<244> ,
         \mem<245> , \mem<246> , \mem<247> , \mem<248> , \mem<249> ,
         \mem<250> , \mem<251> , \mem<252> , \mem<253> , \mem<254> ,
         \mem<255> , N28, n42, n46, n49, n52, n55, n58, n61, n64, n67, n70,
         n73, n76, n79, n82, n85, n88, n90, n91, n92, n94, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n113, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n132, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n151, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n170, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n188, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n206, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n224,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n243, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n261, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n279, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n297, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n316, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n334, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n352, n355, n356, n357, n358, n359, n361, n363, n364, n365,
         n366, n367, n368, n370, n371, n372, n373, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n43, n44, n45, n47, n48, n50, n51, n53, n54, n56, n57, n59, n60, n62,
         n63, n65, n66, n68, n69, n71, n72, n74, n75, n77, n78, n80, n81, n83,
         n84, n86, n87, n89, n93, n95, n112, n114, n130, n131, n133, n149,
         n150, n152, n169, n171, n187, n189, n205, n207, n223, n225, n241,
         n242, n244, n260, n262, n278, n280, n296, n298, n314, n315, n317,
         n333, n335, n351, n353, n354, n360, n362, n369, n374, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988;
  assign N18 = \addr<0> ;
  assign N19 = \addr<1> ;
  assign N20 = \addr<2> ;
  assign N21 = \addr<3> ;
  assign N22 = \addr<4> ;
  assign N23 = \addr<5> ;
  assign N24 = \addr<6> ;
  assign N25 = \addr<7> ;

  DFFPOSX1 \mem_reg<0>  ( .D(n633), .CLK(clk), .Q(\mem<0> ) );
  DFFPOSX1 \mem_reg<1>  ( .D(n632), .CLK(clk), .Q(\mem<1> ) );
  DFFPOSX1 \mem_reg<2>  ( .D(n631), .CLK(clk), .Q(\mem<2> ) );
  DFFPOSX1 \mem_reg<3>  ( .D(n630), .CLK(clk), .Q(\mem<3> ) );
  DFFPOSX1 \mem_reg<4>  ( .D(n629), .CLK(clk), .Q(\mem<4> ) );
  DFFPOSX1 \mem_reg<5>  ( .D(n628), .CLK(clk), .Q(\mem<5> ) );
  DFFPOSX1 \mem_reg<6>  ( .D(n627), .CLK(clk), .Q(\mem<6> ) );
  DFFPOSX1 \mem_reg<7>  ( .D(n626), .CLK(clk), .Q(\mem<7> ) );
  DFFPOSX1 \mem_reg<8>  ( .D(n625), .CLK(clk), .Q(\mem<8> ) );
  DFFPOSX1 \mem_reg<9>  ( .D(n624), .CLK(clk), .Q(\mem<9> ) );
  DFFPOSX1 \mem_reg<10>  ( .D(n623), .CLK(clk), .Q(\mem<10> ) );
  DFFPOSX1 \mem_reg<11>  ( .D(n622), .CLK(clk), .Q(\mem<11> ) );
  DFFPOSX1 \mem_reg<12>  ( .D(n621), .CLK(clk), .Q(\mem<12> ) );
  DFFPOSX1 \mem_reg<13>  ( .D(n620), .CLK(clk), .Q(\mem<13> ) );
  DFFPOSX1 \mem_reg<14>  ( .D(n619), .CLK(clk), .Q(\mem<14> ) );
  DFFPOSX1 \mem_reg<15>  ( .D(n618), .CLK(clk), .Q(\mem<15> ) );
  DFFPOSX1 \mem_reg<16>  ( .D(n617), .CLK(clk), .Q(\mem<16> ) );
  DFFPOSX1 \mem_reg<17>  ( .D(n616), .CLK(clk), .Q(\mem<17> ) );
  DFFPOSX1 \mem_reg<18>  ( .D(n615), .CLK(clk), .Q(\mem<18> ) );
  DFFPOSX1 \mem_reg<19>  ( .D(n614), .CLK(clk), .Q(\mem<19> ) );
  DFFPOSX1 \mem_reg<20>  ( .D(n613), .CLK(clk), .Q(\mem<20> ) );
  DFFPOSX1 \mem_reg<21>  ( .D(n612), .CLK(clk), .Q(\mem<21> ) );
  DFFPOSX1 \mem_reg<22>  ( .D(n611), .CLK(clk), .Q(\mem<22> ) );
  DFFPOSX1 \mem_reg<23>  ( .D(n610), .CLK(clk), .Q(\mem<23> ) );
  DFFPOSX1 \mem_reg<24>  ( .D(n609), .CLK(clk), .Q(\mem<24> ) );
  DFFPOSX1 \mem_reg<25>  ( .D(n608), .CLK(clk), .Q(\mem<25> ) );
  DFFPOSX1 \mem_reg<26>  ( .D(n607), .CLK(clk), .Q(\mem<26> ) );
  DFFPOSX1 \mem_reg<27>  ( .D(n606), .CLK(clk), .Q(\mem<27> ) );
  DFFPOSX1 \mem_reg<28>  ( .D(n605), .CLK(clk), .Q(\mem<28> ) );
  DFFPOSX1 \mem_reg<29>  ( .D(n604), .CLK(clk), .Q(\mem<29> ) );
  DFFPOSX1 \mem_reg<30>  ( .D(n603), .CLK(clk), .Q(\mem<30> ) );
  DFFPOSX1 \mem_reg<31>  ( .D(n602), .CLK(clk), .Q(\mem<31> ) );
  DFFPOSX1 \mem_reg<32>  ( .D(n601), .CLK(clk), .Q(\mem<32> ) );
  DFFPOSX1 \mem_reg<33>  ( .D(n600), .CLK(clk), .Q(\mem<33> ) );
  DFFPOSX1 \mem_reg<34>  ( .D(n599), .CLK(clk), .Q(\mem<34> ) );
  DFFPOSX1 \mem_reg<35>  ( .D(n598), .CLK(clk), .Q(\mem<35> ) );
  DFFPOSX1 \mem_reg<36>  ( .D(n597), .CLK(clk), .Q(\mem<36> ) );
  DFFPOSX1 \mem_reg<37>  ( .D(n596), .CLK(clk), .Q(\mem<37> ) );
  DFFPOSX1 \mem_reg<38>  ( .D(n595), .CLK(clk), .Q(\mem<38> ) );
  DFFPOSX1 \mem_reg<39>  ( .D(n594), .CLK(clk), .Q(\mem<39> ) );
  DFFPOSX1 \mem_reg<40>  ( .D(n593), .CLK(clk), .Q(\mem<40> ) );
  DFFPOSX1 \mem_reg<41>  ( .D(n592), .CLK(clk), .Q(\mem<41> ) );
  DFFPOSX1 \mem_reg<42>  ( .D(n591), .CLK(clk), .Q(\mem<42> ) );
  DFFPOSX1 \mem_reg<43>  ( .D(n590), .CLK(clk), .Q(\mem<43> ) );
  DFFPOSX1 \mem_reg<44>  ( .D(n589), .CLK(clk), .Q(\mem<44> ) );
  DFFPOSX1 \mem_reg<45>  ( .D(n588), .CLK(clk), .Q(\mem<45> ) );
  DFFPOSX1 \mem_reg<46>  ( .D(n587), .CLK(clk), .Q(\mem<46> ) );
  DFFPOSX1 \mem_reg<47>  ( .D(n586), .CLK(clk), .Q(\mem<47> ) );
  DFFPOSX1 \mem_reg<48>  ( .D(n585), .CLK(clk), .Q(\mem<48> ) );
  DFFPOSX1 \mem_reg<49>  ( .D(n584), .CLK(clk), .Q(\mem<49> ) );
  DFFPOSX1 \mem_reg<50>  ( .D(n583), .CLK(clk), .Q(\mem<50> ) );
  DFFPOSX1 \mem_reg<51>  ( .D(n582), .CLK(clk), .Q(\mem<51> ) );
  DFFPOSX1 \mem_reg<52>  ( .D(n581), .CLK(clk), .Q(\mem<52> ) );
  DFFPOSX1 \mem_reg<53>  ( .D(n580), .CLK(clk), .Q(\mem<53> ) );
  DFFPOSX1 \mem_reg<54>  ( .D(n579), .CLK(clk), .Q(\mem<54> ) );
  DFFPOSX1 \mem_reg<55>  ( .D(n578), .CLK(clk), .Q(\mem<55> ) );
  DFFPOSX1 \mem_reg<56>  ( .D(n577), .CLK(clk), .Q(\mem<56> ) );
  DFFPOSX1 \mem_reg<57>  ( .D(n576), .CLK(clk), .Q(\mem<57> ) );
  DFFPOSX1 \mem_reg<58>  ( .D(n575), .CLK(clk), .Q(\mem<58> ) );
  DFFPOSX1 \mem_reg<59>  ( .D(n574), .CLK(clk), .Q(\mem<59> ) );
  DFFPOSX1 \mem_reg<60>  ( .D(n573), .CLK(clk), .Q(\mem<60> ) );
  DFFPOSX1 \mem_reg<61>  ( .D(n572), .CLK(clk), .Q(\mem<61> ) );
  DFFPOSX1 \mem_reg<62>  ( .D(n571), .CLK(clk), .Q(\mem<62> ) );
  DFFPOSX1 \mem_reg<63>  ( .D(n570), .CLK(clk), .Q(\mem<63> ) );
  DFFPOSX1 \mem_reg<64>  ( .D(n569), .CLK(clk), .Q(\mem<64> ) );
  DFFPOSX1 \mem_reg<65>  ( .D(n568), .CLK(clk), .Q(\mem<65> ) );
  DFFPOSX1 \mem_reg<66>  ( .D(n567), .CLK(clk), .Q(\mem<66> ) );
  DFFPOSX1 \mem_reg<67>  ( .D(n566), .CLK(clk), .Q(\mem<67> ) );
  DFFPOSX1 \mem_reg<68>  ( .D(n565), .CLK(clk), .Q(\mem<68> ) );
  DFFPOSX1 \mem_reg<69>  ( .D(n564), .CLK(clk), .Q(\mem<69> ) );
  DFFPOSX1 \mem_reg<70>  ( .D(n563), .CLK(clk), .Q(\mem<70> ) );
  DFFPOSX1 \mem_reg<71>  ( .D(n562), .CLK(clk), .Q(\mem<71> ) );
  DFFPOSX1 \mem_reg<72>  ( .D(n561), .CLK(clk), .Q(\mem<72> ) );
  DFFPOSX1 \mem_reg<73>  ( .D(n560), .CLK(clk), .Q(\mem<73> ) );
  DFFPOSX1 \mem_reg<74>  ( .D(n559), .CLK(clk), .Q(\mem<74> ) );
  DFFPOSX1 \mem_reg<75>  ( .D(n558), .CLK(clk), .Q(\mem<75> ) );
  DFFPOSX1 \mem_reg<76>  ( .D(n557), .CLK(clk), .Q(\mem<76> ) );
  DFFPOSX1 \mem_reg<77>  ( .D(n556), .CLK(clk), .Q(\mem<77> ) );
  DFFPOSX1 \mem_reg<78>  ( .D(n555), .CLK(clk), .Q(\mem<78> ) );
  DFFPOSX1 \mem_reg<79>  ( .D(n554), .CLK(clk), .Q(\mem<79> ) );
  DFFPOSX1 \mem_reg<80>  ( .D(n553), .CLK(clk), .Q(\mem<80> ) );
  DFFPOSX1 \mem_reg<81>  ( .D(n552), .CLK(clk), .Q(\mem<81> ) );
  DFFPOSX1 \mem_reg<82>  ( .D(n551), .CLK(clk), .Q(\mem<82> ) );
  DFFPOSX1 \mem_reg<83>  ( .D(n550), .CLK(clk), .Q(\mem<83> ) );
  DFFPOSX1 \mem_reg<84>  ( .D(n549), .CLK(clk), .Q(\mem<84> ) );
  DFFPOSX1 \mem_reg<85>  ( .D(n548), .CLK(clk), .Q(\mem<85> ) );
  DFFPOSX1 \mem_reg<86>  ( .D(n547), .CLK(clk), .Q(\mem<86> ) );
  DFFPOSX1 \mem_reg<87>  ( .D(n546), .CLK(clk), .Q(\mem<87> ) );
  DFFPOSX1 \mem_reg<88>  ( .D(n545), .CLK(clk), .Q(\mem<88> ) );
  DFFPOSX1 \mem_reg<89>  ( .D(n544), .CLK(clk), .Q(\mem<89> ) );
  DFFPOSX1 \mem_reg<90>  ( .D(n543), .CLK(clk), .Q(\mem<90> ) );
  DFFPOSX1 \mem_reg<91>  ( .D(n542), .CLK(clk), .Q(\mem<91> ) );
  DFFPOSX1 \mem_reg<92>  ( .D(n541), .CLK(clk), .Q(\mem<92> ) );
  DFFPOSX1 \mem_reg<93>  ( .D(n540), .CLK(clk), .Q(\mem<93> ) );
  DFFPOSX1 \mem_reg<94>  ( .D(n539), .CLK(clk), .Q(\mem<94> ) );
  DFFPOSX1 \mem_reg<95>  ( .D(n538), .CLK(clk), .Q(\mem<95> ) );
  DFFPOSX1 \mem_reg<96>  ( .D(n537), .CLK(clk), .Q(\mem<96> ) );
  DFFPOSX1 \mem_reg<97>  ( .D(n536), .CLK(clk), .Q(\mem<97> ) );
  DFFPOSX1 \mem_reg<98>  ( .D(n535), .CLK(clk), .Q(\mem<98> ) );
  DFFPOSX1 \mem_reg<99>  ( .D(n534), .CLK(clk), .Q(\mem<99> ) );
  DFFPOSX1 \mem_reg<100>  ( .D(n533), .CLK(clk), .Q(\mem<100> ) );
  DFFPOSX1 \mem_reg<101>  ( .D(n532), .CLK(clk), .Q(\mem<101> ) );
  DFFPOSX1 \mem_reg<102>  ( .D(n531), .CLK(clk), .Q(\mem<102> ) );
  DFFPOSX1 \mem_reg<103>  ( .D(n530), .CLK(clk), .Q(\mem<103> ) );
  DFFPOSX1 \mem_reg<104>  ( .D(n529), .CLK(clk), .Q(\mem<104> ) );
  DFFPOSX1 \mem_reg<105>  ( .D(n528), .CLK(clk), .Q(\mem<105> ) );
  DFFPOSX1 \mem_reg<106>  ( .D(n527), .CLK(clk), .Q(\mem<106> ) );
  DFFPOSX1 \mem_reg<107>  ( .D(n526), .CLK(clk), .Q(\mem<107> ) );
  DFFPOSX1 \mem_reg<108>  ( .D(n525), .CLK(clk), .Q(\mem<108> ) );
  DFFPOSX1 \mem_reg<109>  ( .D(n524), .CLK(clk), .Q(\mem<109> ) );
  DFFPOSX1 \mem_reg<110>  ( .D(n523), .CLK(clk), .Q(\mem<110> ) );
  DFFPOSX1 \mem_reg<111>  ( .D(n522), .CLK(clk), .Q(\mem<111> ) );
  DFFPOSX1 \mem_reg<112>  ( .D(n521), .CLK(clk), .Q(\mem<112> ) );
  DFFPOSX1 \mem_reg<113>  ( .D(n520), .CLK(clk), .Q(\mem<113> ) );
  DFFPOSX1 \mem_reg<114>  ( .D(n519), .CLK(clk), .Q(\mem<114> ) );
  DFFPOSX1 \mem_reg<115>  ( .D(n518), .CLK(clk), .Q(\mem<115> ) );
  DFFPOSX1 \mem_reg<116>  ( .D(n517), .CLK(clk), .Q(\mem<116> ) );
  DFFPOSX1 \mem_reg<117>  ( .D(n516), .CLK(clk), .Q(\mem<117> ) );
  DFFPOSX1 \mem_reg<118>  ( .D(n515), .CLK(clk), .Q(\mem<118> ) );
  DFFPOSX1 \mem_reg<119>  ( .D(n514), .CLK(clk), .Q(\mem<119> ) );
  DFFPOSX1 \mem_reg<120>  ( .D(n513), .CLK(clk), .Q(\mem<120> ) );
  DFFPOSX1 \mem_reg<121>  ( .D(n512), .CLK(clk), .Q(\mem<121> ) );
  DFFPOSX1 \mem_reg<122>  ( .D(n511), .CLK(clk), .Q(\mem<122> ) );
  DFFPOSX1 \mem_reg<123>  ( .D(n510), .CLK(clk), .Q(\mem<123> ) );
  DFFPOSX1 \mem_reg<124>  ( .D(n509), .CLK(clk), .Q(\mem<124> ) );
  DFFPOSX1 \mem_reg<125>  ( .D(n508), .CLK(clk), .Q(\mem<125> ) );
  DFFPOSX1 \mem_reg<126>  ( .D(n507), .CLK(clk), .Q(\mem<126> ) );
  DFFPOSX1 \mem_reg<127>  ( .D(n506), .CLK(clk), .Q(\mem<127> ) );
  DFFPOSX1 \mem_reg<128>  ( .D(n505), .CLK(clk), .Q(\mem<128> ) );
  DFFPOSX1 \mem_reg<129>  ( .D(n504), .CLK(clk), .Q(\mem<129> ) );
  DFFPOSX1 \mem_reg<130>  ( .D(n503), .CLK(clk), .Q(\mem<130> ) );
  DFFPOSX1 \mem_reg<131>  ( .D(n502), .CLK(clk), .Q(\mem<131> ) );
  DFFPOSX1 \mem_reg<132>  ( .D(n501), .CLK(clk), .Q(\mem<132> ) );
  DFFPOSX1 \mem_reg<133>  ( .D(n500), .CLK(clk), .Q(\mem<133> ) );
  DFFPOSX1 \mem_reg<134>  ( .D(n499), .CLK(clk), .Q(\mem<134> ) );
  DFFPOSX1 \mem_reg<135>  ( .D(n498), .CLK(clk), .Q(\mem<135> ) );
  DFFPOSX1 \mem_reg<136>  ( .D(n497), .CLK(clk), .Q(\mem<136> ) );
  DFFPOSX1 \mem_reg<137>  ( .D(n496), .CLK(clk), .Q(\mem<137> ) );
  DFFPOSX1 \mem_reg<138>  ( .D(n495), .CLK(clk), .Q(\mem<138> ) );
  DFFPOSX1 \mem_reg<139>  ( .D(n494), .CLK(clk), .Q(\mem<139> ) );
  DFFPOSX1 \mem_reg<140>  ( .D(n493), .CLK(clk), .Q(\mem<140> ) );
  DFFPOSX1 \mem_reg<141>  ( .D(n492), .CLK(clk), .Q(\mem<141> ) );
  DFFPOSX1 \mem_reg<142>  ( .D(n491), .CLK(clk), .Q(\mem<142> ) );
  DFFPOSX1 \mem_reg<143>  ( .D(n490), .CLK(clk), .Q(\mem<143> ) );
  DFFPOSX1 \mem_reg<144>  ( .D(n489), .CLK(clk), .Q(\mem<144> ) );
  DFFPOSX1 \mem_reg<145>  ( .D(n488), .CLK(clk), .Q(\mem<145> ) );
  DFFPOSX1 \mem_reg<146>  ( .D(n487), .CLK(clk), .Q(\mem<146> ) );
  DFFPOSX1 \mem_reg<147>  ( .D(n486), .CLK(clk), .Q(\mem<147> ) );
  DFFPOSX1 \mem_reg<148>  ( .D(n485), .CLK(clk), .Q(\mem<148> ) );
  DFFPOSX1 \mem_reg<149>  ( .D(n484), .CLK(clk), .Q(\mem<149> ) );
  DFFPOSX1 \mem_reg<150>  ( .D(n483), .CLK(clk), .Q(\mem<150> ) );
  DFFPOSX1 \mem_reg<151>  ( .D(n482), .CLK(clk), .Q(\mem<151> ) );
  DFFPOSX1 \mem_reg<152>  ( .D(n481), .CLK(clk), .Q(\mem<152> ) );
  DFFPOSX1 \mem_reg<153>  ( .D(n480), .CLK(clk), .Q(\mem<153> ) );
  DFFPOSX1 \mem_reg<154>  ( .D(n479), .CLK(clk), .Q(\mem<154> ) );
  DFFPOSX1 \mem_reg<155>  ( .D(n478), .CLK(clk), .Q(\mem<155> ) );
  DFFPOSX1 \mem_reg<156>  ( .D(n477), .CLK(clk), .Q(\mem<156> ) );
  DFFPOSX1 \mem_reg<157>  ( .D(n476), .CLK(clk), .Q(\mem<157> ) );
  DFFPOSX1 \mem_reg<158>  ( .D(n475), .CLK(clk), .Q(\mem<158> ) );
  DFFPOSX1 \mem_reg<159>  ( .D(n474), .CLK(clk), .Q(\mem<159> ) );
  DFFPOSX1 \mem_reg<160>  ( .D(n473), .CLK(clk), .Q(\mem<160> ) );
  DFFPOSX1 \mem_reg<161>  ( .D(n472), .CLK(clk), .Q(\mem<161> ) );
  DFFPOSX1 \mem_reg<162>  ( .D(n471), .CLK(clk), .Q(\mem<162> ) );
  DFFPOSX1 \mem_reg<163>  ( .D(n470), .CLK(clk), .Q(\mem<163> ) );
  DFFPOSX1 \mem_reg<164>  ( .D(n469), .CLK(clk), .Q(\mem<164> ) );
  DFFPOSX1 \mem_reg<165>  ( .D(n468), .CLK(clk), .Q(\mem<165> ) );
  DFFPOSX1 \mem_reg<166>  ( .D(n467), .CLK(clk), .Q(\mem<166> ) );
  DFFPOSX1 \mem_reg<167>  ( .D(n466), .CLK(clk), .Q(\mem<167> ) );
  DFFPOSX1 \mem_reg<168>  ( .D(n465), .CLK(clk), .Q(\mem<168> ) );
  DFFPOSX1 \mem_reg<169>  ( .D(n464), .CLK(clk), .Q(\mem<169> ) );
  DFFPOSX1 \mem_reg<170>  ( .D(n463), .CLK(clk), .Q(\mem<170> ) );
  DFFPOSX1 \mem_reg<171>  ( .D(n462), .CLK(clk), .Q(\mem<171> ) );
  DFFPOSX1 \mem_reg<172>  ( .D(n461), .CLK(clk), .Q(\mem<172> ) );
  DFFPOSX1 \mem_reg<173>  ( .D(n460), .CLK(clk), .Q(\mem<173> ) );
  DFFPOSX1 \mem_reg<174>  ( .D(n459), .CLK(clk), .Q(\mem<174> ) );
  DFFPOSX1 \mem_reg<175>  ( .D(n458), .CLK(clk), .Q(\mem<175> ) );
  DFFPOSX1 \mem_reg<176>  ( .D(n457), .CLK(clk), .Q(\mem<176> ) );
  DFFPOSX1 \mem_reg<177>  ( .D(n456), .CLK(clk), .Q(\mem<177> ) );
  DFFPOSX1 \mem_reg<178>  ( .D(n455), .CLK(clk), .Q(\mem<178> ) );
  DFFPOSX1 \mem_reg<179>  ( .D(n454), .CLK(clk), .Q(\mem<179> ) );
  DFFPOSX1 \mem_reg<180>  ( .D(n453), .CLK(clk), .Q(\mem<180> ) );
  DFFPOSX1 \mem_reg<181>  ( .D(n452), .CLK(clk), .Q(\mem<181> ) );
  DFFPOSX1 \mem_reg<182>  ( .D(n451), .CLK(clk), .Q(\mem<182> ) );
  DFFPOSX1 \mem_reg<183>  ( .D(n450), .CLK(clk), .Q(\mem<183> ) );
  DFFPOSX1 \mem_reg<184>  ( .D(n449), .CLK(clk), .Q(\mem<184> ) );
  DFFPOSX1 \mem_reg<185>  ( .D(n448), .CLK(clk), .Q(\mem<185> ) );
  DFFPOSX1 \mem_reg<186>  ( .D(n447), .CLK(clk), .Q(\mem<186> ) );
  DFFPOSX1 \mem_reg<187>  ( .D(n446), .CLK(clk), .Q(\mem<187> ) );
  DFFPOSX1 \mem_reg<188>  ( .D(n445), .CLK(clk), .Q(\mem<188> ) );
  DFFPOSX1 \mem_reg<189>  ( .D(n444), .CLK(clk), .Q(\mem<189> ) );
  DFFPOSX1 \mem_reg<190>  ( .D(n443), .CLK(clk), .Q(\mem<190> ) );
  DFFPOSX1 \mem_reg<191>  ( .D(n442), .CLK(clk), .Q(\mem<191> ) );
  DFFPOSX1 \mem_reg<192>  ( .D(n441), .CLK(clk), .Q(\mem<192> ) );
  DFFPOSX1 \mem_reg<193>  ( .D(n440), .CLK(clk), .Q(\mem<193> ) );
  DFFPOSX1 \mem_reg<194>  ( .D(n439), .CLK(clk), .Q(\mem<194> ) );
  DFFPOSX1 \mem_reg<195>  ( .D(n438), .CLK(clk), .Q(\mem<195> ) );
  DFFPOSX1 \mem_reg<196>  ( .D(n437), .CLK(clk), .Q(\mem<196> ) );
  DFFPOSX1 \mem_reg<197>  ( .D(n436), .CLK(clk), .Q(\mem<197> ) );
  DFFPOSX1 \mem_reg<198>  ( .D(n435), .CLK(clk), .Q(\mem<198> ) );
  DFFPOSX1 \mem_reg<199>  ( .D(n434), .CLK(clk), .Q(\mem<199> ) );
  DFFPOSX1 \mem_reg<200>  ( .D(n433), .CLK(clk), .Q(\mem<200> ) );
  DFFPOSX1 \mem_reg<201>  ( .D(n432), .CLK(clk), .Q(\mem<201> ) );
  DFFPOSX1 \mem_reg<202>  ( .D(n431), .CLK(clk), .Q(\mem<202> ) );
  DFFPOSX1 \mem_reg<203>  ( .D(n430), .CLK(clk), .Q(\mem<203> ) );
  DFFPOSX1 \mem_reg<204>  ( .D(n429), .CLK(clk), .Q(\mem<204> ) );
  DFFPOSX1 \mem_reg<205>  ( .D(n428), .CLK(clk), .Q(\mem<205> ) );
  DFFPOSX1 \mem_reg<206>  ( .D(n427), .CLK(clk), .Q(\mem<206> ) );
  DFFPOSX1 \mem_reg<207>  ( .D(n426), .CLK(clk), .Q(\mem<207> ) );
  DFFPOSX1 \mem_reg<208>  ( .D(n425), .CLK(clk), .Q(\mem<208> ) );
  DFFPOSX1 \mem_reg<209>  ( .D(n424), .CLK(clk), .Q(\mem<209> ) );
  DFFPOSX1 \mem_reg<210>  ( .D(n423), .CLK(clk), .Q(\mem<210> ) );
  DFFPOSX1 \mem_reg<211>  ( .D(n422), .CLK(clk), .Q(\mem<211> ) );
  DFFPOSX1 \mem_reg<212>  ( .D(n421), .CLK(clk), .Q(\mem<212> ) );
  DFFPOSX1 \mem_reg<213>  ( .D(n420), .CLK(clk), .Q(\mem<213> ) );
  DFFPOSX1 \mem_reg<214>  ( .D(n419), .CLK(clk), .Q(\mem<214> ) );
  DFFPOSX1 \mem_reg<215>  ( .D(n418), .CLK(clk), .Q(\mem<215> ) );
  DFFPOSX1 \mem_reg<216>  ( .D(n417), .CLK(clk), .Q(\mem<216> ) );
  DFFPOSX1 \mem_reg<217>  ( .D(n416), .CLK(clk), .Q(\mem<217> ) );
  DFFPOSX1 \mem_reg<218>  ( .D(n415), .CLK(clk), .Q(\mem<218> ) );
  DFFPOSX1 \mem_reg<219>  ( .D(n414), .CLK(clk), .Q(\mem<219> ) );
  DFFPOSX1 \mem_reg<220>  ( .D(n413), .CLK(clk), .Q(\mem<220> ) );
  DFFPOSX1 \mem_reg<221>  ( .D(n412), .CLK(clk), .Q(\mem<221> ) );
  DFFPOSX1 \mem_reg<222>  ( .D(n411), .CLK(clk), .Q(\mem<222> ) );
  DFFPOSX1 \mem_reg<223>  ( .D(n410), .CLK(clk), .Q(\mem<223> ) );
  DFFPOSX1 \mem_reg<224>  ( .D(n409), .CLK(clk), .Q(\mem<224> ) );
  DFFPOSX1 \mem_reg<225>  ( .D(n408), .CLK(clk), .Q(\mem<225> ) );
  DFFPOSX1 \mem_reg<226>  ( .D(n407), .CLK(clk), .Q(\mem<226> ) );
  DFFPOSX1 \mem_reg<227>  ( .D(n406), .CLK(clk), .Q(\mem<227> ) );
  DFFPOSX1 \mem_reg<228>  ( .D(n405), .CLK(clk), .Q(\mem<228> ) );
  DFFPOSX1 \mem_reg<229>  ( .D(n404), .CLK(clk), .Q(\mem<229> ) );
  DFFPOSX1 \mem_reg<230>  ( .D(n403), .CLK(clk), .Q(\mem<230> ) );
  DFFPOSX1 \mem_reg<231>  ( .D(n402), .CLK(clk), .Q(\mem<231> ) );
  DFFPOSX1 \mem_reg<232>  ( .D(n401), .CLK(clk), .Q(\mem<232> ) );
  DFFPOSX1 \mem_reg<233>  ( .D(n400), .CLK(clk), .Q(\mem<233> ) );
  DFFPOSX1 \mem_reg<234>  ( .D(n399), .CLK(clk), .Q(\mem<234> ) );
  DFFPOSX1 \mem_reg<235>  ( .D(n398), .CLK(clk), .Q(\mem<235> ) );
  DFFPOSX1 \mem_reg<236>  ( .D(n397), .CLK(clk), .Q(\mem<236> ) );
  DFFPOSX1 \mem_reg<237>  ( .D(n396), .CLK(clk), .Q(\mem<237> ) );
  DFFPOSX1 \mem_reg<238>  ( .D(n395), .CLK(clk), .Q(\mem<238> ) );
  DFFPOSX1 \mem_reg<239>  ( .D(n394), .CLK(clk), .Q(\mem<239> ) );
  DFFPOSX1 \mem_reg<240>  ( .D(n393), .CLK(clk), .Q(\mem<240> ) );
  DFFPOSX1 \mem_reg<241>  ( .D(n392), .CLK(clk), .Q(\mem<241> ) );
  DFFPOSX1 \mem_reg<242>  ( .D(n391), .CLK(clk), .Q(\mem<242> ) );
  DFFPOSX1 \mem_reg<243>  ( .D(n390), .CLK(clk), .Q(\mem<243> ) );
  DFFPOSX1 \mem_reg<244>  ( .D(n389), .CLK(clk), .Q(\mem<244> ) );
  DFFPOSX1 \mem_reg<245>  ( .D(n388), .CLK(clk), .Q(\mem<245> ) );
  DFFPOSX1 \mem_reg<246>  ( .D(n387), .CLK(clk), .Q(\mem<246> ) );
  DFFPOSX1 \mem_reg<247>  ( .D(n386), .CLK(clk), .Q(\mem<247> ) );
  DFFPOSX1 \mem_reg<248>  ( .D(n385), .CLK(clk), .Q(\mem<248> ) );
  DFFPOSX1 \mem_reg<249>  ( .D(n384), .CLK(clk), .Q(\mem<249> ) );
  DFFPOSX1 \mem_reg<250>  ( .D(n383), .CLK(clk), .Q(\mem<250> ) );
  DFFPOSX1 \mem_reg<251>  ( .D(n382), .CLK(clk), .Q(\mem<251> ) );
  DFFPOSX1 \mem_reg<252>  ( .D(n381), .CLK(clk), .Q(\mem<252> ) );
  DFFPOSX1 \mem_reg<253>  ( .D(n380), .CLK(clk), .Q(\mem<253> ) );
  DFFPOSX1 \mem_reg<254>  ( .D(n379), .CLK(clk), .Q(\mem<254> ) );
  DFFPOSX1 \mem_reg<255>  ( .D(n378), .CLK(clk), .Q(\mem<255> ) );
  AND2X2 U6 ( .A(N21), .B(n982), .Y(n355) );
  AND2X2 U7 ( .A(N21), .B(n983), .Y(n364) );
  AND2X2 U8 ( .A(n980), .B(N18), .Y(n356) );
  AND2X2 U9 ( .A(n980), .B(n921), .Y(n358) );
  AND2X2 U10 ( .A(data_in), .B(n68), .Y(n90) );
  OAI21X1 U49 ( .A(n958), .B(n636), .C(n42), .Y(n378) );
  OAI21X1 U50 ( .A(n37), .B(n978), .C(\mem<255> ), .Y(n42) );
  OAI21X1 U51 ( .A(n636), .B(n955), .C(n46), .Y(n379) );
  OAI21X1 U52 ( .A(n979), .B(n35), .C(\mem<254> ), .Y(n46) );
  OAI21X1 U53 ( .A(n636), .B(n954), .C(n49), .Y(n380) );
  OAI21X1 U54 ( .A(n979), .B(n33), .C(\mem<253> ), .Y(n49) );
  OAI21X1 U55 ( .A(n636), .B(n953), .C(n52), .Y(n381) );
  OAI21X1 U56 ( .A(n979), .B(n31), .C(\mem<252> ), .Y(n52) );
  OAI21X1 U57 ( .A(n636), .B(n951), .C(n55), .Y(n382) );
  OAI21X1 U58 ( .A(n979), .B(n29), .C(\mem<251> ), .Y(n55) );
  OAI21X1 U59 ( .A(n636), .B(n949), .C(n58), .Y(n383) );
  OAI21X1 U60 ( .A(n979), .B(n27), .C(\mem<250> ), .Y(n58) );
  OAI21X1 U61 ( .A(n636), .B(n947), .C(n61), .Y(n384) );
  OAI21X1 U62 ( .A(n979), .B(n25), .C(\mem<249> ), .Y(n61) );
  OAI21X1 U63 ( .A(n636), .B(n945), .C(n64), .Y(n385) );
  OAI21X1 U64 ( .A(n979), .B(n23), .C(\mem<248> ), .Y(n64) );
  OAI21X1 U65 ( .A(n636), .B(n944), .C(n67), .Y(n386) );
  OAI21X1 U66 ( .A(n979), .B(n21), .C(\mem<247> ), .Y(n67) );
  OAI21X1 U67 ( .A(n636), .B(n943), .C(n70), .Y(n387) );
  OAI21X1 U68 ( .A(n978), .B(n19), .C(\mem<246> ), .Y(n70) );
  OAI21X1 U69 ( .A(n636), .B(n942), .C(n73), .Y(n388) );
  OAI21X1 U70 ( .A(n978), .B(n17), .C(\mem<245> ), .Y(n73) );
  OAI21X1 U71 ( .A(n636), .B(n941), .C(n76), .Y(n389) );
  OAI21X1 U72 ( .A(n978), .B(n15), .C(\mem<244> ), .Y(n76) );
  OAI21X1 U73 ( .A(n636), .B(n940), .C(n79), .Y(n390) );
  OAI21X1 U74 ( .A(n978), .B(n13), .C(\mem<243> ), .Y(n79) );
  OAI21X1 U75 ( .A(n636), .B(n939), .C(n82), .Y(n391) );
  OAI21X1 U76 ( .A(n978), .B(n11), .C(\mem<242> ), .Y(n82) );
  OAI21X1 U77 ( .A(n636), .B(n938), .C(n85), .Y(n392) );
  OAI21X1 U78 ( .A(n978), .B(n9), .C(\mem<241> ), .Y(n85) );
  OAI21X1 U79 ( .A(n636), .B(n936), .C(n88), .Y(n393) );
  OAI21X1 U80 ( .A(n978), .B(n7), .C(\mem<240> ), .Y(n88) );
  OAI21X1 U83 ( .A(n958), .B(n369), .C(n94), .Y(n394) );
  OAI21X1 U84 ( .A(n37), .B(n977), .C(\mem<239> ), .Y(n94) );
  OAI21X1 U85 ( .A(n956), .B(n369), .C(n96), .Y(n395) );
  OAI21X1 U86 ( .A(n35), .B(n977), .C(\mem<238> ), .Y(n96) );
  OAI21X1 U87 ( .A(n954), .B(n369), .C(n97), .Y(n396) );
  OAI21X1 U88 ( .A(n33), .B(n977), .C(\mem<237> ), .Y(n97) );
  OAI21X1 U89 ( .A(n953), .B(n369), .C(n98), .Y(n397) );
  OAI21X1 U90 ( .A(n31), .B(n977), .C(\mem<236> ), .Y(n98) );
  OAI21X1 U91 ( .A(n952), .B(n369), .C(n99), .Y(n398) );
  OAI21X1 U92 ( .A(n29), .B(n977), .C(\mem<235> ), .Y(n99) );
  OAI21X1 U93 ( .A(n950), .B(n369), .C(n100), .Y(n399) );
  OAI21X1 U94 ( .A(n27), .B(n977), .C(\mem<234> ), .Y(n100) );
  OAI21X1 U95 ( .A(n948), .B(n369), .C(n101), .Y(n400) );
  OAI21X1 U96 ( .A(n25), .B(n977), .C(\mem<233> ), .Y(n101) );
  OAI21X1 U97 ( .A(n946), .B(n369), .C(n102), .Y(n401) );
  OAI21X1 U98 ( .A(n23), .B(n977), .C(\mem<232> ), .Y(n102) );
  OAI21X1 U99 ( .A(n944), .B(n369), .C(n103), .Y(n402) );
  OAI21X1 U100 ( .A(n21), .B(n976), .C(\mem<231> ), .Y(n103) );
  OAI21X1 U101 ( .A(n943), .B(n369), .C(n104), .Y(n403) );
  OAI21X1 U102 ( .A(n19), .B(n976), .C(\mem<230> ), .Y(n104) );
  OAI21X1 U103 ( .A(n942), .B(n369), .C(n105), .Y(n404) );
  OAI21X1 U104 ( .A(n17), .B(n976), .C(\mem<229> ), .Y(n105) );
  OAI21X1 U105 ( .A(n941), .B(n369), .C(n106), .Y(n405) );
  OAI21X1 U106 ( .A(n15), .B(n976), .C(\mem<228> ), .Y(n106) );
  OAI21X1 U107 ( .A(n940), .B(n369), .C(n107), .Y(n406) );
  OAI21X1 U108 ( .A(n13), .B(n976), .C(\mem<227> ), .Y(n107) );
  OAI21X1 U109 ( .A(n939), .B(n369), .C(n108), .Y(n407) );
  OAI21X1 U110 ( .A(n11), .B(n976), .C(\mem<226> ), .Y(n108) );
  OAI21X1 U111 ( .A(n938), .B(n369), .C(n109), .Y(n408) );
  OAI21X1 U112 ( .A(n9), .B(n976), .C(\mem<225> ), .Y(n109) );
  OAI21X1 U113 ( .A(n936), .B(n369), .C(n110), .Y(n409) );
  OAI21X1 U114 ( .A(n7), .B(n976), .C(\mem<224> ), .Y(n110) );
  OAI21X1 U117 ( .A(n958), .B(n353), .C(n113), .Y(n410) );
  OAI21X1 U118 ( .A(n37), .B(n975), .C(\mem<223> ), .Y(n113) );
  OAI21X1 U119 ( .A(n956), .B(n353), .C(n115), .Y(n411) );
  OAI21X1 U120 ( .A(n35), .B(n975), .C(\mem<222> ), .Y(n115) );
  OAI21X1 U121 ( .A(n954), .B(n353), .C(n116), .Y(n412) );
  OAI21X1 U122 ( .A(n33), .B(n975), .C(\mem<221> ), .Y(n116) );
  OAI21X1 U123 ( .A(n953), .B(n353), .C(n117), .Y(n413) );
  OAI21X1 U124 ( .A(n31), .B(n975), .C(\mem<220> ), .Y(n117) );
  OAI21X1 U125 ( .A(n952), .B(n353), .C(n118), .Y(n414) );
  OAI21X1 U126 ( .A(n29), .B(n975), .C(\mem<219> ), .Y(n118) );
  OAI21X1 U127 ( .A(n950), .B(n353), .C(n119), .Y(n415) );
  OAI21X1 U128 ( .A(n27), .B(n975), .C(\mem<218> ), .Y(n119) );
  OAI21X1 U129 ( .A(n948), .B(n353), .C(n120), .Y(n416) );
  OAI21X1 U130 ( .A(n25), .B(n975), .C(\mem<217> ), .Y(n120) );
  OAI21X1 U131 ( .A(n946), .B(n353), .C(n121), .Y(n417) );
  OAI21X1 U132 ( .A(n23), .B(n975), .C(\mem<216> ), .Y(n121) );
  OAI21X1 U133 ( .A(n944), .B(n353), .C(n122), .Y(n418) );
  OAI21X1 U134 ( .A(n21), .B(n975), .C(\mem<215> ), .Y(n122) );
  OAI21X1 U135 ( .A(n943), .B(n353), .C(n123), .Y(n419) );
  OAI21X1 U136 ( .A(n19), .B(n975), .C(\mem<214> ), .Y(n123) );
  OAI21X1 U137 ( .A(n942), .B(n353), .C(n124), .Y(n420) );
  OAI21X1 U138 ( .A(n17), .B(n975), .C(\mem<213> ), .Y(n124) );
  OAI21X1 U139 ( .A(n941), .B(n353), .C(n125), .Y(n421) );
  OAI21X1 U140 ( .A(n15), .B(n975), .C(\mem<212> ), .Y(n125) );
  OAI21X1 U141 ( .A(n940), .B(n353), .C(n126), .Y(n422) );
  OAI21X1 U142 ( .A(n13), .B(n975), .C(\mem<211> ), .Y(n126) );
  OAI21X1 U143 ( .A(n939), .B(n353), .C(n127), .Y(n423) );
  OAI21X1 U144 ( .A(n11), .B(n975), .C(\mem<210> ), .Y(n127) );
  OAI21X1 U145 ( .A(n938), .B(n353), .C(n128), .Y(n424) );
  OAI21X1 U146 ( .A(n9), .B(n975), .C(\mem<209> ), .Y(n128) );
  OAI21X1 U147 ( .A(n936), .B(n353), .C(n129), .Y(n425) );
  OAI21X1 U148 ( .A(n7), .B(n975), .C(\mem<208> ), .Y(n129) );
  OAI21X1 U151 ( .A(n958), .B(n335), .C(n132), .Y(n426) );
  OAI21X1 U152 ( .A(n37), .B(n974), .C(\mem<207> ), .Y(n132) );
  OAI21X1 U153 ( .A(n956), .B(n335), .C(n134), .Y(n427) );
  OAI21X1 U154 ( .A(n35), .B(n974), .C(\mem<206> ), .Y(n134) );
  OAI21X1 U155 ( .A(n954), .B(n335), .C(n135), .Y(n428) );
  OAI21X1 U156 ( .A(n33), .B(n974), .C(\mem<205> ), .Y(n135) );
  OAI21X1 U157 ( .A(n953), .B(n335), .C(n136), .Y(n429) );
  OAI21X1 U158 ( .A(n31), .B(n974), .C(\mem<204> ), .Y(n136) );
  OAI21X1 U159 ( .A(n952), .B(n335), .C(n137), .Y(n430) );
  OAI21X1 U160 ( .A(n29), .B(n974), .C(\mem<203> ), .Y(n137) );
  OAI21X1 U161 ( .A(n950), .B(n335), .C(n138), .Y(n431) );
  OAI21X1 U162 ( .A(n27), .B(n974), .C(\mem<202> ), .Y(n138) );
  OAI21X1 U163 ( .A(n948), .B(n335), .C(n139), .Y(n432) );
  OAI21X1 U164 ( .A(n25), .B(n974), .C(\mem<201> ), .Y(n139) );
  OAI21X1 U165 ( .A(n946), .B(n335), .C(n140), .Y(n433) );
  OAI21X1 U166 ( .A(n23), .B(n974), .C(\mem<200> ), .Y(n140) );
  OAI21X1 U167 ( .A(n944), .B(n335), .C(n141), .Y(n434) );
  OAI21X1 U168 ( .A(n21), .B(n974), .C(\mem<199> ), .Y(n141) );
  OAI21X1 U169 ( .A(n943), .B(n335), .C(n142), .Y(n435) );
  OAI21X1 U170 ( .A(n19), .B(n974), .C(\mem<198> ), .Y(n142) );
  OAI21X1 U171 ( .A(n942), .B(n335), .C(n143), .Y(n436) );
  OAI21X1 U172 ( .A(n17), .B(n974), .C(\mem<197> ), .Y(n143) );
  OAI21X1 U173 ( .A(n941), .B(n335), .C(n144), .Y(n437) );
  OAI21X1 U174 ( .A(n15), .B(n974), .C(\mem<196> ), .Y(n144) );
  OAI21X1 U175 ( .A(n940), .B(n335), .C(n145), .Y(n438) );
  OAI21X1 U176 ( .A(n13), .B(n974), .C(\mem<195> ), .Y(n145) );
  OAI21X1 U177 ( .A(n939), .B(n335), .C(n146), .Y(n439) );
  OAI21X1 U178 ( .A(n11), .B(n974), .C(\mem<194> ), .Y(n146) );
  OAI21X1 U179 ( .A(n938), .B(n335), .C(n147), .Y(n440) );
  OAI21X1 U180 ( .A(n9), .B(n974), .C(\mem<193> ), .Y(n147) );
  OAI21X1 U181 ( .A(n936), .B(n335), .C(n148), .Y(n441) );
  OAI21X1 U182 ( .A(n7), .B(n974), .C(\mem<192> ), .Y(n148) );
  OAI21X1 U185 ( .A(n958), .B(n317), .C(n151), .Y(n442) );
  OAI21X1 U186 ( .A(n37), .B(n973), .C(\mem<191> ), .Y(n151) );
  OAI21X1 U187 ( .A(n956), .B(n317), .C(n153), .Y(n443) );
  OAI21X1 U188 ( .A(n35), .B(n973), .C(\mem<190> ), .Y(n153) );
  OAI21X1 U189 ( .A(n954), .B(n317), .C(n154), .Y(n444) );
  OAI21X1 U190 ( .A(n33), .B(n973), .C(\mem<189> ), .Y(n154) );
  OAI21X1 U191 ( .A(n953), .B(n317), .C(n155), .Y(n445) );
  OAI21X1 U192 ( .A(n31), .B(n973), .C(\mem<188> ), .Y(n155) );
  OAI21X1 U193 ( .A(n952), .B(n317), .C(n156), .Y(n446) );
  OAI21X1 U194 ( .A(n29), .B(n973), .C(\mem<187> ), .Y(n156) );
  OAI21X1 U195 ( .A(n950), .B(n317), .C(n157), .Y(n447) );
  OAI21X1 U196 ( .A(n27), .B(n973), .C(\mem<186> ), .Y(n157) );
  OAI21X1 U197 ( .A(n948), .B(n317), .C(n158), .Y(n448) );
  OAI21X1 U198 ( .A(n25), .B(n973), .C(\mem<185> ), .Y(n158) );
  OAI21X1 U199 ( .A(n946), .B(n317), .C(n159), .Y(n449) );
  OAI21X1 U200 ( .A(n23), .B(n973), .C(\mem<184> ), .Y(n159) );
  OAI21X1 U201 ( .A(n944), .B(n317), .C(n160), .Y(n450) );
  OAI21X1 U202 ( .A(n21), .B(n972), .C(\mem<183> ), .Y(n160) );
  OAI21X1 U203 ( .A(n943), .B(n317), .C(n161), .Y(n451) );
  OAI21X1 U204 ( .A(n19), .B(n972), .C(\mem<182> ), .Y(n161) );
  OAI21X1 U205 ( .A(n942), .B(n317), .C(n162), .Y(n452) );
  OAI21X1 U206 ( .A(n17), .B(n972), .C(\mem<181> ), .Y(n162) );
  OAI21X1 U207 ( .A(n941), .B(n317), .C(n163), .Y(n453) );
  OAI21X1 U208 ( .A(n15), .B(n972), .C(\mem<180> ), .Y(n163) );
  OAI21X1 U209 ( .A(n940), .B(n317), .C(n164), .Y(n454) );
  OAI21X1 U210 ( .A(n13), .B(n972), .C(\mem<179> ), .Y(n164) );
  OAI21X1 U211 ( .A(n939), .B(n317), .C(n165), .Y(n455) );
  OAI21X1 U212 ( .A(n11), .B(n972), .C(\mem<178> ), .Y(n165) );
  OAI21X1 U213 ( .A(n938), .B(n317), .C(n166), .Y(n456) );
  OAI21X1 U214 ( .A(n9), .B(n972), .C(\mem<177> ), .Y(n166) );
  OAI21X1 U215 ( .A(n936), .B(n317), .C(n167), .Y(n457) );
  OAI21X1 U216 ( .A(n7), .B(n972), .C(\mem<176> ), .Y(n167) );
  OAI21X1 U219 ( .A(n958), .B(n296), .C(n170), .Y(n458) );
  OAI21X1 U220 ( .A(n37), .B(n971), .C(\mem<175> ), .Y(n170) );
  OAI21X1 U221 ( .A(n956), .B(n296), .C(n172), .Y(n459) );
  OAI21X1 U222 ( .A(n35), .B(n971), .C(\mem<174> ), .Y(n172) );
  OAI21X1 U223 ( .A(n954), .B(n296), .C(n173), .Y(n460) );
  OAI21X1 U224 ( .A(n33), .B(n971), .C(\mem<173> ), .Y(n173) );
  OAI21X1 U225 ( .A(n953), .B(n296), .C(n174), .Y(n461) );
  OAI21X1 U226 ( .A(n31), .B(n971), .C(\mem<172> ), .Y(n174) );
  OAI21X1 U227 ( .A(n952), .B(n296), .C(n175), .Y(n462) );
  OAI21X1 U228 ( .A(n29), .B(n971), .C(\mem<171> ), .Y(n175) );
  OAI21X1 U229 ( .A(n950), .B(n296), .C(n176), .Y(n463) );
  OAI21X1 U230 ( .A(n27), .B(n971), .C(\mem<170> ), .Y(n176) );
  OAI21X1 U231 ( .A(n948), .B(n296), .C(n177), .Y(n464) );
  OAI21X1 U232 ( .A(n25), .B(n971), .C(\mem<169> ), .Y(n177) );
  OAI21X1 U233 ( .A(n946), .B(n296), .C(n178), .Y(n465) );
  OAI21X1 U234 ( .A(n23), .B(n971), .C(\mem<168> ), .Y(n178) );
  OAI21X1 U235 ( .A(n944), .B(n296), .C(n179), .Y(n466) );
  OAI21X1 U236 ( .A(n21), .B(n970), .C(\mem<167> ), .Y(n179) );
  OAI21X1 U237 ( .A(n943), .B(n296), .C(n180), .Y(n467) );
  OAI21X1 U238 ( .A(n19), .B(n970), .C(\mem<166> ), .Y(n180) );
  OAI21X1 U239 ( .A(n942), .B(n296), .C(n181), .Y(n468) );
  OAI21X1 U240 ( .A(n17), .B(n970), .C(\mem<165> ), .Y(n181) );
  OAI21X1 U241 ( .A(n941), .B(n296), .C(n182), .Y(n469) );
  OAI21X1 U242 ( .A(n15), .B(n970), .C(\mem<164> ), .Y(n182) );
  OAI21X1 U243 ( .A(n940), .B(n296), .C(n183), .Y(n470) );
  OAI21X1 U244 ( .A(n13), .B(n970), .C(\mem<163> ), .Y(n183) );
  OAI21X1 U245 ( .A(n939), .B(n296), .C(n184), .Y(n471) );
  OAI21X1 U246 ( .A(n11), .B(n970), .C(\mem<162> ), .Y(n184) );
  OAI21X1 U247 ( .A(n938), .B(n296), .C(n185), .Y(n472) );
  OAI21X1 U248 ( .A(n9), .B(n970), .C(\mem<161> ), .Y(n185) );
  OAI21X1 U249 ( .A(n936), .B(n296), .C(n186), .Y(n473) );
  OAI21X1 U250 ( .A(n7), .B(n970), .C(\mem<160> ), .Y(n186) );
  OAI21X1 U253 ( .A(n958), .B(n260), .C(n188), .Y(n474) );
  OAI21X1 U254 ( .A(n37), .B(n969), .C(\mem<159> ), .Y(n188) );
  OAI21X1 U255 ( .A(n956), .B(n260), .C(n190), .Y(n475) );
  OAI21X1 U256 ( .A(n35), .B(n969), .C(\mem<158> ), .Y(n190) );
  OAI21X1 U257 ( .A(n954), .B(n260), .C(n191), .Y(n476) );
  OAI21X1 U258 ( .A(n33), .B(n969), .C(\mem<157> ), .Y(n191) );
  OAI21X1 U259 ( .A(n953), .B(n260), .C(n192), .Y(n477) );
  OAI21X1 U260 ( .A(n31), .B(n969), .C(\mem<156> ), .Y(n192) );
  OAI21X1 U261 ( .A(n952), .B(n260), .C(n193), .Y(n478) );
  OAI21X1 U262 ( .A(n29), .B(n969), .C(\mem<155> ), .Y(n193) );
  OAI21X1 U263 ( .A(n950), .B(n260), .C(n194), .Y(n479) );
  OAI21X1 U264 ( .A(n27), .B(n969), .C(\mem<154> ), .Y(n194) );
  OAI21X1 U265 ( .A(n948), .B(n260), .C(n195), .Y(n480) );
  OAI21X1 U266 ( .A(n25), .B(n969), .C(\mem<153> ), .Y(n195) );
  OAI21X1 U267 ( .A(n946), .B(n260), .C(n196), .Y(n481) );
  OAI21X1 U268 ( .A(n23), .B(n969), .C(\mem<152> ), .Y(n196) );
  OAI21X1 U269 ( .A(n944), .B(n260), .C(n197), .Y(n482) );
  OAI21X1 U270 ( .A(n21), .B(n968), .C(\mem<151> ), .Y(n197) );
  OAI21X1 U271 ( .A(n943), .B(n260), .C(n198), .Y(n483) );
  OAI21X1 U272 ( .A(n19), .B(n968), .C(\mem<150> ), .Y(n198) );
  OAI21X1 U273 ( .A(n942), .B(n260), .C(n199), .Y(n484) );
  OAI21X1 U274 ( .A(n17), .B(n968), .C(\mem<149> ), .Y(n199) );
  OAI21X1 U275 ( .A(n941), .B(n260), .C(n200), .Y(n485) );
  OAI21X1 U276 ( .A(n15), .B(n968), .C(\mem<148> ), .Y(n200) );
  OAI21X1 U277 ( .A(n940), .B(n260), .C(n201), .Y(n486) );
  OAI21X1 U278 ( .A(n13), .B(n968), .C(\mem<147> ), .Y(n201) );
  OAI21X1 U279 ( .A(n939), .B(n260), .C(n202), .Y(n487) );
  OAI21X1 U280 ( .A(n11), .B(n968), .C(\mem<146> ), .Y(n202) );
  OAI21X1 U281 ( .A(n938), .B(n260), .C(n203), .Y(n488) );
  OAI21X1 U282 ( .A(n9), .B(n968), .C(\mem<145> ), .Y(n203) );
  OAI21X1 U283 ( .A(n936), .B(n260), .C(n204), .Y(n489) );
  OAI21X1 U284 ( .A(n7), .B(n968), .C(\mem<144> ), .Y(n204) );
  OAI21X1 U287 ( .A(n958), .B(n225), .C(n206), .Y(n490) );
  OAI21X1 U288 ( .A(n37), .B(n967), .C(\mem<143> ), .Y(n206) );
  OAI21X1 U289 ( .A(n956), .B(n225), .C(n208), .Y(n491) );
  OAI21X1 U290 ( .A(n35), .B(n967), .C(\mem<142> ), .Y(n208) );
  OAI21X1 U291 ( .A(n954), .B(n225), .C(n209), .Y(n492) );
  OAI21X1 U292 ( .A(n33), .B(n967), .C(\mem<141> ), .Y(n209) );
  OAI21X1 U293 ( .A(n953), .B(n225), .C(n210), .Y(n493) );
  OAI21X1 U294 ( .A(n31), .B(n967), .C(\mem<140> ), .Y(n210) );
  OAI21X1 U295 ( .A(n952), .B(n225), .C(n211), .Y(n494) );
  OAI21X1 U296 ( .A(n29), .B(n967), .C(\mem<139> ), .Y(n211) );
  OAI21X1 U297 ( .A(n950), .B(n225), .C(n212), .Y(n495) );
  OAI21X1 U298 ( .A(n27), .B(n967), .C(\mem<138> ), .Y(n212) );
  OAI21X1 U299 ( .A(n948), .B(n225), .C(n213), .Y(n496) );
  OAI21X1 U300 ( .A(n25), .B(n967), .C(\mem<137> ), .Y(n213) );
  OAI21X1 U301 ( .A(n946), .B(n225), .C(n214), .Y(n497) );
  OAI21X1 U302 ( .A(n23), .B(n967), .C(\mem<136> ), .Y(n214) );
  OAI21X1 U303 ( .A(n944), .B(n225), .C(n215), .Y(n498) );
  OAI21X1 U304 ( .A(n21), .B(n966), .C(\mem<135> ), .Y(n215) );
  OAI21X1 U305 ( .A(n943), .B(n225), .C(n216), .Y(n499) );
  OAI21X1 U306 ( .A(n19), .B(n966), .C(\mem<134> ), .Y(n216) );
  OAI21X1 U307 ( .A(n942), .B(n225), .C(n217), .Y(n500) );
  OAI21X1 U308 ( .A(n17), .B(n966), .C(\mem<133> ), .Y(n217) );
  OAI21X1 U309 ( .A(n941), .B(n225), .C(n218), .Y(n501) );
  OAI21X1 U310 ( .A(n15), .B(n966), .C(\mem<132> ), .Y(n218) );
  OAI21X1 U311 ( .A(n940), .B(n225), .C(n219), .Y(n502) );
  OAI21X1 U312 ( .A(n13), .B(n966), .C(\mem<131> ), .Y(n219) );
  OAI21X1 U313 ( .A(n939), .B(n225), .C(n220), .Y(n503) );
  OAI21X1 U314 ( .A(n11), .B(n966), .C(\mem<130> ), .Y(n220) );
  OAI21X1 U315 ( .A(n938), .B(n225), .C(n221), .Y(n504) );
  OAI21X1 U316 ( .A(n9), .B(n966), .C(\mem<129> ), .Y(n221) );
  OAI21X1 U317 ( .A(n936), .B(n225), .C(n222), .Y(n505) );
  OAI21X1 U318 ( .A(n7), .B(n966), .C(\mem<128> ), .Y(n222) );
  OAI21X1 U321 ( .A(n957), .B(n189), .C(n224), .Y(n506) );
  OAI21X1 U322 ( .A(n37), .B(n965), .C(\mem<127> ), .Y(n224) );
  OAI21X1 U323 ( .A(n956), .B(n189), .C(n226), .Y(n507) );
  OAI21X1 U324 ( .A(n35), .B(n965), .C(\mem<126> ), .Y(n226) );
  OAI21X1 U325 ( .A(n954), .B(n189), .C(n227), .Y(n508) );
  OAI21X1 U326 ( .A(n33), .B(n965), .C(\mem<125> ), .Y(n227) );
  OAI21X1 U327 ( .A(n953), .B(n189), .C(n228), .Y(n509) );
  OAI21X1 U328 ( .A(n31), .B(n965), .C(\mem<124> ), .Y(n228) );
  OAI21X1 U329 ( .A(n952), .B(n189), .C(n229), .Y(n510) );
  OAI21X1 U330 ( .A(n29), .B(n965), .C(\mem<123> ), .Y(n229) );
  OAI21X1 U331 ( .A(n950), .B(n189), .C(n230), .Y(n511) );
  OAI21X1 U332 ( .A(n27), .B(n965), .C(\mem<122> ), .Y(n230) );
  OAI21X1 U333 ( .A(n948), .B(n189), .C(n231), .Y(n512) );
  OAI21X1 U334 ( .A(n25), .B(n965), .C(\mem<121> ), .Y(n231) );
  OAI21X1 U335 ( .A(n946), .B(n189), .C(n232), .Y(n513) );
  OAI21X1 U336 ( .A(n23), .B(n965), .C(\mem<120> ), .Y(n232) );
  OAI21X1 U337 ( .A(n944), .B(n189), .C(n233), .Y(n514) );
  OAI21X1 U338 ( .A(n21), .B(n965), .C(\mem<119> ), .Y(n233) );
  OAI21X1 U339 ( .A(n943), .B(n189), .C(n234), .Y(n515) );
  OAI21X1 U340 ( .A(n19), .B(n965), .C(\mem<118> ), .Y(n234) );
  OAI21X1 U341 ( .A(n942), .B(n189), .C(n235), .Y(n516) );
  OAI21X1 U342 ( .A(n17), .B(n965), .C(\mem<117> ), .Y(n235) );
  OAI21X1 U343 ( .A(n941), .B(n189), .C(n236), .Y(n517) );
  OAI21X1 U344 ( .A(n15), .B(n965), .C(\mem<116> ), .Y(n236) );
  OAI21X1 U345 ( .A(n940), .B(n189), .C(n237), .Y(n518) );
  OAI21X1 U346 ( .A(n13), .B(n965), .C(\mem<115> ), .Y(n237) );
  OAI21X1 U347 ( .A(n939), .B(n189), .C(n238), .Y(n519) );
  OAI21X1 U348 ( .A(n11), .B(n965), .C(\mem<114> ), .Y(n238) );
  OAI21X1 U349 ( .A(n938), .B(n189), .C(n239), .Y(n520) );
  OAI21X1 U350 ( .A(n9), .B(n965), .C(\mem<113> ), .Y(n239) );
  OAI21X1 U351 ( .A(n936), .B(n189), .C(n240), .Y(n521) );
  OAI21X1 U352 ( .A(n7), .B(n965), .C(\mem<112> ), .Y(n240) );
  OAI21X1 U355 ( .A(n957), .B(n171), .C(n243), .Y(n522) );
  OAI21X1 U356 ( .A(n37), .B(n964), .C(\mem<111> ), .Y(n243) );
  OAI21X1 U357 ( .A(n955), .B(n171), .C(n245), .Y(n523) );
  OAI21X1 U358 ( .A(n35), .B(n964), .C(\mem<110> ), .Y(n245) );
  OAI21X1 U359 ( .A(n954), .B(n171), .C(n246), .Y(n524) );
  OAI21X1 U360 ( .A(n33), .B(n964), .C(\mem<109> ), .Y(n246) );
  OAI21X1 U361 ( .A(n953), .B(n171), .C(n247), .Y(n525) );
  OAI21X1 U362 ( .A(n31), .B(n964), .C(\mem<108> ), .Y(n247) );
  OAI21X1 U363 ( .A(n951), .B(n171), .C(n248), .Y(n526) );
  OAI21X1 U364 ( .A(n29), .B(n964), .C(\mem<107> ), .Y(n248) );
  OAI21X1 U365 ( .A(n949), .B(n171), .C(n249), .Y(n527) );
  OAI21X1 U366 ( .A(n27), .B(n964), .C(\mem<106> ), .Y(n249) );
  OAI21X1 U367 ( .A(n947), .B(n171), .C(n250), .Y(n528) );
  OAI21X1 U368 ( .A(n25), .B(n964), .C(\mem<105> ), .Y(n250) );
  OAI21X1 U369 ( .A(n945), .B(n171), .C(n251), .Y(n529) );
  OAI21X1 U370 ( .A(n23), .B(n964), .C(\mem<104> ), .Y(n251) );
  OAI21X1 U371 ( .A(n944), .B(n171), .C(n252), .Y(n530) );
  OAI21X1 U372 ( .A(n21), .B(n964), .C(\mem<103> ), .Y(n252) );
  OAI21X1 U373 ( .A(n943), .B(n171), .C(n253), .Y(n531) );
  OAI21X1 U374 ( .A(n19), .B(n964), .C(\mem<102> ), .Y(n253) );
  OAI21X1 U375 ( .A(n942), .B(n171), .C(n254), .Y(n532) );
  OAI21X1 U376 ( .A(n17), .B(n964), .C(\mem<101> ), .Y(n254) );
  OAI21X1 U377 ( .A(n941), .B(n171), .C(n255), .Y(n533) );
  OAI21X1 U378 ( .A(n15), .B(n964), .C(\mem<100> ), .Y(n255) );
  OAI21X1 U379 ( .A(n940), .B(n171), .C(n256), .Y(n534) );
  OAI21X1 U380 ( .A(n13), .B(n964), .C(\mem<99> ), .Y(n256) );
  OAI21X1 U381 ( .A(n939), .B(n171), .C(n257), .Y(n535) );
  OAI21X1 U382 ( .A(n11), .B(n964), .C(\mem<98> ), .Y(n257) );
  OAI21X1 U383 ( .A(n938), .B(n171), .C(n258), .Y(n536) );
  OAI21X1 U384 ( .A(n9), .B(n964), .C(\mem<97> ), .Y(n258) );
  OAI21X1 U385 ( .A(n936), .B(n171), .C(n259), .Y(n537) );
  OAI21X1 U386 ( .A(n7), .B(n964), .C(\mem<96> ), .Y(n259) );
  OAI21X1 U389 ( .A(n957), .B(n152), .C(n261), .Y(n538) );
  OAI21X1 U390 ( .A(n37), .B(n963), .C(\mem<95> ), .Y(n261) );
  OAI21X1 U391 ( .A(n955), .B(n152), .C(n263), .Y(n539) );
  OAI21X1 U392 ( .A(n35), .B(n963), .C(\mem<94> ), .Y(n263) );
  OAI21X1 U393 ( .A(n954), .B(n152), .C(n264), .Y(n540) );
  OAI21X1 U394 ( .A(n33), .B(n963), .C(\mem<93> ), .Y(n264) );
  OAI21X1 U395 ( .A(n953), .B(n152), .C(n265), .Y(n541) );
  OAI21X1 U396 ( .A(n31), .B(n963), .C(\mem<92> ), .Y(n265) );
  OAI21X1 U397 ( .A(n951), .B(n152), .C(n266), .Y(n542) );
  OAI21X1 U398 ( .A(n29), .B(n963), .C(\mem<91> ), .Y(n266) );
  OAI21X1 U399 ( .A(n949), .B(n152), .C(n267), .Y(n543) );
  OAI21X1 U400 ( .A(n27), .B(n963), .C(\mem<90> ), .Y(n267) );
  OAI21X1 U401 ( .A(n947), .B(n152), .C(n268), .Y(n544) );
  OAI21X1 U402 ( .A(n25), .B(n963), .C(\mem<89> ), .Y(n268) );
  OAI21X1 U403 ( .A(n945), .B(n152), .C(n269), .Y(n545) );
  OAI21X1 U404 ( .A(n23), .B(n963), .C(\mem<88> ), .Y(n269) );
  OAI21X1 U405 ( .A(n944), .B(n152), .C(n270), .Y(n546) );
  OAI21X1 U406 ( .A(n21), .B(n963), .C(\mem<87> ), .Y(n270) );
  OAI21X1 U407 ( .A(n943), .B(n152), .C(n271), .Y(n547) );
  OAI21X1 U408 ( .A(n19), .B(n963), .C(\mem<86> ), .Y(n271) );
  OAI21X1 U409 ( .A(n942), .B(n152), .C(n272), .Y(n548) );
  OAI21X1 U410 ( .A(n17), .B(n963), .C(\mem<85> ), .Y(n272) );
  OAI21X1 U411 ( .A(n941), .B(n152), .C(n273), .Y(n549) );
  OAI21X1 U412 ( .A(n15), .B(n963), .C(\mem<84> ), .Y(n273) );
  OAI21X1 U413 ( .A(n940), .B(n152), .C(n274), .Y(n550) );
  OAI21X1 U414 ( .A(n13), .B(n963), .C(\mem<83> ), .Y(n274) );
  OAI21X1 U415 ( .A(n939), .B(n152), .C(n275), .Y(n551) );
  OAI21X1 U416 ( .A(n11), .B(n963), .C(\mem<82> ), .Y(n275) );
  OAI21X1 U417 ( .A(n938), .B(n152), .C(n276), .Y(n552) );
  OAI21X1 U418 ( .A(n9), .B(n963), .C(\mem<81> ), .Y(n276) );
  OAI21X1 U419 ( .A(n936), .B(n152), .C(n277), .Y(n553) );
  OAI21X1 U420 ( .A(n7), .B(n963), .C(\mem<80> ), .Y(n277) );
  OAI21X1 U423 ( .A(n957), .B(n149), .C(n279), .Y(n554) );
  OAI21X1 U424 ( .A(n37), .B(n962), .C(\mem<79> ), .Y(n279) );
  OAI21X1 U425 ( .A(n955), .B(n149), .C(n281), .Y(n555) );
  OAI21X1 U426 ( .A(n35), .B(n962), .C(\mem<78> ), .Y(n281) );
  OAI21X1 U427 ( .A(n954), .B(n149), .C(n282), .Y(n556) );
  OAI21X1 U428 ( .A(n33), .B(n962), .C(\mem<77> ), .Y(n282) );
  OAI21X1 U429 ( .A(n953), .B(n149), .C(n283), .Y(n557) );
  OAI21X1 U430 ( .A(n31), .B(n962), .C(\mem<76> ), .Y(n283) );
  OAI21X1 U431 ( .A(n951), .B(n149), .C(n284), .Y(n558) );
  OAI21X1 U432 ( .A(n29), .B(n962), .C(\mem<75> ), .Y(n284) );
  OAI21X1 U433 ( .A(n949), .B(n149), .C(n285), .Y(n559) );
  OAI21X1 U434 ( .A(n27), .B(n962), .C(\mem<74> ), .Y(n285) );
  OAI21X1 U435 ( .A(n947), .B(n149), .C(n286), .Y(n560) );
  OAI21X1 U436 ( .A(n25), .B(n962), .C(\mem<73> ), .Y(n286) );
  OAI21X1 U437 ( .A(n945), .B(n149), .C(n287), .Y(n561) );
  OAI21X1 U438 ( .A(n23), .B(n962), .C(\mem<72> ), .Y(n287) );
  OAI21X1 U439 ( .A(n944), .B(n149), .C(n288), .Y(n562) );
  OAI21X1 U440 ( .A(n21), .B(n962), .C(\mem<71> ), .Y(n288) );
  OAI21X1 U441 ( .A(n943), .B(n149), .C(n289), .Y(n563) );
  OAI21X1 U442 ( .A(n19), .B(n962), .C(\mem<70> ), .Y(n289) );
  OAI21X1 U443 ( .A(n942), .B(n149), .C(n290), .Y(n564) );
  OAI21X1 U444 ( .A(n17), .B(n962), .C(\mem<69> ), .Y(n290) );
  OAI21X1 U445 ( .A(n941), .B(n149), .C(n291), .Y(n565) );
  OAI21X1 U446 ( .A(n15), .B(n962), .C(\mem<68> ), .Y(n291) );
  OAI21X1 U447 ( .A(n940), .B(n149), .C(n292), .Y(n566) );
  OAI21X1 U448 ( .A(n13), .B(n962), .C(\mem<67> ), .Y(n292) );
  OAI21X1 U449 ( .A(n939), .B(n149), .C(n293), .Y(n567) );
  OAI21X1 U450 ( .A(n11), .B(n962), .C(\mem<66> ), .Y(n293) );
  OAI21X1 U451 ( .A(n938), .B(n149), .C(n294), .Y(n568) );
  OAI21X1 U452 ( .A(n9), .B(n962), .C(\mem<65> ), .Y(n294) );
  OAI21X1 U453 ( .A(n936), .B(n149), .C(n295), .Y(n569) );
  OAI21X1 U454 ( .A(n7), .B(n962), .C(\mem<64> ), .Y(n295) );
  OAI21X1 U458 ( .A(n957), .B(n131), .C(n297), .Y(n570) );
  OAI21X1 U459 ( .A(n37), .B(n961), .C(\mem<63> ), .Y(n297) );
  OAI21X1 U460 ( .A(n955), .B(n131), .C(n299), .Y(n571) );
  OAI21X1 U461 ( .A(n35), .B(n961), .C(\mem<62> ), .Y(n299) );
  OAI21X1 U462 ( .A(n954), .B(n131), .C(n300), .Y(n572) );
  OAI21X1 U463 ( .A(n33), .B(n961), .C(\mem<61> ), .Y(n300) );
  OAI21X1 U464 ( .A(n953), .B(n131), .C(n301), .Y(n573) );
  OAI21X1 U465 ( .A(n31), .B(n961), .C(\mem<60> ), .Y(n301) );
  OAI21X1 U466 ( .A(n951), .B(n131), .C(n302), .Y(n574) );
  OAI21X1 U467 ( .A(n29), .B(n961), .C(\mem<59> ), .Y(n302) );
  OAI21X1 U468 ( .A(n949), .B(n131), .C(n303), .Y(n575) );
  OAI21X1 U469 ( .A(n27), .B(n961), .C(\mem<58> ), .Y(n303) );
  OAI21X1 U470 ( .A(n947), .B(n131), .C(n304), .Y(n576) );
  OAI21X1 U471 ( .A(n25), .B(n961), .C(\mem<57> ), .Y(n304) );
  OAI21X1 U472 ( .A(n945), .B(n131), .C(n305), .Y(n577) );
  OAI21X1 U473 ( .A(n23), .B(n961), .C(\mem<56> ), .Y(n305) );
  OAI21X1 U474 ( .A(n944), .B(n131), .C(n306), .Y(n578) );
  OAI21X1 U475 ( .A(n21), .B(n961), .C(\mem<55> ), .Y(n306) );
  OAI21X1 U476 ( .A(n943), .B(n131), .C(n307), .Y(n579) );
  OAI21X1 U477 ( .A(n19), .B(n961), .C(\mem<54> ), .Y(n307) );
  OAI21X1 U478 ( .A(n942), .B(n131), .C(n308), .Y(n580) );
  OAI21X1 U479 ( .A(n17), .B(n961), .C(\mem<53> ), .Y(n308) );
  OAI21X1 U480 ( .A(n941), .B(n131), .C(n309), .Y(n581) );
  OAI21X1 U481 ( .A(n15), .B(n961), .C(\mem<52> ), .Y(n309) );
  OAI21X1 U482 ( .A(n940), .B(n131), .C(n310), .Y(n582) );
  OAI21X1 U483 ( .A(n13), .B(n961), .C(\mem<51> ), .Y(n310) );
  OAI21X1 U484 ( .A(n939), .B(n131), .C(n311), .Y(n583) );
  OAI21X1 U485 ( .A(n11), .B(n961), .C(\mem<50> ), .Y(n311) );
  OAI21X1 U486 ( .A(n938), .B(n131), .C(n312), .Y(n584) );
  OAI21X1 U487 ( .A(n9), .B(n961), .C(\mem<49> ), .Y(n312) );
  OAI21X1 U488 ( .A(n936), .B(n131), .C(n313), .Y(n585) );
  OAI21X1 U489 ( .A(n7), .B(n961), .C(\mem<48> ), .Y(n313) );
  OAI21X1 U492 ( .A(n957), .B(n114), .C(n316), .Y(n586) );
  OAI21X1 U493 ( .A(n37), .B(n960), .C(\mem<47> ), .Y(n316) );
  OAI21X1 U494 ( .A(n955), .B(n114), .C(n318), .Y(n587) );
  OAI21X1 U495 ( .A(n35), .B(n960), .C(\mem<46> ), .Y(n318) );
  OAI21X1 U496 ( .A(n954), .B(n114), .C(n319), .Y(n588) );
  OAI21X1 U497 ( .A(n33), .B(n960), .C(\mem<45> ), .Y(n319) );
  OAI21X1 U498 ( .A(n953), .B(n114), .C(n320), .Y(n589) );
  OAI21X1 U499 ( .A(n31), .B(n960), .C(\mem<44> ), .Y(n320) );
  OAI21X1 U500 ( .A(n951), .B(n114), .C(n321), .Y(n590) );
  OAI21X1 U501 ( .A(n29), .B(n960), .C(\mem<43> ), .Y(n321) );
  OAI21X1 U502 ( .A(n949), .B(n114), .C(n322), .Y(n591) );
  OAI21X1 U503 ( .A(n27), .B(n960), .C(\mem<42> ), .Y(n322) );
  OAI21X1 U504 ( .A(n947), .B(n114), .C(n323), .Y(n592) );
  OAI21X1 U505 ( .A(n25), .B(n960), .C(\mem<41> ), .Y(n323) );
  OAI21X1 U506 ( .A(n945), .B(n114), .C(n324), .Y(n593) );
  OAI21X1 U507 ( .A(n23), .B(n960), .C(\mem<40> ), .Y(n324) );
  OAI21X1 U508 ( .A(n944), .B(n114), .C(n325), .Y(n594) );
  OAI21X1 U509 ( .A(n21), .B(n960), .C(\mem<39> ), .Y(n325) );
  OAI21X1 U510 ( .A(n943), .B(n114), .C(n326), .Y(n595) );
  OAI21X1 U511 ( .A(n19), .B(n960), .C(\mem<38> ), .Y(n326) );
  OAI21X1 U512 ( .A(n942), .B(n114), .C(n327), .Y(n596) );
  OAI21X1 U513 ( .A(n17), .B(n960), .C(\mem<37> ), .Y(n327) );
  OAI21X1 U514 ( .A(n941), .B(n114), .C(n328), .Y(n597) );
  OAI21X1 U515 ( .A(n15), .B(n960), .C(\mem<36> ), .Y(n328) );
  OAI21X1 U516 ( .A(n940), .B(n114), .C(n329), .Y(n598) );
  OAI21X1 U517 ( .A(n13), .B(n960), .C(\mem<35> ), .Y(n329) );
  OAI21X1 U518 ( .A(n939), .B(n114), .C(n330), .Y(n599) );
  OAI21X1 U519 ( .A(n11), .B(n960), .C(\mem<34> ), .Y(n330) );
  OAI21X1 U520 ( .A(n938), .B(n114), .C(n331), .Y(n600) );
  OAI21X1 U521 ( .A(n9), .B(n960), .C(\mem<33> ), .Y(n331) );
  OAI21X1 U522 ( .A(n936), .B(n114), .C(n332), .Y(n601) );
  OAI21X1 U523 ( .A(n7), .B(n960), .C(\mem<32> ), .Y(n332) );
  OAI21X1 U526 ( .A(n957), .B(n95), .C(n334), .Y(n602) );
  OAI21X1 U527 ( .A(n37), .B(n959), .C(\mem<31> ), .Y(n334) );
  OAI21X1 U528 ( .A(n955), .B(n95), .C(n336), .Y(n603) );
  OAI21X1 U529 ( .A(n35), .B(n959), .C(\mem<30> ), .Y(n336) );
  OAI21X1 U530 ( .A(n954), .B(n95), .C(n337), .Y(n604) );
  OAI21X1 U531 ( .A(n33), .B(n959), .C(\mem<29> ), .Y(n337) );
  OAI21X1 U532 ( .A(n953), .B(n95), .C(n338), .Y(n605) );
  OAI21X1 U533 ( .A(n31), .B(n959), .C(\mem<28> ), .Y(n338) );
  OAI21X1 U534 ( .A(n951), .B(n95), .C(n339), .Y(n606) );
  OAI21X1 U535 ( .A(n29), .B(n959), .C(\mem<27> ), .Y(n339) );
  OAI21X1 U536 ( .A(n949), .B(n95), .C(n340), .Y(n607) );
  OAI21X1 U537 ( .A(n27), .B(n959), .C(\mem<26> ), .Y(n340) );
  OAI21X1 U538 ( .A(n947), .B(n95), .C(n341), .Y(n608) );
  OAI21X1 U539 ( .A(n25), .B(n959), .C(\mem<25> ), .Y(n341) );
  OAI21X1 U540 ( .A(n945), .B(n95), .C(n342), .Y(n609) );
  OAI21X1 U541 ( .A(n23), .B(n959), .C(\mem<24> ), .Y(n342) );
  OAI21X1 U542 ( .A(n944), .B(n95), .C(n343), .Y(n610) );
  OAI21X1 U543 ( .A(n21), .B(n959), .C(\mem<23> ), .Y(n343) );
  OAI21X1 U544 ( .A(n943), .B(n95), .C(n344), .Y(n611) );
  OAI21X1 U545 ( .A(n19), .B(n959), .C(\mem<22> ), .Y(n344) );
  OAI21X1 U546 ( .A(n942), .B(n95), .C(n345), .Y(n612) );
  OAI21X1 U547 ( .A(n17), .B(n959), .C(\mem<21> ), .Y(n345) );
  OAI21X1 U548 ( .A(n941), .B(n95), .C(n346), .Y(n613) );
  OAI21X1 U549 ( .A(n15), .B(n959), .C(\mem<20> ), .Y(n346) );
  OAI21X1 U550 ( .A(n940), .B(n95), .C(n347), .Y(n614) );
  OAI21X1 U551 ( .A(n13), .B(n959), .C(\mem<19> ), .Y(n347) );
  OAI21X1 U552 ( .A(n939), .B(n95), .C(n348), .Y(n615) );
  OAI21X1 U553 ( .A(n11), .B(n959), .C(\mem<18> ), .Y(n348) );
  OAI21X1 U554 ( .A(n938), .B(n95), .C(n349), .Y(n616) );
  OAI21X1 U555 ( .A(n9), .B(n959), .C(\mem<17> ), .Y(n349) );
  OAI21X1 U556 ( .A(n936), .B(n95), .C(n350), .Y(n617) );
  OAI21X1 U557 ( .A(n7), .B(n959), .C(\mem<16> ), .Y(n350) );
  OAI21X1 U561 ( .A(n957), .B(n71), .C(n352), .Y(n618) );
  OAI21X1 U562 ( .A(n37), .B(n937), .C(\mem<15> ), .Y(n352) );
  OAI21X1 U565 ( .A(n955), .B(n71), .C(n357), .Y(n619) );
  OAI21X1 U566 ( .A(n35), .B(n937), .C(\mem<14> ), .Y(n357) );
  OAI21X1 U569 ( .A(n954), .B(n71), .C(n359), .Y(n620) );
  OAI21X1 U570 ( .A(n33), .B(n937), .C(\mem<13> ), .Y(n359) );
  OAI21X1 U573 ( .A(n953), .B(n71), .C(n361), .Y(n621) );
  OAI21X1 U574 ( .A(n31), .B(n937), .C(\mem<12> ), .Y(n361) );
  OAI21X1 U577 ( .A(n951), .B(n71), .C(n363), .Y(n622) );
  OAI21X1 U578 ( .A(n29), .B(n937), .C(\mem<11> ), .Y(n363) );
  OAI21X1 U581 ( .A(n949), .B(n71), .C(n365), .Y(n623) );
  OAI21X1 U582 ( .A(n27), .B(n937), .C(\mem<10> ), .Y(n365) );
  OAI21X1 U585 ( .A(n947), .B(n71), .C(n366), .Y(n624) );
  OAI21X1 U586 ( .A(n25), .B(n937), .C(\mem<9> ), .Y(n366) );
  OAI21X1 U589 ( .A(n945), .B(n71), .C(n367), .Y(n625) );
  OAI21X1 U590 ( .A(n23), .B(n937), .C(\mem<8> ), .Y(n367) );
  OAI21X1 U593 ( .A(n944), .B(n71), .C(n368), .Y(n626) );
  OAI21X1 U594 ( .A(n21), .B(n937), .C(\mem<7> ), .Y(n368) );
  OAI21X1 U597 ( .A(n943), .B(n71), .C(n370), .Y(n627) );
  OAI21X1 U598 ( .A(n19), .B(n937), .C(\mem<6> ), .Y(n370) );
  OAI21X1 U601 ( .A(n942), .B(n71), .C(n371), .Y(n628) );
  OAI21X1 U602 ( .A(n17), .B(n937), .C(\mem<5> ), .Y(n371) );
  OAI21X1 U605 ( .A(n941), .B(n71), .C(n372), .Y(n629) );
  OAI21X1 U606 ( .A(n15), .B(n937), .C(\mem<4> ), .Y(n372) );
  OAI21X1 U610 ( .A(n940), .B(n71), .C(n373), .Y(n630) );
  OAI21X1 U611 ( .A(n13), .B(n937), .C(\mem<3> ), .Y(n373) );
  OAI21X1 U614 ( .A(n939), .B(n71), .C(n375), .Y(n631) );
  OAI21X1 U615 ( .A(n11), .B(n937), .C(\mem<2> ), .Y(n375) );
  OAI21X1 U618 ( .A(n938), .B(n71), .C(n376), .Y(n632) );
  OAI21X1 U619 ( .A(n9), .B(n937), .C(\mem<1> ), .Y(n376) );
  OAI21X1 U623 ( .A(n936), .B(n71), .C(n377), .Y(n633) );
  OAI21X1 U624 ( .A(n7), .B(n937), .C(\mem<0> ), .Y(n377) );
  NOR3X1 U634 ( .A(rst), .B(write), .C(n988), .Y(data_out) );
  INVX2 U2 ( .A(n66), .Y(n68) );
  INVX2 U3 ( .A(n187), .Y(n189) );
  INVX2 U4 ( .A(N21), .Y(n907) );
  INVX2 U5 ( .A(n907), .Y(n908) );
  AND2X1 U11 ( .A(N25), .B(n986), .Y(n168) );
  INVX1 U12 ( .A(N22), .Y(n985) );
  AND2X1 U13 ( .A(N25), .B(N24), .Y(n91) );
  AND2X1 U14 ( .A(N23), .B(n984), .Y(n92) );
  AND2X1 U15 ( .A(N23), .B(n985), .Y(n111) );
  BUFX2 U16 ( .A(n634), .Y(n978) );
  BUFX2 U17 ( .A(n360), .Y(n976) );
  BUFX2 U18 ( .A(n314), .Y(n972) );
  BUFX2 U19 ( .A(n278), .Y(n970) );
  BUFX2 U20 ( .A(n242), .Y(n968) );
  BUFX2 U21 ( .A(n207), .Y(n966) );
  BUFX2 U22 ( .A(n89), .Y(n957) );
  BUFX2 U23 ( .A(n86), .Y(n955) );
  BUFX2 U24 ( .A(n83), .Y(n951) );
  BUFX2 U25 ( .A(n80), .Y(n949) );
  BUFX2 U26 ( .A(n77), .Y(n947) );
  BUFX2 U27 ( .A(n74), .Y(n945) );
  INVX4 U28 ( .A(n981), .Y(n980) );
  INVX2 U29 ( .A(n985), .Y(n984) );
  INVX4 U30 ( .A(N18), .Y(n933) );
  INVX4 U31 ( .A(n933), .Y(n930) );
  INVX1 U32 ( .A(n39), .Y(n937) );
  INVX1 U33 ( .A(n53), .Y(n959) );
  INVX1 U34 ( .A(n54), .Y(n960) );
  INVX1 U35 ( .A(n56), .Y(n961) );
  INVX1 U36 ( .A(n57), .Y(n962) );
  INVX1 U37 ( .A(n59), .Y(n963) );
  INVX1 U38 ( .A(n60), .Y(n964) );
  INVX1 U39 ( .A(n62), .Y(n965) );
  INVX1 U40 ( .A(n63), .Y(n974) );
  INVX1 U41 ( .A(n65), .Y(n975) );
  BUFX2 U42 ( .A(n83), .Y(n952) );
  BUFX2 U43 ( .A(n89), .Y(n958) );
  BUFX2 U44 ( .A(n86), .Y(n956) );
  BUFX2 U45 ( .A(n74), .Y(n946) );
  BUFX2 U46 ( .A(n207), .Y(n967) );
  BUFX2 U47 ( .A(n242), .Y(n969) );
  BUFX2 U48 ( .A(n278), .Y(n971) );
  BUFX2 U81 ( .A(n314), .Y(n973) );
  BUFX2 U82 ( .A(n360), .Y(n977) );
  BUFX2 U115 ( .A(n634), .Y(n979) );
  BUFX2 U116 ( .A(n77), .Y(n948) );
  BUFX2 U149 ( .A(n80), .Y(n950) );
  INVX1 U150 ( .A(n38), .Y(n936) );
  INVX1 U183 ( .A(n40), .Y(n938) );
  INVX1 U184 ( .A(n41), .Y(n939) );
  INVX1 U217 ( .A(n43), .Y(n940) );
  INVX1 U218 ( .A(n44), .Y(n941) );
  INVX1 U251 ( .A(n45), .Y(n942) );
  INVX1 U252 ( .A(n47), .Y(n943) );
  INVX1 U285 ( .A(n48), .Y(n944) );
  INVX1 U286 ( .A(n50), .Y(n953) );
  INVX1 U319 ( .A(n51), .Y(n954) );
  INVX1 U320 ( .A(n983), .Y(n982) );
  INVX1 U353 ( .A(N24), .Y(n986) );
  AND2X2 U354 ( .A(n5), .B(n3), .Y(n1) );
  AND2X1 U387 ( .A(n817), .B(n980), .Y(n2) );
  INVX1 U388 ( .A(n2), .Y(n3) );
  AND2X1 U421 ( .A(n816), .B(n653), .Y(n4) );
  INVX1 U422 ( .A(n4), .Y(n5) );
  AND2X1 U455 ( .A(n38), .B(n68), .Y(n6) );
  INVX1 U456 ( .A(n6), .Y(n7) );
  AND2X1 U457 ( .A(n40), .B(n68), .Y(n8) );
  INVX1 U490 ( .A(n8), .Y(n9) );
  AND2X1 U491 ( .A(n41), .B(n68), .Y(n10) );
  INVX1 U524 ( .A(n10), .Y(n11) );
  AND2X1 U525 ( .A(n43), .B(n68), .Y(n12) );
  INVX1 U558 ( .A(n12), .Y(n13) );
  AND2X1 U559 ( .A(n44), .B(n68), .Y(n14) );
  INVX1 U560 ( .A(n14), .Y(n15) );
  AND2X1 U563 ( .A(n45), .B(n68), .Y(n16) );
  INVX1 U564 ( .A(n16), .Y(n17) );
  AND2X1 U567 ( .A(n47), .B(n68), .Y(n18) );
  INVX1 U568 ( .A(n18), .Y(n19) );
  AND2X1 U571 ( .A(n48), .B(n68), .Y(n20) );
  INVX1 U572 ( .A(n20), .Y(n21) );
  AND2X1 U575 ( .A(n72), .B(n68), .Y(n22) );
  INVX1 U576 ( .A(n22), .Y(n23) );
  AND2X1 U579 ( .A(n75), .B(n68), .Y(n24) );
  INVX1 U580 ( .A(n24), .Y(n25) );
  AND2X1 U583 ( .A(n78), .B(n68), .Y(n26) );
  INVX1 U584 ( .A(n26), .Y(n27) );
  AND2X1 U587 ( .A(n81), .B(n68), .Y(n28) );
  INVX1 U588 ( .A(n28), .Y(n29) );
  AND2X1 U591 ( .A(n50), .B(n68), .Y(n30) );
  INVX1 U592 ( .A(n30), .Y(n31) );
  AND2X1 U595 ( .A(n51), .B(n68), .Y(n32) );
  INVX1 U596 ( .A(n32), .Y(n33) );
  AND2X1 U599 ( .A(n84), .B(n68), .Y(n34) );
  INVX1 U600 ( .A(n34), .Y(n35) );
  AND2X1 U603 ( .A(n87), .B(n68), .Y(n36) );
  INVX1 U604 ( .A(n36), .Y(n37) );
  AND2X1 U607 ( .A(n646), .B(n638), .Y(n38) );
  AND2X1 U608 ( .A(n648), .B(n640), .Y(n39) );
  AND2X1 U609 ( .A(n646), .B(n642), .Y(n40) );
  AND2X1 U612 ( .A(n646), .B(n358), .Y(n41) );
  AND2X1 U613 ( .A(n646), .B(n356), .Y(n43) );
  AND2X1 U616 ( .A(n650), .B(n638), .Y(n44) );
  AND2X1 U617 ( .A(n650), .B(n642), .Y(n45) );
  AND2X1 U620 ( .A(n650), .B(n358), .Y(n47) );
  AND2X1 U621 ( .A(n650), .B(n356), .Y(n48) );
  AND2X1 U622 ( .A(n638), .B(n355), .Y(n50) );
  AND2X1 U625 ( .A(n642), .B(n355), .Y(n51) );
  AND2X1 U626 ( .A(n648), .B(n644), .Y(n53) );
  AND2X1 U627 ( .A(n648), .B(n111), .Y(n54) );
  AND2X1 U628 ( .A(n648), .B(n92), .Y(n56) );
  AND2X1 U629 ( .A(n652), .B(n640), .Y(n57) );
  AND2X1 U630 ( .A(n652), .B(n644), .Y(n59) );
  AND2X1 U631 ( .A(n652), .B(n111), .Y(n60) );
  AND2X1 U632 ( .A(n652), .B(n92), .Y(n62) );
  AND2X1 U633 ( .A(n640), .B(n91), .Y(n63) );
  AND2X1 U635 ( .A(n644), .B(n91), .Y(n65) );
  OR2X1 U636 ( .A(n987), .B(rst), .Y(n66) );
  AND2X1 U637 ( .A(n39), .B(n90), .Y(n69) );
  INVX1 U638 ( .A(n69), .Y(n71) );
  AND2X1 U639 ( .A(n364), .B(n638), .Y(n72) );
  INVX1 U640 ( .A(n72), .Y(n74) );
  AND2X1 U641 ( .A(n364), .B(n642), .Y(n75) );
  INVX1 U642 ( .A(n75), .Y(n77) );
  AND2X1 U643 ( .A(n364), .B(n358), .Y(n78) );
  INVX1 U644 ( .A(n78), .Y(n80) );
  AND2X1 U645 ( .A(n364), .B(n356), .Y(n81) );
  INVX1 U646 ( .A(n81), .Y(n83) );
  AND2X1 U647 ( .A(n358), .B(n355), .Y(n84) );
  INVX1 U648 ( .A(n84), .Y(n86) );
  AND2X1 U649 ( .A(n355), .B(n356), .Y(n87) );
  INVX1 U650 ( .A(n87), .Y(n89) );
  AND2X1 U651 ( .A(n53), .B(n90), .Y(n93) );
  INVX1 U652 ( .A(n93), .Y(n95) );
  AND2X1 U653 ( .A(n54), .B(n90), .Y(n112) );
  INVX1 U654 ( .A(n112), .Y(n114) );
  AND2X1 U655 ( .A(n56), .B(n90), .Y(n130) );
  INVX1 U656 ( .A(n130), .Y(n131) );
  AND2X1 U657 ( .A(n57), .B(n90), .Y(n133) );
  INVX1 U658 ( .A(n133), .Y(n149) );
  AND2X1 U659 ( .A(n59), .B(n90), .Y(n150) );
  INVX1 U660 ( .A(n150), .Y(n152) );
  AND2X1 U661 ( .A(n60), .B(n90), .Y(n169) );
  INVX1 U662 ( .A(n169), .Y(n171) );
  AND2X1 U663 ( .A(n62), .B(n90), .Y(n187) );
  AND2X1 U664 ( .A(n168), .B(n640), .Y(n205) );
  INVX1 U665 ( .A(n205), .Y(n207) );
  AND2X1 U666 ( .A(n205), .B(n90), .Y(n223) );
  INVX1 U667 ( .A(n223), .Y(n225) );
  AND2X1 U668 ( .A(n168), .B(n644), .Y(n241) );
  INVX1 U669 ( .A(n241), .Y(n242) );
  AND2X1 U670 ( .A(n241), .B(n90), .Y(n244) );
  INVX1 U671 ( .A(n244), .Y(n260) );
  AND2X1 U672 ( .A(n168), .B(n111), .Y(n262) );
  INVX1 U673 ( .A(n262), .Y(n278) );
  AND2X1 U674 ( .A(n262), .B(n90), .Y(n280) );
  INVX1 U675 ( .A(n280), .Y(n296) );
  AND2X1 U676 ( .A(n168), .B(n92), .Y(n298) );
  INVX1 U677 ( .A(n298), .Y(n314) );
  AND2X1 U678 ( .A(n298), .B(n90), .Y(n315) );
  INVX1 U679 ( .A(n315), .Y(n317) );
  AND2X1 U680 ( .A(n63), .B(n90), .Y(n333) );
  INVX1 U681 ( .A(n333), .Y(n335) );
  AND2X1 U682 ( .A(n65), .B(n90), .Y(n351) );
  INVX1 U683 ( .A(n351), .Y(n353) );
  AND2X1 U684 ( .A(n111), .B(n91), .Y(n354) );
  INVX1 U685 ( .A(n354), .Y(n360) );
  AND2X1 U686 ( .A(n354), .B(n90), .Y(n362) );
  INVX1 U687 ( .A(n362), .Y(n369) );
  AND2X1 U688 ( .A(n91), .B(n92), .Y(n374) );
  INVX1 U689 ( .A(n374), .Y(n634) );
  AND2X1 U690 ( .A(n90), .B(n374), .Y(n635) );
  INVX1 U691 ( .A(n635), .Y(n636) );
  OR2X1 U692 ( .A(N18), .B(n980), .Y(n637) );
  INVX1 U693 ( .A(n637), .Y(n638) );
  OR2X1 U694 ( .A(n984), .B(N23), .Y(n639) );
  INVX1 U695 ( .A(n639), .Y(n640) );
  OR2X1 U696 ( .A(n921), .B(n980), .Y(n641) );
  INVX1 U697 ( .A(n641), .Y(n642) );
  OR2X1 U698 ( .A(n985), .B(N23), .Y(n643) );
  INVX1 U699 ( .A(n643), .Y(n644) );
  OR2X1 U700 ( .A(n982), .B(N21), .Y(n645) );
  INVX1 U701 ( .A(n645), .Y(n646) );
  OR2X1 U702 ( .A(N24), .B(N25), .Y(n647) );
  INVX1 U703 ( .A(n647), .Y(n648) );
  OR2X1 U704 ( .A(n983), .B(N21), .Y(n649) );
  INVX1 U705 ( .A(n649), .Y(n650) );
  OR2X1 U706 ( .A(n986), .B(N25), .Y(n651) );
  INVX1 U707 ( .A(n651), .Y(n652) );
  INVX1 U708 ( .A(n980), .Y(n653) );
  INVX1 U709 ( .A(N28), .Y(n988) );
  MUX2X1 U710 ( .B(n655), .A(n656), .S(n919), .Y(n654) );
  MUX2X1 U711 ( .B(n658), .A(n659), .S(n919), .Y(n657) );
  MUX2X1 U712 ( .B(n661), .A(n662), .S(n919), .Y(n660) );
  MUX2X1 U713 ( .B(n664), .A(n665), .S(n919), .Y(n663) );
  MUX2X1 U714 ( .B(n667), .A(n668), .S(n909), .Y(n666) );
  MUX2X1 U715 ( .B(n670), .A(n671), .S(n919), .Y(n669) );
  MUX2X1 U716 ( .B(n673), .A(n674), .S(n919), .Y(n672) );
  MUX2X1 U717 ( .B(n676), .A(n677), .S(n919), .Y(n675) );
  MUX2X1 U718 ( .B(n679), .A(n680), .S(n919), .Y(n678) );
  MUX2X1 U719 ( .B(n682), .A(n683), .S(n909), .Y(n681) );
  MUX2X1 U720 ( .B(n685), .A(n686), .S(n919), .Y(n684) );
  MUX2X1 U721 ( .B(n688), .A(n689), .S(n919), .Y(n687) );
  MUX2X1 U722 ( .B(n691), .A(n692), .S(n919), .Y(n690) );
  MUX2X1 U723 ( .B(n694), .A(n695), .S(n919), .Y(n693) );
  MUX2X1 U724 ( .B(n697), .A(n698), .S(n909), .Y(n696) );
  MUX2X1 U725 ( .B(n700), .A(n701), .S(n918), .Y(n699) );
  MUX2X1 U726 ( .B(n703), .A(n704), .S(n918), .Y(n702) );
  MUX2X1 U727 ( .B(n706), .A(n707), .S(n918), .Y(n705) );
  MUX2X1 U728 ( .B(n709), .A(n710), .S(n918), .Y(n708) );
  MUX2X1 U729 ( .B(n712), .A(n713), .S(n909), .Y(n711) );
  MUX2X1 U730 ( .B(n715), .A(n716), .S(N23), .Y(n714) );
  MUX2X1 U731 ( .B(n718), .A(n719), .S(n918), .Y(n717) );
  MUX2X1 U732 ( .B(n721), .A(n722), .S(n918), .Y(n720) );
  MUX2X1 U733 ( .B(n724), .A(n725), .S(n918), .Y(n723) );
  MUX2X1 U734 ( .B(n727), .A(n728), .S(n918), .Y(n726) );
  MUX2X1 U735 ( .B(n730), .A(n731), .S(n909), .Y(n729) );
  MUX2X1 U736 ( .B(n733), .A(n734), .S(n918), .Y(n732) );
  MUX2X1 U737 ( .B(n736), .A(n737), .S(n918), .Y(n735) );
  MUX2X1 U738 ( .B(n739), .A(n740), .S(n918), .Y(n738) );
  MUX2X1 U739 ( .B(n742), .A(n743), .S(n918), .Y(n741) );
  MUX2X1 U740 ( .B(n745), .A(n746), .S(n909), .Y(n744) );
  MUX2X1 U741 ( .B(n748), .A(n749), .S(n917), .Y(n747) );
  MUX2X1 U742 ( .B(n751), .A(n752), .S(n917), .Y(n750) );
  MUX2X1 U743 ( .B(n754), .A(n755), .S(n917), .Y(n753) );
  MUX2X1 U744 ( .B(n757), .A(n758), .S(n917), .Y(n756) );
  MUX2X1 U745 ( .B(n760), .A(n761), .S(n909), .Y(n759) );
  MUX2X1 U746 ( .B(n763), .A(n764), .S(n917), .Y(n762) );
  MUX2X1 U747 ( .B(n766), .A(n767), .S(n917), .Y(n765) );
  MUX2X1 U748 ( .B(n769), .A(n770), .S(n917), .Y(n768) );
  MUX2X1 U749 ( .B(n772), .A(n773), .S(n917), .Y(n771) );
  MUX2X1 U750 ( .B(n775), .A(n776), .S(n909), .Y(n774) );
  MUX2X1 U751 ( .B(n778), .A(n779), .S(N23), .Y(n777) );
  MUX2X1 U752 ( .B(n781), .A(n782), .S(n917), .Y(n780) );
  MUX2X1 U753 ( .B(n784), .A(n785), .S(n917), .Y(n783) );
  MUX2X1 U754 ( .B(n787), .A(n788), .S(n917), .Y(n786) );
  MUX2X1 U755 ( .B(n790), .A(n791), .S(n917), .Y(n789) );
  MUX2X1 U756 ( .B(n793), .A(n794), .S(n909), .Y(n792) );
  MUX2X1 U757 ( .B(n796), .A(n797), .S(n917), .Y(n795) );
  MUX2X1 U758 ( .B(n799), .A(n800), .S(n915), .Y(n798) );
  MUX2X1 U759 ( .B(n802), .A(n803), .S(n915), .Y(n801) );
  MUX2X1 U760 ( .B(n805), .A(n806), .S(n918), .Y(n804) );
  MUX2X1 U761 ( .B(n808), .A(n809), .S(n909), .Y(n807) );
  MUX2X1 U762 ( .B(n811), .A(n812), .S(n915), .Y(n810) );
  MUX2X1 U763 ( .B(n814), .A(n815), .S(n918), .Y(n813) );
  MUX2X1 U764 ( .B(n819), .A(n820), .S(n915), .Y(n818) );
  MUX2X1 U765 ( .B(n822), .A(n823), .S(n909), .Y(n821) );
  MUX2X1 U766 ( .B(n825), .A(n826), .S(n915), .Y(n824) );
  MUX2X1 U767 ( .B(n828), .A(n829), .S(n919), .Y(n827) );
  MUX2X1 U768 ( .B(n831), .A(n832), .S(n915), .Y(n830) );
  MUX2X1 U769 ( .B(n834), .A(n835), .S(n915), .Y(n833) );
  MUX2X1 U770 ( .B(n837), .A(n838), .S(n909), .Y(n836) );
  MUX2X1 U771 ( .B(n840), .A(n841), .S(N23), .Y(n839) );
  MUX2X1 U772 ( .B(n843), .A(n844), .S(n916), .Y(n842) );
  MUX2X1 U773 ( .B(n846), .A(n847), .S(n916), .Y(n845) );
  MUX2X1 U774 ( .B(n849), .A(n850), .S(n916), .Y(n848) );
  MUX2X1 U775 ( .B(n852), .A(n853), .S(n916), .Y(n851) );
  MUX2X1 U776 ( .B(n855), .A(n856), .S(n908), .Y(n854) );
  MUX2X1 U777 ( .B(n858), .A(n859), .S(n916), .Y(n857) );
  MUX2X1 U778 ( .B(n861), .A(n862), .S(n916), .Y(n860) );
  MUX2X1 U779 ( .B(n864), .A(n865), .S(n916), .Y(n863) );
  MUX2X1 U780 ( .B(n867), .A(n868), .S(n916), .Y(n866) );
  MUX2X1 U781 ( .B(n870), .A(n871), .S(n908), .Y(n869) );
  MUX2X1 U782 ( .B(n873), .A(n874), .S(n916), .Y(n872) );
  MUX2X1 U783 ( .B(n876), .A(n877), .S(n916), .Y(n875) );
  MUX2X1 U784 ( .B(n879), .A(n880), .S(n916), .Y(n878) );
  MUX2X1 U785 ( .B(n882), .A(n883), .S(n916), .Y(n881) );
  MUX2X1 U786 ( .B(n885), .A(n886), .S(n908), .Y(n884) );
  MUX2X1 U787 ( .B(n888), .A(n889), .S(n915), .Y(n887) );
  MUX2X1 U788 ( .B(n891), .A(n892), .S(n915), .Y(n890) );
  MUX2X1 U789 ( .B(n894), .A(n895), .S(n915), .Y(n893) );
  MUX2X1 U790 ( .B(n897), .A(n898), .S(n915), .Y(n896) );
  MUX2X1 U791 ( .B(n900), .A(n901), .S(n908), .Y(n899) );
  MUX2X1 U792 ( .B(n903), .A(n904), .S(N23), .Y(n902) );
  MUX2X1 U793 ( .B(n905), .A(n906), .S(N25), .Y(N28) );
  MUX2X1 U794 ( .B(\mem<254> ), .A(\mem<255> ), .S(n923), .Y(n656) );
  MUX2X1 U795 ( .B(\mem<252> ), .A(\mem<253> ), .S(n923), .Y(n655) );
  MUX2X1 U796 ( .B(\mem<250> ), .A(\mem<251> ), .S(n923), .Y(n659) );
  MUX2X1 U797 ( .B(\mem<248> ), .A(\mem<249> ), .S(n923), .Y(n658) );
  MUX2X1 U798 ( .B(n657), .A(n654), .S(n912), .Y(n668) );
  MUX2X1 U799 ( .B(\mem<246> ), .A(\mem<247> ), .S(n923), .Y(n662) );
  MUX2X1 U800 ( .B(\mem<244> ), .A(\mem<245> ), .S(n923), .Y(n661) );
  MUX2X1 U801 ( .B(\mem<242> ), .A(\mem<243> ), .S(n923), .Y(n665) );
  MUX2X1 U802 ( .B(\mem<240> ), .A(\mem<241> ), .S(n923), .Y(n664) );
  MUX2X1 U803 ( .B(n663), .A(n660), .S(n912), .Y(n667) );
  MUX2X1 U804 ( .B(\mem<238> ), .A(\mem<239> ), .S(n924), .Y(n671) );
  MUX2X1 U805 ( .B(\mem<236> ), .A(\mem<237> ), .S(n924), .Y(n670) );
  MUX2X1 U806 ( .B(\mem<234> ), .A(\mem<235> ), .S(n924), .Y(n674) );
  MUX2X1 U807 ( .B(\mem<232> ), .A(\mem<233> ), .S(n924), .Y(n673) );
  MUX2X1 U808 ( .B(n672), .A(n669), .S(n912), .Y(n683) );
  MUX2X1 U809 ( .B(\mem<230> ), .A(\mem<231> ), .S(n924), .Y(n677) );
  MUX2X1 U810 ( .B(\mem<228> ), .A(\mem<229> ), .S(n924), .Y(n676) );
  MUX2X1 U811 ( .B(\mem<226> ), .A(\mem<227> ), .S(n924), .Y(n680) );
  MUX2X1 U812 ( .B(\mem<224> ), .A(\mem<225> ), .S(n924), .Y(n679) );
  MUX2X1 U813 ( .B(n678), .A(n675), .S(n912), .Y(n682) );
  MUX2X1 U814 ( .B(n681), .A(n666), .S(n984), .Y(n716) );
  MUX2X1 U815 ( .B(\mem<222> ), .A(\mem<223> ), .S(n924), .Y(n686) );
  MUX2X1 U816 ( .B(\mem<220> ), .A(\mem<221> ), .S(n924), .Y(n685) );
  MUX2X1 U817 ( .B(\mem<218> ), .A(\mem<219> ), .S(n924), .Y(n689) );
  MUX2X1 U818 ( .B(\mem<216> ), .A(\mem<217> ), .S(n924), .Y(n688) );
  MUX2X1 U819 ( .B(n687), .A(n684), .S(n912), .Y(n698) );
  MUX2X1 U820 ( .B(\mem<214> ), .A(\mem<215> ), .S(n925), .Y(n692) );
  MUX2X1 U821 ( .B(\mem<212> ), .A(\mem<213> ), .S(n925), .Y(n691) );
  MUX2X1 U822 ( .B(\mem<210> ), .A(\mem<211> ), .S(n925), .Y(n695) );
  MUX2X1 U823 ( .B(\mem<208> ), .A(\mem<209> ), .S(n925), .Y(n694) );
  MUX2X1 U824 ( .B(n693), .A(n690), .S(n912), .Y(n697) );
  MUX2X1 U825 ( .B(\mem<206> ), .A(\mem<207> ), .S(n925), .Y(n701) );
  MUX2X1 U826 ( .B(\mem<204> ), .A(\mem<205> ), .S(n925), .Y(n700) );
  MUX2X1 U827 ( .B(\mem<202> ), .A(\mem<203> ), .S(n925), .Y(n704) );
  MUX2X1 U828 ( .B(\mem<200> ), .A(\mem<201> ), .S(n925), .Y(n703) );
  MUX2X1 U829 ( .B(n702), .A(n699), .S(n912), .Y(n713) );
  MUX2X1 U830 ( .B(\mem<198> ), .A(\mem<199> ), .S(n925), .Y(n707) );
  MUX2X1 U831 ( .B(\mem<196> ), .A(\mem<197> ), .S(n925), .Y(n706) );
  MUX2X1 U832 ( .B(\mem<194> ), .A(\mem<195> ), .S(n925), .Y(n710) );
  MUX2X1 U833 ( .B(\mem<192> ), .A(\mem<193> ), .S(n925), .Y(n709) );
  MUX2X1 U834 ( .B(n708), .A(n705), .S(n912), .Y(n712) );
  MUX2X1 U835 ( .B(n711), .A(n696), .S(n984), .Y(n715) );
  MUX2X1 U836 ( .B(\mem<190> ), .A(\mem<191> ), .S(n926), .Y(n719) );
  MUX2X1 U837 ( .B(\mem<188> ), .A(\mem<189> ), .S(n926), .Y(n718) );
  MUX2X1 U838 ( .B(\mem<186> ), .A(\mem<187> ), .S(n926), .Y(n722) );
  MUX2X1 U839 ( .B(\mem<184> ), .A(\mem<185> ), .S(n926), .Y(n721) );
  MUX2X1 U840 ( .B(n720), .A(n717), .S(n912), .Y(n731) );
  MUX2X1 U841 ( .B(\mem<182> ), .A(\mem<183> ), .S(n926), .Y(n725) );
  MUX2X1 U842 ( .B(\mem<180> ), .A(\mem<181> ), .S(n926), .Y(n724) );
  MUX2X1 U843 ( .B(\mem<178> ), .A(\mem<179> ), .S(n926), .Y(n728) );
  MUX2X1 U844 ( .B(\mem<176> ), .A(\mem<177> ), .S(n926), .Y(n727) );
  MUX2X1 U845 ( .B(n726), .A(n723), .S(n912), .Y(n730) );
  MUX2X1 U846 ( .B(\mem<174> ), .A(\mem<175> ), .S(n926), .Y(n734) );
  MUX2X1 U847 ( .B(\mem<172> ), .A(\mem<173> ), .S(n926), .Y(n733) );
  MUX2X1 U848 ( .B(\mem<170> ), .A(\mem<171> ), .S(n926), .Y(n737) );
  MUX2X1 U849 ( .B(\mem<168> ), .A(\mem<169> ), .S(n926), .Y(n736) );
  MUX2X1 U850 ( .B(n735), .A(n732), .S(n912), .Y(n746) );
  MUX2X1 U851 ( .B(\mem<166> ), .A(\mem<167> ), .S(n927), .Y(n740) );
  MUX2X1 U852 ( .B(\mem<164> ), .A(\mem<165> ), .S(n927), .Y(n739) );
  MUX2X1 U853 ( .B(\mem<162> ), .A(\mem<163> ), .S(n927), .Y(n743) );
  MUX2X1 U854 ( .B(\mem<160> ), .A(\mem<161> ), .S(n927), .Y(n742) );
  MUX2X1 U855 ( .B(n741), .A(n738), .S(n912), .Y(n745) );
  MUX2X1 U856 ( .B(n744), .A(n729), .S(n984), .Y(n779) );
  MUX2X1 U857 ( .B(\mem<158> ), .A(\mem<159> ), .S(n927), .Y(n749) );
  MUX2X1 U858 ( .B(\mem<156> ), .A(\mem<157> ), .S(n927), .Y(n748) );
  MUX2X1 U859 ( .B(\mem<154> ), .A(\mem<155> ), .S(n927), .Y(n752) );
  MUX2X1 U860 ( .B(\mem<152> ), .A(\mem<153> ), .S(n927), .Y(n751) );
  MUX2X1 U861 ( .B(n750), .A(n747), .S(n911), .Y(n761) );
  MUX2X1 U862 ( .B(\mem<150> ), .A(\mem<151> ), .S(n927), .Y(n755) );
  MUX2X1 U863 ( .B(\mem<148> ), .A(\mem<149> ), .S(n927), .Y(n754) );
  MUX2X1 U864 ( .B(\mem<146> ), .A(\mem<147> ), .S(n927), .Y(n758) );
  MUX2X1 U865 ( .B(\mem<144> ), .A(\mem<145> ), .S(n927), .Y(n757) );
  MUX2X1 U866 ( .B(n756), .A(n753), .S(n911), .Y(n760) );
  MUX2X1 U867 ( .B(\mem<142> ), .A(\mem<143> ), .S(n928), .Y(n764) );
  MUX2X1 U868 ( .B(\mem<140> ), .A(\mem<141> ), .S(n928), .Y(n763) );
  MUX2X1 U869 ( .B(\mem<138> ), .A(\mem<139> ), .S(n928), .Y(n767) );
  MUX2X1 U870 ( .B(\mem<136> ), .A(\mem<137> ), .S(n928), .Y(n766) );
  MUX2X1 U871 ( .B(n765), .A(n762), .S(n911), .Y(n776) );
  MUX2X1 U872 ( .B(\mem<134> ), .A(\mem<135> ), .S(n928), .Y(n770) );
  MUX2X1 U873 ( .B(\mem<132> ), .A(\mem<133> ), .S(n928), .Y(n769) );
  MUX2X1 U874 ( .B(\mem<130> ), .A(\mem<131> ), .S(n928), .Y(n773) );
  MUX2X1 U875 ( .B(\mem<128> ), .A(\mem<129> ), .S(n928), .Y(n772) );
  MUX2X1 U876 ( .B(n771), .A(n768), .S(n911), .Y(n775) );
  MUX2X1 U877 ( .B(n774), .A(n759), .S(n984), .Y(n778) );
  MUX2X1 U878 ( .B(n777), .A(n714), .S(N24), .Y(n906) );
  MUX2X1 U879 ( .B(\mem<126> ), .A(\mem<127> ), .S(n928), .Y(n782) );
  MUX2X1 U880 ( .B(\mem<124> ), .A(\mem<125> ), .S(n928), .Y(n781) );
  MUX2X1 U881 ( .B(\mem<122> ), .A(\mem<123> ), .S(n928), .Y(n785) );
  MUX2X1 U882 ( .B(\mem<120> ), .A(\mem<121> ), .S(n928), .Y(n784) );
  MUX2X1 U883 ( .B(n783), .A(n780), .S(n911), .Y(n794) );
  MUX2X1 U884 ( .B(\mem<118> ), .A(\mem<119> ), .S(n929), .Y(n788) );
  MUX2X1 U885 ( .B(\mem<116> ), .A(\mem<117> ), .S(n929), .Y(n787) );
  MUX2X1 U886 ( .B(\mem<114> ), .A(\mem<115> ), .S(n929), .Y(n791) );
  MUX2X1 U887 ( .B(\mem<112> ), .A(\mem<113> ), .S(n929), .Y(n790) );
  MUX2X1 U888 ( .B(n789), .A(n786), .S(n911), .Y(n793) );
  MUX2X1 U889 ( .B(\mem<110> ), .A(\mem<111> ), .S(n929), .Y(n797) );
  MUX2X1 U890 ( .B(\mem<108> ), .A(\mem<109> ), .S(n929), .Y(n796) );
  MUX2X1 U891 ( .B(\mem<106> ), .A(\mem<107> ), .S(n929), .Y(n800) );
  MUX2X1 U892 ( .B(\mem<104> ), .A(\mem<105> ), .S(n929), .Y(n799) );
  MUX2X1 U893 ( .B(n798), .A(n795), .S(n911), .Y(n809) );
  MUX2X1 U894 ( .B(\mem<102> ), .A(\mem<103> ), .S(n929), .Y(n803) );
  MUX2X1 U895 ( .B(\mem<100> ), .A(\mem<101> ), .S(n929), .Y(n802) );
  MUX2X1 U896 ( .B(\mem<98> ), .A(\mem<99> ), .S(n929), .Y(n806) );
  MUX2X1 U897 ( .B(\mem<96> ), .A(\mem<97> ), .S(n929), .Y(n805) );
  MUX2X1 U898 ( .B(n804), .A(n801), .S(n911), .Y(n808) );
  MUX2X1 U899 ( .B(n807), .A(n792), .S(n984), .Y(n841) );
  MUX2X1 U900 ( .B(\mem<94> ), .A(\mem<95> ), .S(n930), .Y(n812) );
  MUX2X1 U901 ( .B(\mem<92> ), .A(\mem<93> ), .S(n930), .Y(n811) );
  MUX2X1 U902 ( .B(\mem<90> ), .A(\mem<91> ), .S(n930), .Y(n815) );
  MUX2X1 U903 ( .B(\mem<88> ), .A(\mem<89> ), .S(n930), .Y(n814) );
  MUX2X1 U904 ( .B(n813), .A(n810), .S(n911), .Y(n823) );
  MUX2X1 U905 ( .B(\mem<86> ), .A(\mem<87> ), .S(n930), .Y(n817) );
  MUX2X1 U906 ( .B(\mem<84> ), .A(\mem<85> ), .S(n930), .Y(n816) );
  MUX2X1 U907 ( .B(\mem<82> ), .A(\mem<83> ), .S(n930), .Y(n820) );
  MUX2X1 U908 ( .B(\mem<80> ), .A(\mem<81> ), .S(n930), .Y(n819) );
  MUX2X1 U909 ( .B(n818), .A(n1), .S(n911), .Y(n822) );
  MUX2X1 U910 ( .B(\mem<78> ), .A(\mem<79> ), .S(n930), .Y(n826) );
  MUX2X1 U911 ( .B(\mem<76> ), .A(\mem<77> ), .S(n930), .Y(n825) );
  MUX2X1 U912 ( .B(\mem<74> ), .A(\mem<75> ), .S(n930), .Y(n829) );
  MUX2X1 U913 ( .B(\mem<72> ), .A(\mem<73> ), .S(n930), .Y(n828) );
  MUX2X1 U914 ( .B(n827), .A(n824), .S(n911), .Y(n838) );
  MUX2X1 U915 ( .B(\mem<70> ), .A(\mem<71> ), .S(n929), .Y(n832) );
  MUX2X1 U916 ( .B(\mem<68> ), .A(\mem<69> ), .S(n929), .Y(n831) );
  MUX2X1 U917 ( .B(\mem<66> ), .A(\mem<67> ), .S(n929), .Y(n835) );
  MUX2X1 U918 ( .B(\mem<64> ), .A(\mem<65> ), .S(n929), .Y(n834) );
  MUX2X1 U919 ( .B(n833), .A(n830), .S(n911), .Y(n837) );
  MUX2X1 U920 ( .B(n836), .A(n821), .S(n984), .Y(n840) );
  MUX2X1 U921 ( .B(\mem<62> ), .A(\mem<63> ), .S(n930), .Y(n844) );
  MUX2X1 U922 ( .B(\mem<60> ), .A(\mem<61> ), .S(n929), .Y(n843) );
  MUX2X1 U923 ( .B(\mem<58> ), .A(\mem<59> ), .S(n929), .Y(n847) );
  MUX2X1 U924 ( .B(\mem<56> ), .A(\mem<57> ), .S(n930), .Y(n846) );
  MUX2X1 U925 ( .B(n845), .A(n842), .S(n910), .Y(n856) );
  MUX2X1 U926 ( .B(\mem<54> ), .A(\mem<55> ), .S(n929), .Y(n850) );
  MUX2X1 U927 ( .B(\mem<52> ), .A(\mem<53> ), .S(n929), .Y(n849) );
  MUX2X1 U928 ( .B(\mem<50> ), .A(\mem<51> ), .S(n929), .Y(n853) );
  MUX2X1 U929 ( .B(\mem<48> ), .A(\mem<49> ), .S(n929), .Y(n852) );
  MUX2X1 U930 ( .B(n851), .A(n848), .S(n910), .Y(n855) );
  MUX2X1 U931 ( .B(\mem<46> ), .A(\mem<47> ), .S(n931), .Y(n859) );
  MUX2X1 U932 ( .B(\mem<44> ), .A(\mem<45> ), .S(n931), .Y(n858) );
  MUX2X1 U933 ( .B(\mem<42> ), .A(\mem<43> ), .S(n931), .Y(n862) );
  MUX2X1 U934 ( .B(\mem<40> ), .A(\mem<41> ), .S(n931), .Y(n861) );
  MUX2X1 U935 ( .B(n860), .A(n857), .S(n910), .Y(n871) );
  MUX2X1 U936 ( .B(\mem<38> ), .A(\mem<39> ), .S(n931), .Y(n865) );
  MUX2X1 U937 ( .B(\mem<36> ), .A(\mem<37> ), .S(n931), .Y(n864) );
  MUX2X1 U938 ( .B(\mem<34> ), .A(\mem<35> ), .S(n931), .Y(n868) );
  MUX2X1 U939 ( .B(\mem<32> ), .A(\mem<33> ), .S(n931), .Y(n867) );
  MUX2X1 U940 ( .B(n866), .A(n863), .S(n910), .Y(n870) );
  MUX2X1 U941 ( .B(n869), .A(n854), .S(n984), .Y(n904) );
  MUX2X1 U942 ( .B(\mem<30> ), .A(\mem<31> ), .S(n931), .Y(n874) );
  MUX2X1 U943 ( .B(\mem<28> ), .A(\mem<29> ), .S(n931), .Y(n873) );
  MUX2X1 U944 ( .B(\mem<26> ), .A(\mem<27> ), .S(n931), .Y(n877) );
  MUX2X1 U945 ( .B(\mem<24> ), .A(\mem<25> ), .S(n931), .Y(n876) );
  MUX2X1 U946 ( .B(n875), .A(n872), .S(n910), .Y(n886) );
  MUX2X1 U947 ( .B(\mem<22> ), .A(\mem<23> ), .S(n932), .Y(n880) );
  MUX2X1 U948 ( .B(\mem<20> ), .A(\mem<21> ), .S(n932), .Y(n879) );
  MUX2X1 U949 ( .B(\mem<18> ), .A(\mem<19> ), .S(n932), .Y(n883) );
  MUX2X1 U950 ( .B(\mem<16> ), .A(\mem<17> ), .S(n932), .Y(n882) );
  MUX2X1 U951 ( .B(n881), .A(n878), .S(n910), .Y(n885) );
  MUX2X1 U952 ( .B(\mem<14> ), .A(\mem<15> ), .S(n932), .Y(n889) );
  MUX2X1 U953 ( .B(\mem<12> ), .A(\mem<13> ), .S(n932), .Y(n888) );
  MUX2X1 U954 ( .B(\mem<10> ), .A(\mem<11> ), .S(n932), .Y(n892) );
  MUX2X1 U955 ( .B(\mem<8> ), .A(\mem<9> ), .S(n932), .Y(n891) );
  MUX2X1 U956 ( .B(n890), .A(n887), .S(n910), .Y(n901) );
  MUX2X1 U957 ( .B(\mem<6> ), .A(\mem<7> ), .S(n932), .Y(n895) );
  MUX2X1 U958 ( .B(\mem<4> ), .A(\mem<5> ), .S(n932), .Y(n894) );
  MUX2X1 U959 ( .B(\mem<2> ), .A(\mem<3> ), .S(n932), .Y(n898) );
  MUX2X1 U960 ( .B(\mem<0> ), .A(\mem<1> ), .S(n932), .Y(n897) );
  MUX2X1 U961 ( .B(n896), .A(n893), .S(n910), .Y(n900) );
  MUX2X1 U962 ( .B(n899), .A(n884), .S(n984), .Y(n903) );
  MUX2X1 U963 ( .B(n902), .A(n839), .S(N24), .Y(n905) );
  INVX8 U964 ( .A(n907), .Y(n909) );
  INVX8 U965 ( .A(n983), .Y(n910) );
  INVX8 U966 ( .A(n983), .Y(n911) );
  INVX8 U967 ( .A(n983), .Y(n912) );
  INVX8 U968 ( .A(n980), .Y(n913) );
  INVX8 U969 ( .A(n980), .Y(n914) );
  INVX8 U970 ( .A(n914), .Y(n915) );
  INVX8 U971 ( .A(n914), .Y(n916) );
  INVX8 U972 ( .A(n913), .Y(n917) );
  INVX8 U973 ( .A(n913), .Y(n918) );
  INVX8 U974 ( .A(n913), .Y(n919) );
  INVX8 U975 ( .A(n934), .Y(n920) );
  INVX8 U976 ( .A(n935), .Y(n921) );
  INVX8 U977 ( .A(n935), .Y(n922) );
  INVX8 U978 ( .A(n922), .Y(n923) );
  INVX8 U979 ( .A(n922), .Y(n924) );
  INVX8 U980 ( .A(n922), .Y(n925) );
  INVX8 U981 ( .A(n921), .Y(n926) );
  INVX8 U982 ( .A(n921), .Y(n927) );
  INVX8 U983 ( .A(n921), .Y(n928) );
  INVX8 U984 ( .A(n933), .Y(n929) );
  INVX8 U985 ( .A(n920), .Y(n931) );
  INVX8 U986 ( .A(n920), .Y(n932) );
  INVX8 U987 ( .A(n933), .Y(n934) );
  INVX8 U988 ( .A(n933), .Y(n935) );
  INVX1 U989 ( .A(N19), .Y(n981) );
  INVX1 U990 ( .A(write), .Y(n987) );
  INVX8 U991 ( .A(N20), .Y(n983) );
endmodule


module memc_Size16_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1926), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1927), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1928), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1929), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1930), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1931), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1932), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1933), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1934), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1935), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1936), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1937), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1938), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1939), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1940), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1941), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1942), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1943), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1944), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1945), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1946), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1947), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1948), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1949), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1950), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1951), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1952), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1953), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1954), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1955), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1956), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1957), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1958), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1959), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1960), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1961), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1962), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1963), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1964), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1965), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1966), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1967), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1968), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1969), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1970), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1971), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1972), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1973), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1974), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1975), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1976), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1977), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1978), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1979), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1980), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1981), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1982), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1983), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1984), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1985), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1986), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1987), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1988), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1989), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1990), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1991), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1992), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1993), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1994), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1995), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1996), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1997), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1998), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1999), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2000), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2001), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2002), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2003), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2004), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2005), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2006), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2007), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2008), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2009), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2010), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2011), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2012), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2013), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2014), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2015), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2016), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2017), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2018), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2019), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2020), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2021), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2022), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2023), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2024), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2025), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2026), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2027), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2028), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2029), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2030), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2031), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2032), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2033), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2034), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2035), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2036), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2037), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2038), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2039), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2040), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2041), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2042), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2043), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2044), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2045), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2046), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2047), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2048), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2049), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2050), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2051), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2052), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2053), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2054), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2055), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2056), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2057), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2058), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2059), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2060), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2061), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2062), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2063), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2064), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2065), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2066), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2067), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2068), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2069), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2070), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2071), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2072), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2073), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2074), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2075), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2076), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2077), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2078), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2079), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2080), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2081), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2082), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2083), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2084), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2085), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2086), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2087), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2088), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2089), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2090), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2091), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2092), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2093), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2094), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2095), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2096), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2097), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2098), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2099), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2100), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2101), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2102), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2103), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2104), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2105), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2106), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2107), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2108), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2109), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2110), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2111), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2112), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2113), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2114), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2115), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2116), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2117), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2118), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2119), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2120), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2121), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2122), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2123), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2124), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2125), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2126), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2127), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2128), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2129), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2130), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2131), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2132), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2133), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2134), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2135), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2136), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2137), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2138), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2139), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2140), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2141), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2142), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2143), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2144), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2145), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2146), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2147), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2148), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2149), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2150), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2151), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2152), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2153), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2154), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2155), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2156), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2157), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2166), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2167), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2168), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2169), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2170), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2171), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2172), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2173), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2174), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2175), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2176), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2177), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2178), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2179), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2180), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2181), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2182), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2183), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2184), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2185), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2186), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2187), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2188), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2189), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2190), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2191), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2192), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2193), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2194), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2195), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2196), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2197), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2198), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2199), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2200), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2201), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2202), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2203), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2204), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2205), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2206), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2207), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2208), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2209), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2210), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2211), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2212), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2213), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2214), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2215), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2216), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2217), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2218), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2219), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2220), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2221), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2222), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2223), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2224), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2225), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2226), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2227), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2228), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2229), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2230), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2231), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2232), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2233), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2234), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2235), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2236), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2237), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2238), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2239), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2240), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2241), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2242), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2243), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2244), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2245), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2246), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2247), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2248), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2249), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2250), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2251), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2252), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2253), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2254), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2255), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2256), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2257), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2258), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2259), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2260), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2261), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2262), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2263), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2264), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2265), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2266), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2267), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2268), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2269), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2270), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2271), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2272), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2273), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2274), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2275), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2276), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2277), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2278), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2279), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2280), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2281), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2282), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2283), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2284), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2285), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2286), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2287), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2288), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2289), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2290), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2291), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2292), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2293), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2294), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2295), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2296), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2297), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2298), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2299), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2300), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2301), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2302), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2303), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2304), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2305), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2306), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2307), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2308), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2309), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2310), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2311), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2312), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2313), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2314), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2315), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2316), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2317), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2318), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2319), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2320), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2321), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2322), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2323), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2324), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2325), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2326), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2327), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2328), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2329), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2330), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2331), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2332), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2333), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2334), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2335), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2336), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2337), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2338), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2339), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2340), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2341), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2342), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2343), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2344), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2345), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2346), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2347), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2348), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2349), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2350), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2351), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2352), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2353), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2354), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2355), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2356), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2357), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2358), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2359), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2360), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2361), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2362), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2363), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2364), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2365), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2366), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2367), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2368), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2369), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2370), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2371), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2372), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2373), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2374), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2375), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2376), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2377), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2378), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2379), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2380), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2381), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2382), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2383), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2384), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2385), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2386), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2387), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2388), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2389), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2390), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2391), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2392), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2393), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2394), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2395), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2396), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2397), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2398), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2399), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2400), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2401), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2402), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2403), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2404), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2405), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2406), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2407), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2408), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2409), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2410), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2411), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2412), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2413), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2414), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2415), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2416), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2417), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2418), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2419), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2420), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2421), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2422), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2423), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2424), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2425), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2426), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2427), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2428), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2429), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2430), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2431), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2432), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2433), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2434), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2435), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2436), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2437), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2438) );
  BUFX2 U2 ( .A(n24), .Y(n1) );
  INVX2 U3 ( .A(n6), .Y(n2) );
  INVX1 U4 ( .A(n6), .Y(n5) );
  INVX8 U5 ( .A(n97), .Y(n1366) );
  INVX8 U6 ( .A(n94), .Y(n1358) );
  AND2X2 U7 ( .A(\data_in<12> ), .B(n1227), .Y(n100) );
  AND2X2 U8 ( .A(\data_in<1> ), .B(n1227), .Y(n93) );
  AND2X2 U9 ( .A(\data_in<5> ), .B(n1351), .Y(n96) );
  INVX4 U10 ( .A(n73), .Y(n1353) );
  INVX1 U11 ( .A(write), .Y(n3) );
  INVX1 U12 ( .A(n3), .Y(n4) );
  INVX1 U13 ( .A(n1176), .Y(n1183) );
  INVX1 U14 ( .A(n1176), .Y(n1182) );
  INVX1 U15 ( .A(n1176), .Y(n1181) );
  INVX1 U16 ( .A(n1177), .Y(n1180) );
  INVX1 U17 ( .A(n1177), .Y(n1179) );
  INVX1 U18 ( .A(n1177), .Y(n1178) );
  INVX1 U19 ( .A(n1392), .Y(n1176) );
  INVX1 U20 ( .A(n1390), .Y(n1185) );
  INVX1 U21 ( .A(n1392), .Y(n1177) );
  INVX1 U22 ( .A(n1201), .Y(n1203) );
  INVX1 U23 ( .A(n1201), .Y(n1202) );
  INVX1 U24 ( .A(n1185), .Y(n1186) );
  INVX1 U25 ( .A(n1201), .Y(n1204) );
  INVX1 U26 ( .A(n1201), .Y(n1205) );
  INVX1 U27 ( .A(n1185), .Y(n1187) );
  INVX1 U28 ( .A(n1201), .Y(n1206) );
  INVX1 U29 ( .A(n1201), .Y(n1207) );
  INVX1 U30 ( .A(n1185), .Y(n1188) );
  INVX1 U31 ( .A(n1200), .Y(n1208) );
  INVX1 U32 ( .A(n1200), .Y(n1209) );
  INVX1 U33 ( .A(n1184), .Y(n1189) );
  INVX1 U34 ( .A(n1200), .Y(n1210) );
  INVX1 U35 ( .A(n1199), .Y(n1211) );
  INVX1 U36 ( .A(n1184), .Y(n1190) );
  INVX1 U37 ( .A(n1199), .Y(n1212) );
  INVX1 U38 ( .A(n1199), .Y(n1213) );
  INVX1 U39 ( .A(n1184), .Y(n1191) );
  INVX1 U40 ( .A(n1198), .Y(n1214) );
  INVX1 U41 ( .A(n1198), .Y(n1215) );
  INVX1 U42 ( .A(n1185), .Y(n1192) );
  INVX1 U43 ( .A(n1198), .Y(n1216) );
  INVX2 U44 ( .A(n1200), .Y(n1217) );
  INVX1 U45 ( .A(n1185), .Y(n1193) );
  INVX2 U46 ( .A(n1198), .Y(n1218) );
  INVX2 U47 ( .A(n1199), .Y(n1219) );
  INVX1 U48 ( .A(n1185), .Y(n1194) );
  INVX1 U49 ( .A(n1197), .Y(n1220) );
  INVX1 U50 ( .A(n1197), .Y(n1221) );
  INVX2 U51 ( .A(n1184), .Y(n1195) );
  INVX1 U52 ( .A(n1197), .Y(n1222) );
  INVX2 U53 ( .A(n1197), .Y(n1223) );
  INVX2 U54 ( .A(n1184), .Y(n1196) );
  INVX1 U55 ( .A(n645), .Y(N32) );
  INVX1 U56 ( .A(n646), .Y(N31) );
  INVX1 U57 ( .A(n647), .Y(N30) );
  INVX1 U58 ( .A(n648), .Y(N29) );
  INVX1 U59 ( .A(n649), .Y(N28) );
  INVX1 U60 ( .A(n650), .Y(N27) );
  INVX1 U61 ( .A(n1163), .Y(N26) );
  INVX1 U62 ( .A(n1164), .Y(N25) );
  INVX1 U63 ( .A(n1165), .Y(N24) );
  INVX1 U64 ( .A(n1166), .Y(N23) );
  INVX1 U65 ( .A(n1167), .Y(N22) );
  INVX1 U66 ( .A(n1168), .Y(N21) );
  INVX1 U67 ( .A(n1169), .Y(N20) );
  INVX1 U68 ( .A(n1170), .Y(N19) );
  INVX1 U69 ( .A(n1171), .Y(N18) );
  INVX1 U70 ( .A(n1172), .Y(N17) );
  BUFX2 U71 ( .A(n108), .Y(n1228) );
  BUFX2 U72 ( .A(n110), .Y(n1232) );
  BUFX2 U73 ( .A(n112), .Y(n1236) );
  BUFX2 U74 ( .A(n114), .Y(n1240) );
  BUFX2 U75 ( .A(n116), .Y(n1242) );
  BUFX2 U76 ( .A(n118), .Y(n1246) );
  BUFX2 U77 ( .A(n120), .Y(n1250) );
  BUFX2 U78 ( .A(n122), .Y(n1257) );
  BUFX2 U79 ( .A(n124), .Y(n1261) );
  BUFX2 U80 ( .A(n126), .Y(n1265) );
  BUFX2 U81 ( .A(n128), .Y(n1269) );
  BUFX2 U82 ( .A(n130), .Y(n1273) );
  BUFX2 U83 ( .A(n132), .Y(n1277) );
  BUFX2 U84 ( .A(n134), .Y(n1281) );
  BUFX2 U85 ( .A(n136), .Y(n1288) );
  BUFX2 U86 ( .A(n138), .Y(n1292) );
  BUFX2 U87 ( .A(n140), .Y(n1296) );
  BUFX2 U88 ( .A(n142), .Y(n1300) );
  BUFX2 U89 ( .A(n144), .Y(n1304) );
  BUFX2 U90 ( .A(n146), .Y(n1308) );
  BUFX2 U91 ( .A(n148), .Y(n1312) );
  BUFX2 U92 ( .A(n150), .Y(n1319) );
  BUFX2 U93 ( .A(n152), .Y(n1323) );
  BUFX2 U94 ( .A(n154), .Y(n1327) );
  BUFX2 U95 ( .A(n156), .Y(n1331) );
  BUFX2 U96 ( .A(n158), .Y(n1335) );
  BUFX2 U97 ( .A(n160), .Y(n1339) );
  BUFX2 U98 ( .A(n162), .Y(n1343) );
  INVX1 U99 ( .A(n1395), .Y(n1175) );
  INVX1 U100 ( .A(n1395), .Y(n1174) );
  INVX1 U101 ( .A(n1397), .Y(n1396) );
  INVX1 U102 ( .A(N14), .Y(n1397) );
  INVX1 U103 ( .A(N10), .Y(n1201) );
  INVX1 U104 ( .A(n1388), .Y(n1198) );
  INVX1 U105 ( .A(n1388), .Y(n1199) );
  INVX1 U106 ( .A(n1388), .Y(n1200) );
  INVX1 U107 ( .A(n1397), .Y(n1173) );
  INVX1 U108 ( .A(n1388), .Y(n1197) );
  INVX1 U109 ( .A(n1395), .Y(n1394) );
  INVX1 U110 ( .A(N13), .Y(n1395) );
  INVX1 U111 ( .A(n1390), .Y(n1184) );
  BUFX2 U112 ( .A(n108), .Y(n1229) );
  BUFX2 U113 ( .A(n110), .Y(n1233) );
  BUFX2 U114 ( .A(n112), .Y(n1237) );
  BUFX2 U115 ( .A(n120), .Y(n1251) );
  INVX1 U116 ( .A(rst), .Y(n1387) );
  INVX1 U117 ( .A(n105), .Y(n1316) );
  INVX1 U118 ( .A(n106), .Y(n1347) );
  BUFX2 U119 ( .A(n126), .Y(n1266) );
  BUFX2 U120 ( .A(n128), .Y(n1270) );
  BUFX2 U121 ( .A(n130), .Y(n1274) );
  BUFX2 U122 ( .A(n132), .Y(n1278) );
  BUFX2 U123 ( .A(n134), .Y(n1282) );
  BUFX2 U124 ( .A(n140), .Y(n1297) );
  BUFX2 U125 ( .A(n144), .Y(n1305) );
  BUFX2 U126 ( .A(n146), .Y(n1309) );
  BUFX2 U127 ( .A(n148), .Y(n1313) );
  BUFX2 U128 ( .A(n154), .Y(n1328) );
  BUFX2 U129 ( .A(n158), .Y(n1336) );
  BUFX2 U130 ( .A(n160), .Y(n1340) );
  BUFX2 U131 ( .A(n162), .Y(n1344) );
  BUFX2 U132 ( .A(n116), .Y(n1243) );
  BUFX2 U133 ( .A(n118), .Y(n1247) );
  BUFX2 U134 ( .A(n122), .Y(n1258) );
  BUFX2 U135 ( .A(n124), .Y(n1262) );
  BUFX2 U136 ( .A(n136), .Y(n1289) );
  BUFX2 U137 ( .A(n138), .Y(n1293) );
  BUFX2 U138 ( .A(n142), .Y(n1301) );
  BUFX2 U139 ( .A(n150), .Y(n1320) );
  BUFX2 U140 ( .A(n152), .Y(n1324) );
  BUFX2 U141 ( .A(n156), .Y(n1332) );
  BUFX2 U142 ( .A(n114), .Y(n1241) );
  INVX1 U143 ( .A(n103), .Y(n1254) );
  INVX1 U144 ( .A(n104), .Y(n1285) );
  INVX2 U145 ( .A(n6), .Y(n7) );
  OR2X2 U146 ( .A(write), .B(rst), .Y(n6) );
  AND2X2 U147 ( .A(\data_in<0> ), .B(n1351), .Y(n8) );
  AND2X2 U148 ( .A(n1350), .B(n107), .Y(n9) );
  INVX1 U149 ( .A(n9), .Y(n10) );
  AND2X2 U150 ( .A(\data_in<8> ), .B(n1227), .Y(n11) );
  AND2X2 U151 ( .A(\data_in<10> ), .B(n1227), .Y(n12) );
  AND2X2 U152 ( .A(n1350), .B(n109), .Y(n13) );
  INVX1 U153 ( .A(n13), .Y(n14) );
  AND2X2 U154 ( .A(n1350), .B(n111), .Y(n15) );
  INVX1 U155 ( .A(n15), .Y(n16) );
  AND2X2 U156 ( .A(n1350), .B(n115), .Y(n17) );
  INVX1 U157 ( .A(n17), .Y(n18) );
  AND2X2 U158 ( .A(n1350), .B(n117), .Y(n19) );
  INVX1 U159 ( .A(n19), .Y(n20) );
  AND2X2 U160 ( .A(n1350), .B(n119), .Y(n21) );
  INVX1 U161 ( .A(n21), .Y(n22) );
  AND2X2 U162 ( .A(n1350), .B(n103), .Y(n23) );
  INVX1 U163 ( .A(n23), .Y(n24) );
  AND2X2 U164 ( .A(n1350), .B(n121), .Y(n25) );
  INVX1 U165 ( .A(n25), .Y(n26) );
  AND2X2 U166 ( .A(n1350), .B(n123), .Y(n27) );
  INVX1 U167 ( .A(n27), .Y(n28) );
  AND2X2 U168 ( .A(n1350), .B(n125), .Y(n29) );
  INVX1 U169 ( .A(n29), .Y(n30) );
  AND2X2 U170 ( .A(n1350), .B(n127), .Y(n31) );
  INVX1 U171 ( .A(n31), .Y(n32) );
  AND2X2 U172 ( .A(n1352), .B(n129), .Y(n33) );
  INVX1 U173 ( .A(n33), .Y(n34) );
  AND2X2 U174 ( .A(n1352), .B(n131), .Y(n35) );
  INVX1 U175 ( .A(n35), .Y(n36) );
  AND2X2 U176 ( .A(n1352), .B(n133), .Y(n37) );
  INVX1 U177 ( .A(n37), .Y(n38) );
  AND2X2 U178 ( .A(n1352), .B(n104), .Y(n39) );
  INVX1 U179 ( .A(n39), .Y(n40) );
  AND2X2 U180 ( .A(n1352), .B(n135), .Y(n41) );
  INVX1 U181 ( .A(n41), .Y(n42) );
  AND2X2 U182 ( .A(n1352), .B(n137), .Y(n43) );
  INVX1 U183 ( .A(n43), .Y(n44) );
  AND2X2 U184 ( .A(n1352), .B(n139), .Y(n45) );
  INVX1 U185 ( .A(n45), .Y(n46) );
  AND2X2 U186 ( .A(n1352), .B(n141), .Y(n47) );
  INVX1 U187 ( .A(n47), .Y(n48) );
  AND2X2 U188 ( .A(n1352), .B(n143), .Y(n49) );
  INVX1 U189 ( .A(n49), .Y(n50) );
  AND2X2 U190 ( .A(n1352), .B(n145), .Y(n51) );
  INVX1 U191 ( .A(n51), .Y(n52) );
  AND2X2 U192 ( .A(n1352), .B(n147), .Y(n53) );
  INVX1 U193 ( .A(n53), .Y(n54) );
  AND2X2 U194 ( .A(n1352), .B(n105), .Y(n55) );
  INVX1 U195 ( .A(n55), .Y(n56) );
  AND2X2 U196 ( .A(n1352), .B(n149), .Y(n57) );
  INVX1 U197 ( .A(n57), .Y(n58) );
  AND2X2 U198 ( .A(n1352), .B(n151), .Y(n59) );
  INVX1 U199 ( .A(n59), .Y(n60) );
  AND2X2 U200 ( .A(n1352), .B(n153), .Y(n61) );
  INVX1 U201 ( .A(n61), .Y(n62) );
  AND2X2 U202 ( .A(n1352), .B(n155), .Y(n63) );
  INVX1 U203 ( .A(n63), .Y(n64) );
  AND2X2 U204 ( .A(n1352), .B(n157), .Y(n65) );
  INVX1 U205 ( .A(n65), .Y(n66) );
  AND2X2 U206 ( .A(n1352), .B(n159), .Y(n67) );
  INVX1 U207 ( .A(n67), .Y(n68) );
  AND2X2 U208 ( .A(n1352), .B(n161), .Y(n69) );
  INVX1 U209 ( .A(n69), .Y(n70) );
  AND2X2 U210 ( .A(n1352), .B(n106), .Y(n71) );
  INVX1 U211 ( .A(n71), .Y(n72) );
  BUFX2 U212 ( .A(n34), .Y(n1275) );
  BUFX2 U213 ( .A(n38), .Y(n1283) );
  BUFX2 U214 ( .A(n40), .Y(n1286) );
  BUFX2 U215 ( .A(n40), .Y(n1287) );
  BUFX2 U216 ( .A(n44), .Y(n1294) );
  BUFX2 U217 ( .A(n48), .Y(n1302) );
  BUFX2 U218 ( .A(n52), .Y(n1310) );
  BUFX2 U219 ( .A(n56), .Y(n1317) );
  BUFX2 U220 ( .A(n56), .Y(n1318) );
  BUFX2 U221 ( .A(n58), .Y(n1321) );
  BUFX2 U222 ( .A(n58), .Y(n1322) );
  BUFX2 U223 ( .A(n60), .Y(n1325) );
  BUFX2 U224 ( .A(n60), .Y(n1326) );
  BUFX2 U225 ( .A(n62), .Y(n1329) );
  BUFX2 U226 ( .A(n62), .Y(n1330) );
  BUFX2 U227 ( .A(n64), .Y(n1333) );
  BUFX2 U228 ( .A(n64), .Y(n1334) );
  BUFX2 U229 ( .A(n66), .Y(n1337) );
  BUFX2 U230 ( .A(n66), .Y(n1338) );
  BUFX2 U231 ( .A(n68), .Y(n1341) );
  BUFX2 U232 ( .A(n68), .Y(n1342) );
  BUFX2 U233 ( .A(n70), .Y(n1345) );
  BUFX2 U234 ( .A(n70), .Y(n1346) );
  BUFX2 U235 ( .A(n72), .Y(n1348) );
  BUFX2 U236 ( .A(n72), .Y(n1349) );
  AND2X2 U237 ( .A(n4), .B(n1387), .Y(n73) );
  INVX1 U238 ( .A(n1393), .Y(n1392) );
  INVX1 U239 ( .A(n1389), .Y(n1388) );
  INVX1 U240 ( .A(N12), .Y(n1393) );
  AND2X1 U241 ( .A(n1392), .B(n1390), .Y(n74) );
  INVX1 U242 ( .A(n1391), .Y(n1390) );
  AND2X1 U243 ( .A(n2438), .B(n1396), .Y(n75) );
  AND2X2 U244 ( .A(\data_in<4> ), .B(n1351), .Y(n76) );
  INVX1 U245 ( .A(n76), .Y(n77) );
  AND2X2 U246 ( .A(\data_in<9> ), .B(n1351), .Y(n78) );
  INVX1 U247 ( .A(n78), .Y(n79) );
  AND2X2 U248 ( .A(\data_in<15> ), .B(n1351), .Y(n80) );
  INVX1 U249 ( .A(n80), .Y(n81) );
  INVX1 U250 ( .A(n1353), .Y(n1351) );
  INVX2 U251 ( .A(n163), .Y(n1463) );
  BUFX2 U252 ( .A(n1430), .Y(n82) );
  INVX1 U253 ( .A(n82), .Y(n1823) );
  BUFX2 U254 ( .A(n1447), .Y(n83) );
  INVX1 U255 ( .A(n83), .Y(n1840) );
  BUFX2 U256 ( .A(n1465), .Y(n84) );
  INVX1 U257 ( .A(n84), .Y(n1857) );
  BUFX2 U258 ( .A(n1482), .Y(n85) );
  INVX1 U259 ( .A(n85), .Y(n1874) );
  BUFX2 U260 ( .A(n1499), .Y(n86) );
  INVX1 U261 ( .A(n86), .Y(n1891) );
  BUFX2 U262 ( .A(n1660), .Y(n87) );
  INVX1 U263 ( .A(n87), .Y(n1773) );
  BUFX2 U264 ( .A(n1790), .Y(n88) );
  INVX1 U265 ( .A(n88), .Y(n1908) );
  AND2X1 U266 ( .A(n1388), .B(n74), .Y(n89) );
  AND2X1 U267 ( .A(n1394), .B(n75), .Y(n90) );
  AND2X1 U268 ( .A(n1389), .B(n74), .Y(n91) );
  AND2X1 U269 ( .A(n1395), .B(n75), .Y(n92) );
  AND2X2 U270 ( .A(\data_in<2> ), .B(n1352), .Y(n94) );
  AND2X2 U271 ( .A(\data_in<3> ), .B(n1352), .Y(n95) );
  AND2X2 U272 ( .A(\data_in<6> ), .B(n1352), .Y(n97) );
  AND2X2 U273 ( .A(\data_in<7> ), .B(n1227), .Y(n98) );
  AND2X2 U274 ( .A(\data_in<11> ), .B(n1351), .Y(n99) );
  AND2X2 U275 ( .A(\data_in<13> ), .B(n1351), .Y(n101) );
  AND2X2 U276 ( .A(\data_in<14> ), .B(n1227), .Y(n102) );
  AND2X1 U277 ( .A(n90), .B(n1909), .Y(n103) );
  AND2X1 U278 ( .A(n1909), .B(n92), .Y(n104) );
  AND2X1 U279 ( .A(n1909), .B(n1773), .Y(n105) );
  AND2X1 U280 ( .A(n1909), .B(n1908), .Y(n106) );
  AND2X1 U281 ( .A(n89), .B(n90), .Y(n107) );
  INVX1 U282 ( .A(n107), .Y(n108) );
  AND2X1 U283 ( .A(n90), .B(n91), .Y(n109) );
  INVX1 U284 ( .A(n109), .Y(n110) );
  AND2X1 U285 ( .A(n90), .B(n1823), .Y(n111) );
  INVX1 U286 ( .A(n111), .Y(n112) );
  AND2X1 U287 ( .A(n90), .B(n1840), .Y(n113) );
  INVX1 U288 ( .A(n113), .Y(n114) );
  AND2X1 U289 ( .A(n90), .B(n1857), .Y(n115) );
  INVX1 U290 ( .A(n115), .Y(n116) );
  AND2X1 U291 ( .A(n90), .B(n1874), .Y(n117) );
  INVX1 U292 ( .A(n117), .Y(n118) );
  AND2X1 U293 ( .A(n90), .B(n1891), .Y(n119) );
  INVX1 U294 ( .A(n119), .Y(n120) );
  AND2X1 U295 ( .A(n89), .B(n92), .Y(n121) );
  INVX1 U296 ( .A(n121), .Y(n122) );
  AND2X1 U297 ( .A(n91), .B(n92), .Y(n123) );
  INVX1 U298 ( .A(n123), .Y(n124) );
  AND2X1 U299 ( .A(n1823), .B(n92), .Y(n125) );
  INVX1 U300 ( .A(n125), .Y(n126) );
  AND2X1 U301 ( .A(n1840), .B(n92), .Y(n127) );
  INVX1 U302 ( .A(n127), .Y(n128) );
  AND2X1 U303 ( .A(n1857), .B(n92), .Y(n129) );
  INVX1 U304 ( .A(n129), .Y(n130) );
  AND2X1 U305 ( .A(n1874), .B(n92), .Y(n131) );
  INVX1 U306 ( .A(n131), .Y(n132) );
  AND2X1 U307 ( .A(n1891), .B(n92), .Y(n133) );
  INVX1 U308 ( .A(n133), .Y(n134) );
  AND2X1 U309 ( .A(n89), .B(n1773), .Y(n135) );
  INVX1 U310 ( .A(n135), .Y(n136) );
  AND2X1 U311 ( .A(n91), .B(n1773), .Y(n137) );
  INVX1 U312 ( .A(n137), .Y(n138) );
  AND2X1 U313 ( .A(n1823), .B(n1773), .Y(n139) );
  INVX1 U314 ( .A(n139), .Y(n140) );
  AND2X1 U315 ( .A(n1840), .B(n1773), .Y(n141) );
  INVX1 U316 ( .A(n141), .Y(n142) );
  AND2X1 U317 ( .A(n1857), .B(n1773), .Y(n143) );
  INVX1 U318 ( .A(n143), .Y(n144) );
  AND2X1 U319 ( .A(n1874), .B(n1773), .Y(n145) );
  INVX1 U320 ( .A(n145), .Y(n146) );
  AND2X1 U321 ( .A(n1891), .B(n1773), .Y(n147) );
  INVX1 U322 ( .A(n147), .Y(n148) );
  AND2X1 U323 ( .A(n89), .B(n1908), .Y(n149) );
  INVX1 U324 ( .A(n149), .Y(n150) );
  AND2X1 U325 ( .A(n91), .B(n1908), .Y(n151) );
  INVX1 U326 ( .A(n151), .Y(n152) );
  AND2X1 U327 ( .A(n1823), .B(n1908), .Y(n153) );
  INVX1 U328 ( .A(n153), .Y(n154) );
  AND2X1 U329 ( .A(n1840), .B(n1908), .Y(n155) );
  INVX1 U330 ( .A(n155), .Y(n156) );
  AND2X1 U331 ( .A(n1857), .B(n1908), .Y(n157) );
  INVX1 U332 ( .A(n157), .Y(n158) );
  AND2X1 U333 ( .A(n1874), .B(n1908), .Y(n159) );
  INVX1 U334 ( .A(n159), .Y(n160) );
  AND2X1 U335 ( .A(n1891), .B(n1908), .Y(n161) );
  INVX1 U336 ( .A(n161), .Y(n162) );
  BUFX2 U337 ( .A(n32), .Y(n1271) );
  BUFX2 U338 ( .A(n28), .Y(n1263) );
  BUFX2 U339 ( .A(n22), .Y(n1252) );
  BUFX2 U340 ( .A(n18), .Y(n1244) );
  AND2X2 U341 ( .A(n1350), .B(n113), .Y(n163) );
  BUFX2 U342 ( .A(n10), .Y(n1231) );
  BUFX2 U343 ( .A(n24), .Y(n1256) );
  BUFX2 U344 ( .A(n24), .Y(n1255) );
  BUFX2 U345 ( .A(n32), .Y(n1272) );
  BUFX2 U346 ( .A(n30), .Y(n1267) );
  BUFX2 U347 ( .A(n30), .Y(n1268) );
  BUFX2 U348 ( .A(n28), .Y(n1264) );
  BUFX2 U349 ( .A(n26), .Y(n1259) );
  BUFX2 U350 ( .A(n26), .Y(n1260) );
  BUFX2 U351 ( .A(n22), .Y(n1253) );
  BUFX2 U352 ( .A(n20), .Y(n1248) );
  BUFX2 U353 ( .A(n20), .Y(n1249) );
  BUFX2 U354 ( .A(n18), .Y(n1245) );
  BUFX2 U355 ( .A(n16), .Y(n1238) );
  BUFX2 U356 ( .A(n16), .Y(n1239) );
  BUFX2 U357 ( .A(n14), .Y(n1234) );
  BUFX2 U358 ( .A(n14), .Y(n1235) );
  BUFX2 U359 ( .A(n10), .Y(n1230) );
  INVX4 U360 ( .A(n1353), .Y(n1350) );
  INVX1 U361 ( .A(N11), .Y(n1391) );
  MUX2X1 U362 ( .B(n165), .A(n166), .S(n1186), .Y(n164) );
  MUX2X1 U363 ( .B(n168), .A(n169), .S(n1186), .Y(n167) );
  MUX2X1 U364 ( .B(n171), .A(n172), .S(n1186), .Y(n170) );
  MUX2X1 U365 ( .B(n174), .A(n175), .S(n1186), .Y(n173) );
  MUX2X1 U366 ( .B(n177), .A(n178), .S(n1175), .Y(n176) );
  MUX2X1 U367 ( .B(n180), .A(n181), .S(n1186), .Y(n179) );
  MUX2X1 U368 ( .B(n183), .A(n184), .S(n1186), .Y(n182) );
  MUX2X1 U369 ( .B(n186), .A(n187), .S(n1186), .Y(n185) );
  MUX2X1 U370 ( .B(n189), .A(n190), .S(n1186), .Y(n188) );
  MUX2X1 U371 ( .B(n192), .A(n193), .S(n1175), .Y(n191) );
  MUX2X1 U372 ( .B(n195), .A(n196), .S(n1187), .Y(n194) );
  MUX2X1 U373 ( .B(n198), .A(n199), .S(n1187), .Y(n197) );
  MUX2X1 U374 ( .B(n201), .A(n202), .S(n1187), .Y(n200) );
  MUX2X1 U375 ( .B(n204), .A(n205), .S(n1187), .Y(n203) );
  MUX2X1 U376 ( .B(n207), .A(n208), .S(n1175), .Y(n206) );
  MUX2X1 U377 ( .B(n210), .A(n211), .S(n1187), .Y(n209) );
  MUX2X1 U378 ( .B(n213), .A(n215), .S(n1187), .Y(n212) );
  MUX2X1 U379 ( .B(n217), .A(n218), .S(n1187), .Y(n216) );
  MUX2X1 U380 ( .B(n220), .A(n221), .S(n1187), .Y(n219) );
  MUX2X1 U381 ( .B(n223), .A(n224), .S(n1175), .Y(n222) );
  MUX2X1 U382 ( .B(n226), .A(n227), .S(n1187), .Y(n225) );
  MUX2X1 U383 ( .B(n229), .A(n230), .S(n1187), .Y(n228) );
  MUX2X1 U384 ( .B(n232), .A(n233), .S(n1187), .Y(n231) );
  MUX2X1 U385 ( .B(n235), .A(n236), .S(n1187), .Y(n234) );
  MUX2X1 U386 ( .B(n238), .A(n239), .S(n1175), .Y(n237) );
  MUX2X1 U387 ( .B(n241), .A(n242), .S(n1188), .Y(n240) );
  MUX2X1 U388 ( .B(n244), .A(n245), .S(n1188), .Y(n243) );
  MUX2X1 U389 ( .B(n247), .A(n248), .S(n1188), .Y(n246) );
  MUX2X1 U390 ( .B(n250), .A(n251), .S(n1188), .Y(n249) );
  MUX2X1 U391 ( .B(n253), .A(n254), .S(n1175), .Y(n252) );
  MUX2X1 U392 ( .B(n256), .A(n257), .S(n1188), .Y(n255) );
  MUX2X1 U393 ( .B(n259), .A(n260), .S(n1188), .Y(n258) );
  MUX2X1 U394 ( .B(n262), .A(n263), .S(n1188), .Y(n261) );
  MUX2X1 U395 ( .B(n265), .A(n266), .S(n1188), .Y(n264) );
  MUX2X1 U396 ( .B(n268), .A(n269), .S(n1175), .Y(n267) );
  MUX2X1 U397 ( .B(n271), .A(n272), .S(n1188), .Y(n270) );
  MUX2X1 U398 ( .B(n274), .A(n275), .S(n1188), .Y(n273) );
  MUX2X1 U399 ( .B(n277), .A(n278), .S(n1188), .Y(n276) );
  MUX2X1 U400 ( .B(n280), .A(n281), .S(n1188), .Y(n279) );
  MUX2X1 U401 ( .B(n283), .A(n284), .S(n1175), .Y(n282) );
  MUX2X1 U402 ( .B(n286), .A(n287), .S(n1189), .Y(n285) );
  MUX2X1 U403 ( .B(n289), .A(n290), .S(n1189), .Y(n288) );
  MUX2X1 U404 ( .B(n292), .A(n293), .S(n1189), .Y(n291) );
  MUX2X1 U405 ( .B(n295), .A(n296), .S(n1189), .Y(n294) );
  MUX2X1 U406 ( .B(n298), .A(n299), .S(n1175), .Y(n297) );
  MUX2X1 U407 ( .B(n301), .A(n302), .S(n1189), .Y(n300) );
  MUX2X1 U408 ( .B(n304), .A(n305), .S(n1189), .Y(n303) );
  MUX2X1 U409 ( .B(n307), .A(n308), .S(n1189), .Y(n306) );
  MUX2X1 U410 ( .B(n310), .A(n311), .S(n1189), .Y(n309) );
  MUX2X1 U411 ( .B(n313), .A(n314), .S(n1175), .Y(n312) );
  MUX2X1 U412 ( .B(n316), .A(n317), .S(n1189), .Y(n315) );
  MUX2X1 U413 ( .B(n319), .A(n320), .S(n1189), .Y(n318) );
  MUX2X1 U414 ( .B(n322), .A(n323), .S(n1189), .Y(n321) );
  MUX2X1 U415 ( .B(n325), .A(n326), .S(n1189), .Y(n324) );
  MUX2X1 U416 ( .B(n328), .A(n329), .S(n1175), .Y(n327) );
  MUX2X1 U417 ( .B(n331), .A(n332), .S(n1190), .Y(n330) );
  MUX2X1 U418 ( .B(n334), .A(n335), .S(n1190), .Y(n333) );
  MUX2X1 U419 ( .B(n337), .A(n338), .S(n1190), .Y(n336) );
  MUX2X1 U420 ( .B(n340), .A(n341), .S(n1190), .Y(n339) );
  MUX2X1 U421 ( .B(n343), .A(n344), .S(n1175), .Y(n342) );
  MUX2X1 U422 ( .B(n346), .A(n347), .S(n1190), .Y(n345) );
  MUX2X1 U423 ( .B(n349), .A(n350), .S(n1190), .Y(n348) );
  MUX2X1 U424 ( .B(n352), .A(n353), .S(n1190), .Y(n351) );
  MUX2X1 U425 ( .B(n355), .A(n356), .S(n1190), .Y(n354) );
  MUX2X1 U426 ( .B(n358), .A(n359), .S(n1174), .Y(n357) );
  MUX2X1 U427 ( .B(n361), .A(n362), .S(n1190), .Y(n360) );
  MUX2X1 U428 ( .B(n364), .A(n365), .S(n1190), .Y(n363) );
  MUX2X1 U429 ( .B(n367), .A(n368), .S(n1190), .Y(n366) );
  MUX2X1 U430 ( .B(n370), .A(n371), .S(n1190), .Y(n369) );
  MUX2X1 U431 ( .B(n373), .A(n374), .S(n1174), .Y(n372) );
  MUX2X1 U432 ( .B(n376), .A(n377), .S(n1191), .Y(n375) );
  MUX2X1 U433 ( .B(n379), .A(n380), .S(n1191), .Y(n378) );
  MUX2X1 U434 ( .B(n382), .A(n383), .S(n1191), .Y(n381) );
  MUX2X1 U435 ( .B(n385), .A(n386), .S(n1191), .Y(n384) );
  MUX2X1 U436 ( .B(n388), .A(n389), .S(n1174), .Y(n387) );
  MUX2X1 U437 ( .B(n391), .A(n392), .S(n1191), .Y(n390) );
  MUX2X1 U438 ( .B(n394), .A(n395), .S(n1191), .Y(n393) );
  MUX2X1 U439 ( .B(n397), .A(n398), .S(n1191), .Y(n396) );
  MUX2X1 U440 ( .B(n400), .A(n401), .S(n1191), .Y(n399) );
  MUX2X1 U441 ( .B(n403), .A(n404), .S(n1174), .Y(n402) );
  MUX2X1 U442 ( .B(n406), .A(n407), .S(n1191), .Y(n405) );
  MUX2X1 U443 ( .B(n409), .A(n410), .S(n1191), .Y(n408) );
  MUX2X1 U444 ( .B(n412), .A(n413), .S(n1191), .Y(n411) );
  MUX2X1 U445 ( .B(n415), .A(n416), .S(n1191), .Y(n414) );
  MUX2X1 U446 ( .B(n418), .A(n419), .S(n1174), .Y(n417) );
  MUX2X1 U447 ( .B(n421), .A(n422), .S(n1192), .Y(n420) );
  MUX2X1 U448 ( .B(n424), .A(n425), .S(n1192), .Y(n423) );
  MUX2X1 U449 ( .B(n427), .A(n428), .S(n1192), .Y(n426) );
  MUX2X1 U450 ( .B(n430), .A(n431), .S(n1192), .Y(n429) );
  MUX2X1 U451 ( .B(n433), .A(n434), .S(n1174), .Y(n432) );
  MUX2X1 U452 ( .B(n436), .A(n437), .S(n1192), .Y(n435) );
  MUX2X1 U453 ( .B(n439), .A(n440), .S(n1192), .Y(n438) );
  MUX2X1 U454 ( .B(n442), .A(n443), .S(n1192), .Y(n441) );
  MUX2X1 U455 ( .B(n445), .A(n446), .S(n1192), .Y(n444) );
  MUX2X1 U456 ( .B(n448), .A(n449), .S(n1174), .Y(n447) );
  MUX2X1 U457 ( .B(n451), .A(n452), .S(n1192), .Y(n450) );
  MUX2X1 U458 ( .B(n454), .A(n455), .S(n1192), .Y(n453) );
  MUX2X1 U459 ( .B(n457), .A(n458), .S(n1192), .Y(n456) );
  MUX2X1 U460 ( .B(n460), .A(n461), .S(n1192), .Y(n459) );
  MUX2X1 U461 ( .B(n463), .A(n464), .S(n1174), .Y(n462) );
  MUX2X1 U462 ( .B(n466), .A(n467), .S(n1193), .Y(n465) );
  MUX2X1 U463 ( .B(n469), .A(n470), .S(n1193), .Y(n468) );
  MUX2X1 U464 ( .B(n472), .A(n473), .S(n1193), .Y(n471) );
  MUX2X1 U465 ( .B(n475), .A(n476), .S(n1193), .Y(n474) );
  MUX2X1 U466 ( .B(n478), .A(n479), .S(n1174), .Y(n477) );
  MUX2X1 U467 ( .B(n481), .A(n482), .S(n1193), .Y(n480) );
  MUX2X1 U468 ( .B(n484), .A(n485), .S(n1193), .Y(n483) );
  MUX2X1 U469 ( .B(n487), .A(n488), .S(n1193), .Y(n486) );
  MUX2X1 U470 ( .B(n490), .A(n491), .S(n1193), .Y(n489) );
  MUX2X1 U471 ( .B(n493), .A(n494), .S(n1174), .Y(n492) );
  MUX2X1 U472 ( .B(n496), .A(n497), .S(n1193), .Y(n495) );
  MUX2X1 U473 ( .B(n499), .A(n500), .S(n1193), .Y(n498) );
  MUX2X1 U474 ( .B(n502), .A(n503), .S(n1193), .Y(n501) );
  MUX2X1 U475 ( .B(n505), .A(n506), .S(n1193), .Y(n504) );
  MUX2X1 U476 ( .B(n508), .A(n509), .S(n1174), .Y(n507) );
  MUX2X1 U477 ( .B(n511), .A(n512), .S(n1194), .Y(n510) );
  MUX2X1 U478 ( .B(n514), .A(n515), .S(n1194), .Y(n513) );
  MUX2X1 U479 ( .B(n517), .A(n518), .S(n1194), .Y(n516) );
  MUX2X1 U480 ( .B(n520), .A(n521), .S(n1194), .Y(n519) );
  MUX2X1 U481 ( .B(n523), .A(n524), .S(n1174), .Y(n522) );
  MUX2X1 U482 ( .B(n526), .A(n527), .S(n1194), .Y(n525) );
  MUX2X1 U483 ( .B(n529), .A(n530), .S(n1194), .Y(n528) );
  MUX2X1 U484 ( .B(n532), .A(n533), .S(n1194), .Y(n531) );
  MUX2X1 U485 ( .B(n535), .A(n536), .S(n1194), .Y(n534) );
  MUX2X1 U486 ( .B(n538), .A(n539), .S(n1174), .Y(n537) );
  MUX2X1 U487 ( .B(n541), .A(n542), .S(n1194), .Y(n540) );
  MUX2X1 U488 ( .B(n544), .A(n545), .S(n1194), .Y(n543) );
  MUX2X1 U489 ( .B(n547), .A(n548), .S(n1194), .Y(n546) );
  MUX2X1 U490 ( .B(n550), .A(n551), .S(n1194), .Y(n549) );
  MUX2X1 U491 ( .B(n553), .A(n554), .S(n1174), .Y(n552) );
  MUX2X1 U492 ( .B(n556), .A(n557), .S(n1195), .Y(n555) );
  MUX2X1 U493 ( .B(n559), .A(n560), .S(n1195), .Y(n558) );
  MUX2X1 U494 ( .B(n562), .A(n563), .S(n1195), .Y(n561) );
  MUX2X1 U495 ( .B(n565), .A(n566), .S(n1195), .Y(n564) );
  MUX2X1 U496 ( .B(n568), .A(n569), .S(n1175), .Y(n567) );
  MUX2X1 U497 ( .B(n571), .A(n572), .S(n1195), .Y(n570) );
  MUX2X1 U498 ( .B(n574), .A(n575), .S(n1195), .Y(n573) );
  MUX2X1 U499 ( .B(n577), .A(n578), .S(n1195), .Y(n576) );
  MUX2X1 U500 ( .B(n580), .A(n581), .S(n1195), .Y(n579) );
  MUX2X1 U501 ( .B(n583), .A(n584), .S(n1175), .Y(n582) );
  MUX2X1 U502 ( .B(n586), .A(n587), .S(n1195), .Y(n585) );
  MUX2X1 U503 ( .B(n589), .A(n590), .S(n1195), .Y(n588) );
  MUX2X1 U504 ( .B(n592), .A(n593), .S(n1195), .Y(n591) );
  MUX2X1 U505 ( .B(n595), .A(n596), .S(n1195), .Y(n594) );
  MUX2X1 U506 ( .B(n598), .A(n599), .S(n1174), .Y(n597) );
  MUX2X1 U507 ( .B(n601), .A(n602), .S(n1196), .Y(n600) );
  MUX2X1 U508 ( .B(n604), .A(n605), .S(n1196), .Y(n603) );
  MUX2X1 U509 ( .B(n607), .A(n608), .S(n1196), .Y(n606) );
  MUX2X1 U510 ( .B(n610), .A(n611), .S(n1196), .Y(n609) );
  MUX2X1 U511 ( .B(n613), .A(n614), .S(n1174), .Y(n612) );
  MUX2X1 U512 ( .B(n616), .A(n617), .S(n1196), .Y(n615) );
  MUX2X1 U513 ( .B(n619), .A(n620), .S(n1196), .Y(n618) );
  MUX2X1 U514 ( .B(n622), .A(n623), .S(n1196), .Y(n621) );
  MUX2X1 U515 ( .B(n625), .A(n626), .S(n1196), .Y(n624) );
  MUX2X1 U516 ( .B(n628), .A(n629), .S(n1175), .Y(n627) );
  MUX2X1 U517 ( .B(n631), .A(n632), .S(n1196), .Y(n630) );
  MUX2X1 U518 ( .B(n634), .A(n635), .S(n1196), .Y(n633) );
  MUX2X1 U519 ( .B(n637), .A(n638), .S(n1196), .Y(n636) );
  MUX2X1 U520 ( .B(n640), .A(n641), .S(n1196), .Y(n639) );
  MUX2X1 U521 ( .B(n643), .A(n644), .S(n1175), .Y(n642) );
  MUX2X1 U522 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1202), .Y(n166) );
  MUX2X1 U523 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1202), .Y(n165) );
  MUX2X1 U524 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1202), .Y(n169) );
  MUX2X1 U525 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1202), .Y(n168) );
  MUX2X1 U526 ( .B(n167), .A(n164), .S(n1183), .Y(n178) );
  MUX2X1 U527 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1203), .Y(n172) );
  MUX2X1 U528 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1203), .Y(n171) );
  MUX2X1 U529 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1203), .Y(n175) );
  MUX2X1 U530 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1203), .Y(n174) );
  MUX2X1 U531 ( .B(n173), .A(n170), .S(n1183), .Y(n177) );
  MUX2X1 U532 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1203), .Y(n181) );
  MUX2X1 U533 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1203), .Y(n180) );
  MUX2X1 U534 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1203), .Y(n184) );
  MUX2X1 U535 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1203), .Y(n183) );
  MUX2X1 U536 ( .B(n182), .A(n179), .S(n1183), .Y(n193) );
  MUX2X1 U537 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1203), .Y(n187) );
  MUX2X1 U538 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1203), .Y(n186) );
  MUX2X1 U539 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1203), .Y(n190) );
  MUX2X1 U540 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1203), .Y(n189) );
  MUX2X1 U541 ( .B(n188), .A(n185), .S(n1183), .Y(n192) );
  MUX2X1 U542 ( .B(n191), .A(n176), .S(n1173), .Y(n645) );
  MUX2X1 U543 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1204), .Y(n196) );
  MUX2X1 U544 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1204), .Y(n195) );
  MUX2X1 U545 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1204), .Y(n199) );
  MUX2X1 U546 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1204), .Y(n198) );
  MUX2X1 U547 ( .B(n197), .A(n194), .S(n1183), .Y(n208) );
  MUX2X1 U548 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1204), .Y(n202) );
  MUX2X1 U549 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1204), .Y(n201) );
  MUX2X1 U550 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1204), .Y(n205) );
  MUX2X1 U551 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1204), .Y(n204) );
  MUX2X1 U552 ( .B(n203), .A(n200), .S(n1183), .Y(n207) );
  MUX2X1 U553 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1204), .Y(n211) );
  MUX2X1 U554 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1204), .Y(n210) );
  MUX2X1 U555 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1204), .Y(n215) );
  MUX2X1 U556 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1204), .Y(n213) );
  MUX2X1 U557 ( .B(n212), .A(n209), .S(n1183), .Y(n224) );
  MUX2X1 U558 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1205), .Y(n218) );
  MUX2X1 U559 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1205), .Y(n217) );
  MUX2X1 U560 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1205), .Y(n221) );
  MUX2X1 U561 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1205), .Y(n220) );
  MUX2X1 U562 ( .B(n219), .A(n216), .S(n1183), .Y(n223) );
  MUX2X1 U563 ( .B(n222), .A(n206), .S(n1173), .Y(n646) );
  MUX2X1 U564 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1205), .Y(n227) );
  MUX2X1 U565 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1205), .Y(n226) );
  MUX2X1 U566 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1205), .Y(n230) );
  MUX2X1 U567 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1205), .Y(n229) );
  MUX2X1 U568 ( .B(n228), .A(n225), .S(n1183), .Y(n239) );
  MUX2X1 U569 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1205), .Y(n233) );
  MUX2X1 U570 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1205), .Y(n232) );
  MUX2X1 U571 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1205), .Y(n236) );
  MUX2X1 U572 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1205), .Y(n235) );
  MUX2X1 U573 ( .B(n234), .A(n231), .S(n1183), .Y(n238) );
  MUX2X1 U574 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1206), .Y(n242) );
  MUX2X1 U575 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1206), .Y(n241) );
  MUX2X1 U576 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1206), .Y(n245) );
  MUX2X1 U577 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1206), .Y(n244) );
  MUX2X1 U578 ( .B(n243), .A(n240), .S(n1183), .Y(n254) );
  MUX2X1 U579 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1206), .Y(n248) );
  MUX2X1 U580 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1206), .Y(n247) );
  MUX2X1 U581 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1206), .Y(n251) );
  MUX2X1 U582 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1206), .Y(n250) );
  MUX2X1 U583 ( .B(n249), .A(n246), .S(n1183), .Y(n253) );
  MUX2X1 U584 ( .B(n252), .A(n237), .S(n1173), .Y(n647) );
  MUX2X1 U585 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1206), .Y(n257) );
  MUX2X1 U586 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1206), .Y(n256) );
  MUX2X1 U587 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1206), .Y(n260) );
  MUX2X1 U588 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1206), .Y(n259) );
  MUX2X1 U589 ( .B(n258), .A(n255), .S(n1182), .Y(n269) );
  MUX2X1 U590 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1207), .Y(n263) );
  MUX2X1 U591 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1207), .Y(n262) );
  MUX2X1 U592 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1207), .Y(n266) );
  MUX2X1 U593 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1207), .Y(n265) );
  MUX2X1 U594 ( .B(n264), .A(n261), .S(n1182), .Y(n268) );
  MUX2X1 U595 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1207), .Y(n272) );
  MUX2X1 U596 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1207), .Y(n271) );
  MUX2X1 U597 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1207), .Y(n275) );
  MUX2X1 U598 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1207), .Y(n274) );
  MUX2X1 U599 ( .B(n273), .A(n270), .S(n1182), .Y(n284) );
  MUX2X1 U600 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1207), .Y(n278) );
  MUX2X1 U601 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1207), .Y(n277) );
  MUX2X1 U602 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1207), .Y(n281) );
  MUX2X1 U603 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1207), .Y(n280) );
  MUX2X1 U604 ( .B(n279), .A(n276), .S(n1182), .Y(n283) );
  MUX2X1 U605 ( .B(n282), .A(n267), .S(n1173), .Y(n648) );
  MUX2X1 U606 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1208), .Y(n287) );
  MUX2X1 U607 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1208), .Y(n286) );
  MUX2X1 U608 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1208), .Y(n290) );
  MUX2X1 U609 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1208), .Y(n289) );
  MUX2X1 U610 ( .B(n288), .A(n285), .S(n1182), .Y(n299) );
  MUX2X1 U611 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1208), .Y(n293) );
  MUX2X1 U612 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1208), .Y(n292) );
  MUX2X1 U613 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1208), .Y(n296) );
  MUX2X1 U614 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1208), .Y(n295) );
  MUX2X1 U615 ( .B(n294), .A(n291), .S(n1182), .Y(n298) );
  MUX2X1 U616 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1208), .Y(n302) );
  MUX2X1 U617 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1208), .Y(n301) );
  MUX2X1 U618 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1208), .Y(n305) );
  MUX2X1 U619 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1208), .Y(n304) );
  MUX2X1 U620 ( .B(n303), .A(n300), .S(n1182), .Y(n314) );
  MUX2X1 U621 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1209), .Y(n308) );
  MUX2X1 U622 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1209), .Y(n307) );
  MUX2X1 U623 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1209), .Y(n311) );
  MUX2X1 U624 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1209), .Y(n310) );
  MUX2X1 U625 ( .B(n309), .A(n306), .S(n1182), .Y(n313) );
  MUX2X1 U626 ( .B(n312), .A(n297), .S(n1173), .Y(n649) );
  MUX2X1 U627 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1209), .Y(n317) );
  MUX2X1 U628 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1209), .Y(n316) );
  MUX2X1 U629 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1209), .Y(n320) );
  MUX2X1 U630 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1209), .Y(n319) );
  MUX2X1 U631 ( .B(n318), .A(n315), .S(n1182), .Y(n329) );
  MUX2X1 U632 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1209), .Y(n323) );
  MUX2X1 U633 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1209), .Y(n322) );
  MUX2X1 U634 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1209), .Y(n326) );
  MUX2X1 U635 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1209), .Y(n325) );
  MUX2X1 U636 ( .B(n324), .A(n321), .S(n1182), .Y(n328) );
  MUX2X1 U637 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1210), .Y(n332) );
  MUX2X1 U638 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1210), .Y(n331) );
  MUX2X1 U639 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1210), .Y(n335) );
  MUX2X1 U640 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1210), .Y(n334) );
  MUX2X1 U641 ( .B(n333), .A(n330), .S(n1182), .Y(n344) );
  MUX2X1 U642 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1210), .Y(n338) );
  MUX2X1 U643 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1210), .Y(n337) );
  MUX2X1 U644 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1210), .Y(n341) );
  MUX2X1 U645 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1210), .Y(n340) );
  MUX2X1 U646 ( .B(n339), .A(n336), .S(n1182), .Y(n343) );
  MUX2X1 U647 ( .B(n342), .A(n327), .S(n1173), .Y(n650) );
  MUX2X1 U648 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1210), .Y(n347) );
  MUX2X1 U649 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1210), .Y(n346) );
  MUX2X1 U650 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1210), .Y(n350) );
  MUX2X1 U651 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1210), .Y(n349) );
  MUX2X1 U652 ( .B(n348), .A(n345), .S(n1181), .Y(n359) );
  MUX2X1 U653 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1211), .Y(n353) );
  MUX2X1 U654 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1211), .Y(n352) );
  MUX2X1 U655 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1211), .Y(n356) );
  MUX2X1 U656 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1211), .Y(n355) );
  MUX2X1 U657 ( .B(n354), .A(n351), .S(n1181), .Y(n358) );
  MUX2X1 U658 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1211), .Y(n362) );
  MUX2X1 U659 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1211), .Y(n361) );
  MUX2X1 U660 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1211), .Y(n365) );
  MUX2X1 U661 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1211), .Y(n364) );
  MUX2X1 U662 ( .B(n363), .A(n360), .S(n1181), .Y(n374) );
  MUX2X1 U663 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1211), .Y(n368) );
  MUX2X1 U664 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1211), .Y(n367) );
  MUX2X1 U665 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1211), .Y(n371) );
  MUX2X1 U666 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1211), .Y(n370) );
  MUX2X1 U667 ( .B(n369), .A(n366), .S(n1181), .Y(n373) );
  MUX2X1 U668 ( .B(n372), .A(n357), .S(n1173), .Y(n1163) );
  MUX2X1 U669 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1212), .Y(n377) );
  MUX2X1 U670 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1212), .Y(n376) );
  MUX2X1 U671 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1212), .Y(n380) );
  MUX2X1 U672 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1212), .Y(n379) );
  MUX2X1 U673 ( .B(n378), .A(n375), .S(n1181), .Y(n389) );
  MUX2X1 U674 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1212), .Y(n383) );
  MUX2X1 U675 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1212), .Y(n382) );
  MUX2X1 U676 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1212), .Y(n386) );
  MUX2X1 U677 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1212), .Y(n385) );
  MUX2X1 U678 ( .B(n384), .A(n381), .S(n1181), .Y(n388) );
  MUX2X1 U679 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1212), .Y(n392) );
  MUX2X1 U680 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1212), .Y(n391) );
  MUX2X1 U681 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1212), .Y(n395) );
  MUX2X1 U682 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1212), .Y(n394) );
  MUX2X1 U683 ( .B(n393), .A(n390), .S(n1181), .Y(n404) );
  MUX2X1 U684 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1213), .Y(n398) );
  MUX2X1 U685 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1213), .Y(n397) );
  MUX2X1 U686 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1213), .Y(n401) );
  MUX2X1 U687 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1213), .Y(n400) );
  MUX2X1 U688 ( .B(n399), .A(n396), .S(n1181), .Y(n403) );
  MUX2X1 U689 ( .B(n402), .A(n387), .S(n1173), .Y(n1164) );
  MUX2X1 U690 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1213), .Y(n407) );
  MUX2X1 U691 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1213), .Y(n406) );
  MUX2X1 U692 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1213), .Y(n410) );
  MUX2X1 U693 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1213), .Y(n409) );
  MUX2X1 U694 ( .B(n408), .A(n405), .S(n1181), .Y(n419) );
  MUX2X1 U695 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1213), .Y(n413) );
  MUX2X1 U696 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1213), .Y(n412) );
  MUX2X1 U697 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1213), .Y(n416) );
  MUX2X1 U698 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1213), .Y(n415) );
  MUX2X1 U699 ( .B(n414), .A(n411), .S(n1181), .Y(n418) );
  MUX2X1 U700 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1214), .Y(n422) );
  MUX2X1 U701 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1214), .Y(n421) );
  MUX2X1 U702 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1214), .Y(n425) );
  MUX2X1 U703 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1214), .Y(n424) );
  MUX2X1 U704 ( .B(n423), .A(n420), .S(n1181), .Y(n434) );
  MUX2X1 U705 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1214), .Y(n428) );
  MUX2X1 U706 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1214), .Y(n427) );
  MUX2X1 U707 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1214), .Y(n431) );
  MUX2X1 U708 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1214), .Y(n430) );
  MUX2X1 U709 ( .B(n429), .A(n426), .S(n1181), .Y(n433) );
  MUX2X1 U710 ( .B(n432), .A(n417), .S(n1173), .Y(n1165) );
  MUX2X1 U711 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1214), .Y(n437) );
  MUX2X1 U712 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1214), .Y(n436) );
  MUX2X1 U713 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1214), .Y(n440) );
  MUX2X1 U714 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1214), .Y(n439) );
  MUX2X1 U715 ( .B(n438), .A(n435), .S(n1180), .Y(n449) );
  MUX2X1 U716 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1215), .Y(n443) );
  MUX2X1 U717 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1215), .Y(n442) );
  MUX2X1 U718 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1215), .Y(n446) );
  MUX2X1 U719 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1215), .Y(n445) );
  MUX2X1 U720 ( .B(n444), .A(n441), .S(n1180), .Y(n448) );
  MUX2X1 U721 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1215), .Y(n452) );
  MUX2X1 U722 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1215), .Y(n451) );
  MUX2X1 U723 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1215), .Y(n455) );
  MUX2X1 U724 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1215), .Y(n454) );
  MUX2X1 U725 ( .B(n453), .A(n450), .S(n1180), .Y(n464) );
  MUX2X1 U726 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1215), .Y(n458) );
  MUX2X1 U727 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1215), .Y(n457) );
  MUX2X1 U728 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1215), .Y(n461) );
  MUX2X1 U729 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1215), .Y(n460) );
  MUX2X1 U730 ( .B(n459), .A(n456), .S(n1180), .Y(n463) );
  MUX2X1 U731 ( .B(n462), .A(n447), .S(n1173), .Y(n1166) );
  MUX2X1 U732 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1216), .Y(n467) );
  MUX2X1 U733 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1216), .Y(n466) );
  MUX2X1 U734 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1216), .Y(n470) );
  MUX2X1 U735 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1216), .Y(n469) );
  MUX2X1 U736 ( .B(n468), .A(n465), .S(n1180), .Y(n479) );
  MUX2X1 U737 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1216), .Y(n473) );
  MUX2X1 U738 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1216), .Y(n472) );
  MUX2X1 U739 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1216), .Y(n476) );
  MUX2X1 U740 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1216), .Y(n475) );
  MUX2X1 U741 ( .B(n474), .A(n471), .S(n1180), .Y(n478) );
  MUX2X1 U742 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1216), .Y(n482) );
  MUX2X1 U743 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1216), .Y(n481) );
  MUX2X1 U744 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1216), .Y(n485) );
  MUX2X1 U745 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1216), .Y(n484) );
  MUX2X1 U746 ( .B(n483), .A(n480), .S(n1180), .Y(n494) );
  MUX2X1 U747 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1217), .Y(n488) );
  MUX2X1 U748 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1217), .Y(n487) );
  MUX2X1 U749 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1217), .Y(n491) );
  MUX2X1 U750 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1217), .Y(n490) );
  MUX2X1 U751 ( .B(n489), .A(n486), .S(n1180), .Y(n493) );
  MUX2X1 U752 ( .B(n492), .A(n477), .S(n1173), .Y(n1167) );
  MUX2X1 U753 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1217), .Y(n497) );
  MUX2X1 U754 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1217), .Y(n496) );
  MUX2X1 U755 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1217), .Y(n500) );
  MUX2X1 U756 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1217), .Y(n499) );
  MUX2X1 U757 ( .B(n498), .A(n495), .S(n1180), .Y(n509) );
  MUX2X1 U758 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1217), .Y(n503) );
  MUX2X1 U759 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1217), .Y(n502) );
  MUX2X1 U760 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1217), .Y(n506) );
  MUX2X1 U761 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1217), .Y(n505) );
  MUX2X1 U762 ( .B(n504), .A(n501), .S(n1180), .Y(n508) );
  MUX2X1 U763 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1218), .Y(n512) );
  MUX2X1 U764 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1218), .Y(n511) );
  MUX2X1 U765 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1218), .Y(n515) );
  MUX2X1 U766 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1218), .Y(n514) );
  MUX2X1 U767 ( .B(n513), .A(n510), .S(n1180), .Y(n524) );
  MUX2X1 U768 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1218), .Y(n518) );
  MUX2X1 U769 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1218), .Y(n517) );
  MUX2X1 U770 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1218), .Y(n521) );
  MUX2X1 U771 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1218), .Y(n520) );
  MUX2X1 U772 ( .B(n519), .A(n516), .S(n1180), .Y(n523) );
  MUX2X1 U773 ( .B(n522), .A(n507), .S(n1173), .Y(n1168) );
  MUX2X1 U774 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1218), .Y(n527) );
  MUX2X1 U775 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1218), .Y(n526) );
  MUX2X1 U776 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1218), .Y(n530) );
  MUX2X1 U777 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1218), .Y(n529) );
  MUX2X1 U778 ( .B(n528), .A(n525), .S(n1179), .Y(n539) );
  MUX2X1 U779 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1219), .Y(n533) );
  MUX2X1 U780 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1219), .Y(n532) );
  MUX2X1 U781 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1219), .Y(n536) );
  MUX2X1 U782 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1219), .Y(n535) );
  MUX2X1 U783 ( .B(n534), .A(n531), .S(n1179), .Y(n538) );
  MUX2X1 U784 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1219), .Y(n542) );
  MUX2X1 U785 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1219), .Y(n541) );
  MUX2X1 U786 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1219), .Y(n545) );
  MUX2X1 U787 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1219), .Y(n544) );
  MUX2X1 U788 ( .B(n543), .A(n540), .S(n1179), .Y(n554) );
  MUX2X1 U789 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1219), .Y(n548) );
  MUX2X1 U790 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1219), .Y(n547) );
  MUX2X1 U791 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1219), .Y(n551) );
  MUX2X1 U792 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1219), .Y(n550) );
  MUX2X1 U793 ( .B(n549), .A(n546), .S(n1179), .Y(n553) );
  MUX2X1 U794 ( .B(n552), .A(n537), .S(n1173), .Y(n1169) );
  MUX2X1 U795 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1220), .Y(n557) );
  MUX2X1 U796 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1220), .Y(n556) );
  MUX2X1 U797 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1220), .Y(n560) );
  MUX2X1 U798 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1220), .Y(n559) );
  MUX2X1 U799 ( .B(n558), .A(n555), .S(n1179), .Y(n569) );
  MUX2X1 U800 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1220), .Y(n563) );
  MUX2X1 U801 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1220), .Y(n562) );
  MUX2X1 U802 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1220), .Y(n566) );
  MUX2X1 U803 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1220), .Y(n565) );
  MUX2X1 U804 ( .B(n564), .A(n561), .S(n1179), .Y(n568) );
  MUX2X1 U805 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1220), .Y(n572) );
  MUX2X1 U806 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1220), .Y(n571) );
  MUX2X1 U807 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1220), .Y(n575) );
  MUX2X1 U808 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1220), .Y(n574) );
  MUX2X1 U809 ( .B(n573), .A(n570), .S(n1179), .Y(n584) );
  MUX2X1 U810 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1221), .Y(n578) );
  MUX2X1 U811 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1221), .Y(n577) );
  MUX2X1 U812 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1221), .Y(n581) );
  MUX2X1 U813 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1221), .Y(n580) );
  MUX2X1 U814 ( .B(n579), .A(n576), .S(n1179), .Y(n583) );
  MUX2X1 U815 ( .B(n582), .A(n567), .S(n1173), .Y(n1170) );
  MUX2X1 U816 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1221), .Y(n587) );
  MUX2X1 U817 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1221), .Y(n586) );
  MUX2X1 U818 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1221), .Y(n590) );
  MUX2X1 U819 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1221), .Y(n589) );
  MUX2X1 U820 ( .B(n588), .A(n585), .S(n1179), .Y(n599) );
  MUX2X1 U821 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1221), .Y(n593) );
  MUX2X1 U822 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1221), .Y(n592) );
  MUX2X1 U823 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1221), .Y(n596) );
  MUX2X1 U824 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1221), .Y(n595) );
  MUX2X1 U825 ( .B(n594), .A(n591), .S(n1179), .Y(n598) );
  MUX2X1 U826 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1222), .Y(n602) );
  MUX2X1 U827 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1222), .Y(n601) );
  MUX2X1 U828 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1222), .Y(n605) );
  MUX2X1 U829 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1222), .Y(n604) );
  MUX2X1 U830 ( .B(n603), .A(n600), .S(n1179), .Y(n614) );
  MUX2X1 U831 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1222), .Y(n608) );
  MUX2X1 U832 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1222), .Y(n607) );
  MUX2X1 U833 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1222), .Y(n611) );
  MUX2X1 U834 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1222), .Y(n610) );
  MUX2X1 U835 ( .B(n609), .A(n606), .S(n1179), .Y(n613) );
  MUX2X1 U836 ( .B(n612), .A(n597), .S(n1173), .Y(n1171) );
  MUX2X1 U837 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1222), .Y(n617) );
  MUX2X1 U838 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1222), .Y(n616) );
  MUX2X1 U839 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1222), .Y(n620) );
  MUX2X1 U840 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1222), .Y(n619) );
  MUX2X1 U841 ( .B(n618), .A(n615), .S(n1178), .Y(n629) );
  MUX2X1 U842 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1223), .Y(n623) );
  MUX2X1 U843 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1223), .Y(n622) );
  MUX2X1 U844 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1223), .Y(n626) );
  MUX2X1 U845 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1223), .Y(n625) );
  MUX2X1 U846 ( .B(n624), .A(n621), .S(n1178), .Y(n628) );
  MUX2X1 U847 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1223), .Y(n632) );
  MUX2X1 U848 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1223), .Y(n631) );
  MUX2X1 U849 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1223), .Y(n635) );
  MUX2X1 U850 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1223), .Y(n634) );
  MUX2X1 U851 ( .B(n633), .A(n630), .S(n1178), .Y(n644) );
  MUX2X1 U852 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1223), .Y(n638) );
  MUX2X1 U853 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1223), .Y(n637) );
  MUX2X1 U854 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1223), .Y(n641) );
  MUX2X1 U855 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1223), .Y(n640) );
  MUX2X1 U856 ( .B(n639), .A(n636), .S(n1178), .Y(n643) );
  MUX2X1 U857 ( .B(n642), .A(n627), .S(n1173), .Y(n1172) );
  INVX2 U858 ( .A(n77), .Y(n1224) );
  INVX2 U859 ( .A(n77), .Y(n1363) );
  INVX2 U860 ( .A(n81), .Y(n1225) );
  INVX2 U861 ( .A(n81), .Y(n1386) );
  INVX2 U862 ( .A(n79), .Y(n1226) );
  INVX2 U863 ( .A(n79), .Y(n1373) );
  INVX1 U864 ( .A(n1353), .Y(n1227) );
  BUFX2 U865 ( .A(n54), .Y(n1314) );
  BUFX2 U866 ( .A(n54), .Y(n1315) );
  BUFX2 U867 ( .A(n52), .Y(n1311) );
  BUFX2 U868 ( .A(n50), .Y(n1306) );
  BUFX2 U869 ( .A(n50), .Y(n1307) );
  BUFX2 U870 ( .A(n48), .Y(n1303) );
  BUFX2 U871 ( .A(n46), .Y(n1298) );
  BUFX2 U872 ( .A(n46), .Y(n1299) );
  BUFX2 U873 ( .A(n44), .Y(n1295) );
  BUFX2 U874 ( .A(n42), .Y(n1290) );
  BUFX2 U875 ( .A(n42), .Y(n1291) );
  BUFX2 U876 ( .A(n38), .Y(n1284) );
  BUFX2 U877 ( .A(n36), .Y(n1279) );
  BUFX2 U878 ( .A(n36), .Y(n1280) );
  BUFX2 U879 ( .A(n34), .Y(n1276) );
  INVX1 U880 ( .A(N10), .Y(n1389) );
  INVX8 U881 ( .A(n1353), .Y(n1352) );
  INVX8 U882 ( .A(n8), .Y(n1354) );
  INVX8 U883 ( .A(n8), .Y(n1355) );
  INVX8 U884 ( .A(n93), .Y(n1356) );
  INVX8 U885 ( .A(n93), .Y(n1357) );
  INVX8 U886 ( .A(n95), .Y(n1359) );
  INVX8 U887 ( .A(n95), .Y(n1360) );
  INVX8 U888 ( .A(n1224), .Y(n1361) );
  INVX8 U889 ( .A(n1363), .Y(n1362) );
  INVX8 U890 ( .A(n96), .Y(n1364) );
  INVX8 U891 ( .A(n96), .Y(n1365) );
  INVX8 U892 ( .A(n98), .Y(n1367) );
  INVX8 U893 ( .A(n98), .Y(n1368) );
  INVX8 U894 ( .A(n11), .Y(n1369) );
  INVX8 U895 ( .A(n11), .Y(n1370) );
  INVX8 U896 ( .A(n1226), .Y(n1371) );
  INVX8 U897 ( .A(n1373), .Y(n1372) );
  INVX8 U898 ( .A(n12), .Y(n1374) );
  INVX8 U899 ( .A(n12), .Y(n1375) );
  INVX8 U900 ( .A(n99), .Y(n1376) );
  INVX8 U901 ( .A(n99), .Y(n1377) );
  INVX8 U902 ( .A(n100), .Y(n1378) );
  INVX8 U903 ( .A(n100), .Y(n1379) );
  INVX8 U904 ( .A(n101), .Y(n1380) );
  INVX8 U905 ( .A(n101), .Y(n1381) );
  INVX8 U906 ( .A(n102), .Y(n1382) );
  INVX8 U907 ( .A(n102), .Y(n1383) );
  INVX8 U908 ( .A(n1225), .Y(n1384) );
  INVX8 U909 ( .A(n1386), .Y(n1385) );
  AND2X2 U910 ( .A(n2), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U911 ( .A(n7), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U912 ( .A(N30), .B(n5), .Y(\data_out<2> ) );
  AND2X2 U913 ( .A(n2), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U914 ( .A(N28), .B(n5), .Y(\data_out<4> ) );
  AND2X2 U915 ( .A(N27), .B(n2), .Y(\data_out<5> ) );
  AND2X2 U916 ( .A(n7), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U917 ( .A(N25), .B(n7), .Y(\data_out<7> ) );
  AND2X2 U918 ( .A(n7), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U919 ( .A(n7), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U920 ( .A(n2), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U921 ( .A(n7), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U922 ( .A(n7), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U923 ( .A(n2), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U924 ( .A(N18), .B(n2), .Y(\data_out<14> ) );
  AND2X2 U925 ( .A(n5), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U926 ( .A(\mem<31><0> ), .B(n1230), .Y(n1398) );
  OAI21X1 U927 ( .A(n1229), .B(n1354), .C(n1398), .Y(n2437) );
  NAND2X1 U928 ( .A(\mem<31><1> ), .B(n1230), .Y(n1399) );
  OAI21X1 U929 ( .A(n1356), .B(n1228), .C(n1399), .Y(n2436) );
  NAND2X1 U930 ( .A(\mem<31><2> ), .B(n1230), .Y(n1400) );
  OAI21X1 U931 ( .A(n1358), .B(n1228), .C(n1400), .Y(n2435) );
  NAND2X1 U932 ( .A(\mem<31><3> ), .B(n1230), .Y(n1401) );
  OAI21X1 U933 ( .A(n1360), .B(n1228), .C(n1401), .Y(n2434) );
  NAND2X1 U934 ( .A(\mem<31><4> ), .B(n1230), .Y(n1402) );
  OAI21X1 U935 ( .A(n1362), .B(n1228), .C(n1402), .Y(n2433) );
  NAND2X1 U936 ( .A(\mem<31><5> ), .B(n1230), .Y(n1403) );
  OAI21X1 U937 ( .A(n1365), .B(n1228), .C(n1403), .Y(n2432) );
  NAND2X1 U938 ( .A(\mem<31><6> ), .B(n1230), .Y(n1404) );
  OAI21X1 U939 ( .A(n1366), .B(n1228), .C(n1404), .Y(n2431) );
  NAND2X1 U940 ( .A(\mem<31><7> ), .B(n1230), .Y(n1405) );
  OAI21X1 U941 ( .A(n1367), .B(n1228), .C(n1405), .Y(n2430) );
  NAND2X1 U942 ( .A(\mem<31><8> ), .B(n1231), .Y(n1406) );
  OAI21X1 U943 ( .A(n1370), .B(n1228), .C(n1406), .Y(n2429) );
  NAND2X1 U944 ( .A(\mem<31><9> ), .B(n1231), .Y(n1407) );
  OAI21X1 U945 ( .A(n1372), .B(n1229), .C(n1407), .Y(n2428) );
  NAND2X1 U946 ( .A(\mem<31><10> ), .B(n1231), .Y(n1408) );
  OAI21X1 U947 ( .A(n1375), .B(n1229), .C(n1408), .Y(n2427) );
  NAND2X1 U948 ( .A(\mem<31><11> ), .B(n1231), .Y(n1409) );
  OAI21X1 U949 ( .A(n1376), .B(n1229), .C(n1409), .Y(n2426) );
  NAND2X1 U950 ( .A(\mem<31><12> ), .B(n1231), .Y(n1410) );
  OAI21X1 U951 ( .A(n1378), .B(n1229), .C(n1410), .Y(n2425) );
  NAND2X1 U952 ( .A(\mem<31><13> ), .B(n1231), .Y(n1411) );
  OAI21X1 U953 ( .A(n1380), .B(n1229), .C(n1411), .Y(n2424) );
  NAND2X1 U954 ( .A(\mem<31><14> ), .B(n1231), .Y(n1412) );
  OAI21X1 U955 ( .A(n1383), .B(n1229), .C(n1412), .Y(n2423) );
  NAND2X1 U956 ( .A(\mem<31><15> ), .B(n1231), .Y(n1413) );
  OAI21X1 U957 ( .A(n1385), .B(n1229), .C(n1413), .Y(n2422) );
  NAND2X1 U958 ( .A(\mem<30><0> ), .B(n1234), .Y(n1414) );
  OAI21X1 U959 ( .A(n1232), .B(n1354), .C(n1414), .Y(n2421) );
  NAND2X1 U960 ( .A(\mem<30><1> ), .B(n1234), .Y(n1415) );
  OAI21X1 U961 ( .A(n1232), .B(n1357), .C(n1415), .Y(n2420) );
  NAND2X1 U962 ( .A(\mem<30><2> ), .B(n1234), .Y(n1416) );
  OAI21X1 U963 ( .A(n1232), .B(n1358), .C(n1416), .Y(n2419) );
  NAND2X1 U964 ( .A(\mem<30><3> ), .B(n1234), .Y(n1417) );
  OAI21X1 U965 ( .A(n1232), .B(n1360), .C(n1417), .Y(n2418) );
  NAND2X1 U966 ( .A(\mem<30><4> ), .B(n1234), .Y(n1418) );
  OAI21X1 U967 ( .A(n1232), .B(n1362), .C(n1418), .Y(n2417) );
  NAND2X1 U968 ( .A(\mem<30><5> ), .B(n1234), .Y(n1419) );
  OAI21X1 U969 ( .A(n1232), .B(n1365), .C(n1419), .Y(n2416) );
  NAND2X1 U970 ( .A(\mem<30><6> ), .B(n1234), .Y(n1420) );
  OAI21X1 U971 ( .A(n1232), .B(n1366), .C(n1420), .Y(n2415) );
  NAND2X1 U972 ( .A(\mem<30><7> ), .B(n1234), .Y(n1421) );
  OAI21X1 U973 ( .A(n1232), .B(n1368), .C(n1421), .Y(n2414) );
  NAND2X1 U974 ( .A(\mem<30><8> ), .B(n1235), .Y(n1422) );
  OAI21X1 U975 ( .A(n1233), .B(n1370), .C(n1422), .Y(n2413) );
  NAND2X1 U976 ( .A(\mem<30><9> ), .B(n1235), .Y(n1423) );
  OAI21X1 U977 ( .A(n1233), .B(n1372), .C(n1423), .Y(n2412) );
  NAND2X1 U978 ( .A(\mem<30><10> ), .B(n1235), .Y(n1424) );
  OAI21X1 U979 ( .A(n1233), .B(n1375), .C(n1424), .Y(n2411) );
  NAND2X1 U980 ( .A(\mem<30><11> ), .B(n1235), .Y(n1425) );
  OAI21X1 U981 ( .A(n1233), .B(n1377), .C(n1425), .Y(n2410) );
  NAND2X1 U982 ( .A(\mem<30><12> ), .B(n1235), .Y(n1426) );
  OAI21X1 U983 ( .A(n1233), .B(n1379), .C(n1426), .Y(n2409) );
  NAND2X1 U984 ( .A(\mem<30><13> ), .B(n1235), .Y(n1427) );
  OAI21X1 U985 ( .A(n1233), .B(n1380), .C(n1427), .Y(n2408) );
  NAND2X1 U986 ( .A(\mem<30><14> ), .B(n1235), .Y(n1428) );
  OAI21X1 U987 ( .A(n1233), .B(n1382), .C(n1428), .Y(n2407) );
  NAND2X1 U988 ( .A(\mem<30><15> ), .B(n1235), .Y(n1429) );
  OAI21X1 U989 ( .A(n1233), .B(n1385), .C(n1429), .Y(n2406) );
  NAND3X1 U990 ( .A(n1388), .B(n1392), .C(n1391), .Y(n1430) );
  NAND2X1 U991 ( .A(\mem<29><0> ), .B(n1238), .Y(n1431) );
  OAI21X1 U992 ( .A(n1236), .B(n1354), .C(n1431), .Y(n2405) );
  NAND2X1 U993 ( .A(\mem<29><1> ), .B(n1238), .Y(n1432) );
  OAI21X1 U994 ( .A(n1236), .B(n1356), .C(n1432), .Y(n2404) );
  NAND2X1 U995 ( .A(\mem<29><2> ), .B(n1238), .Y(n1433) );
  OAI21X1 U996 ( .A(n1236), .B(n1358), .C(n1433), .Y(n2403) );
  NAND2X1 U997 ( .A(\mem<29><3> ), .B(n1238), .Y(n1434) );
  OAI21X1 U998 ( .A(n1236), .B(n1360), .C(n1434), .Y(n2402) );
  NAND2X1 U999 ( .A(\mem<29><4> ), .B(n1238), .Y(n1435) );
  OAI21X1 U1000 ( .A(n1236), .B(n1362), .C(n1435), .Y(n2401) );
  NAND2X1 U1001 ( .A(\mem<29><5> ), .B(n1238), .Y(n1436) );
  OAI21X1 U1002 ( .A(n1236), .B(n1365), .C(n1436), .Y(n2400) );
  NAND2X1 U1003 ( .A(\mem<29><6> ), .B(n1238), .Y(n1437) );
  OAI21X1 U1004 ( .A(n1236), .B(n1366), .C(n1437), .Y(n2399) );
  NAND2X1 U1005 ( .A(\mem<29><7> ), .B(n1238), .Y(n1438) );
  OAI21X1 U1006 ( .A(n1236), .B(n1367), .C(n1438), .Y(n2398) );
  NAND2X1 U1007 ( .A(\mem<29><8> ), .B(n1239), .Y(n1439) );
  OAI21X1 U1008 ( .A(n1237), .B(n1370), .C(n1439), .Y(n2397) );
  NAND2X1 U1009 ( .A(\mem<29><9> ), .B(n1239), .Y(n1440) );
  OAI21X1 U1010 ( .A(n1237), .B(n1372), .C(n1440), .Y(n2396) );
  NAND2X1 U1011 ( .A(\mem<29><10> ), .B(n1239), .Y(n1441) );
  OAI21X1 U1012 ( .A(n1237), .B(n1375), .C(n1441), .Y(n2395) );
  NAND2X1 U1013 ( .A(\mem<29><11> ), .B(n1239), .Y(n1442) );
  OAI21X1 U1014 ( .A(n1237), .B(n1376), .C(n1442), .Y(n2394) );
  NAND2X1 U1015 ( .A(\mem<29><12> ), .B(n1239), .Y(n1443) );
  OAI21X1 U1016 ( .A(n1237), .B(n1378), .C(n1443), .Y(n2393) );
  NAND2X1 U1017 ( .A(\mem<29><13> ), .B(n1239), .Y(n1444) );
  OAI21X1 U1018 ( .A(n1237), .B(n1381), .C(n1444), .Y(n2392) );
  NAND2X1 U1019 ( .A(\mem<29><14> ), .B(n1239), .Y(n1445) );
  OAI21X1 U1020 ( .A(n1237), .B(n1383), .C(n1445), .Y(n2391) );
  NAND2X1 U1021 ( .A(\mem<29><15> ), .B(n1239), .Y(n1446) );
  OAI21X1 U1022 ( .A(n1237), .B(n1385), .C(n1446), .Y(n2390) );
  NAND3X1 U1023 ( .A(n1392), .B(n1391), .C(n1389), .Y(n1447) );
  NAND2X1 U1024 ( .A(\mem<28><0> ), .B(n1463), .Y(n1448) );
  OAI21X1 U1025 ( .A(n1240), .B(n1354), .C(n1448), .Y(n2389) );
  NAND2X1 U1026 ( .A(\mem<28><1> ), .B(n1463), .Y(n1449) );
  OAI21X1 U1027 ( .A(n1240), .B(n1356), .C(n1449), .Y(n2388) );
  NAND2X1 U1028 ( .A(\mem<28><2> ), .B(n1463), .Y(n1450) );
  OAI21X1 U1029 ( .A(n1240), .B(n1358), .C(n1450), .Y(n2387) );
  NAND2X1 U1030 ( .A(\mem<28><3> ), .B(n1463), .Y(n1451) );
  OAI21X1 U1031 ( .A(n1240), .B(n1360), .C(n1451), .Y(n2386) );
  NAND2X1 U1032 ( .A(\mem<28><4> ), .B(n1463), .Y(n1452) );
  OAI21X1 U1033 ( .A(n1240), .B(n1362), .C(n1452), .Y(n2385) );
  NAND2X1 U1034 ( .A(\mem<28><5> ), .B(n1463), .Y(n1453) );
  OAI21X1 U1035 ( .A(n1240), .B(n1365), .C(n1453), .Y(n2384) );
  NAND2X1 U1036 ( .A(\mem<28><6> ), .B(n1463), .Y(n1454) );
  OAI21X1 U1037 ( .A(n1240), .B(n1366), .C(n1454), .Y(n2383) );
  NAND2X1 U1038 ( .A(\mem<28><7> ), .B(n1463), .Y(n1455) );
  OAI21X1 U1039 ( .A(n1240), .B(n1367), .C(n1455), .Y(n2382) );
  NAND2X1 U1040 ( .A(\mem<28><8> ), .B(n1463), .Y(n1456) );
  OAI21X1 U1041 ( .A(n1241), .B(n1370), .C(n1456), .Y(n2381) );
  NAND2X1 U1042 ( .A(\mem<28><9> ), .B(n1463), .Y(n1457) );
  OAI21X1 U1043 ( .A(n1241), .B(n1372), .C(n1457), .Y(n2380) );
  NAND2X1 U1044 ( .A(\mem<28><10> ), .B(n1463), .Y(n1458) );
  OAI21X1 U1045 ( .A(n1241), .B(n1375), .C(n1458), .Y(n2379) );
  NAND2X1 U1046 ( .A(\mem<28><11> ), .B(n1463), .Y(n1459) );
  OAI21X1 U1047 ( .A(n1241), .B(n1376), .C(n1459), .Y(n2378) );
  NAND2X1 U1048 ( .A(\mem<28><12> ), .B(n1463), .Y(n1460) );
  OAI21X1 U1049 ( .A(n1241), .B(n1378), .C(n1460), .Y(n2377) );
  NAND2X1 U1050 ( .A(\mem<28><13> ), .B(n1463), .Y(n1461) );
  OAI21X1 U1051 ( .A(n1241), .B(n1381), .C(n1461), .Y(n2376) );
  NAND2X1 U1052 ( .A(\mem<28><14> ), .B(n1463), .Y(n1462) );
  OAI21X1 U1053 ( .A(n1241), .B(n1383), .C(n1462), .Y(n2375) );
  NAND2X1 U1054 ( .A(\mem<28><15> ), .B(n1463), .Y(n1464) );
  OAI21X1 U1055 ( .A(n1241), .B(n1385), .C(n1464), .Y(n2374) );
  NAND3X1 U1056 ( .A(n1388), .B(n1390), .C(n1393), .Y(n1465) );
  NAND2X1 U1057 ( .A(\mem<27><0> ), .B(n1244), .Y(n1466) );
  OAI21X1 U1058 ( .A(n1242), .B(n1354), .C(n1466), .Y(n2373) );
  NAND2X1 U1059 ( .A(\mem<27><1> ), .B(n1244), .Y(n1467) );
  OAI21X1 U1060 ( .A(n1242), .B(n1357), .C(n1467), .Y(n2372) );
  NAND2X1 U1061 ( .A(\mem<27><2> ), .B(n1244), .Y(n1468) );
  OAI21X1 U1062 ( .A(n1242), .B(n1358), .C(n1468), .Y(n2371) );
  NAND2X1 U1063 ( .A(\mem<27><3> ), .B(n1244), .Y(n1469) );
  OAI21X1 U1064 ( .A(n1242), .B(n1360), .C(n1469), .Y(n2370) );
  NAND2X1 U1065 ( .A(\mem<27><4> ), .B(n1244), .Y(n1470) );
  OAI21X1 U1066 ( .A(n1242), .B(n1362), .C(n1470), .Y(n2369) );
  NAND2X1 U1067 ( .A(\mem<27><5> ), .B(n1244), .Y(n1471) );
  OAI21X1 U1068 ( .A(n1242), .B(n1365), .C(n1471), .Y(n2368) );
  NAND2X1 U1069 ( .A(\mem<27><6> ), .B(n1244), .Y(n1472) );
  OAI21X1 U1070 ( .A(n1242), .B(n1366), .C(n1472), .Y(n2367) );
  NAND2X1 U1071 ( .A(\mem<27><7> ), .B(n1244), .Y(n1473) );
  OAI21X1 U1072 ( .A(n1242), .B(n1368), .C(n1473), .Y(n2366) );
  NAND2X1 U1073 ( .A(\mem<27><8> ), .B(n1245), .Y(n1474) );
  OAI21X1 U1074 ( .A(n1243), .B(n1370), .C(n1474), .Y(n2365) );
  NAND2X1 U1075 ( .A(\mem<27><9> ), .B(n1245), .Y(n1475) );
  OAI21X1 U1076 ( .A(n1243), .B(n1372), .C(n1475), .Y(n2364) );
  NAND2X1 U1077 ( .A(\mem<27><10> ), .B(n1245), .Y(n1476) );
  OAI21X1 U1078 ( .A(n1243), .B(n1375), .C(n1476), .Y(n2363) );
  NAND2X1 U1079 ( .A(\mem<27><11> ), .B(n1245), .Y(n1477) );
  OAI21X1 U1080 ( .A(n1243), .B(n1377), .C(n1477), .Y(n2362) );
  NAND2X1 U1081 ( .A(\mem<27><12> ), .B(n1245), .Y(n1478) );
  OAI21X1 U1082 ( .A(n1243), .B(n1379), .C(n1478), .Y(n2361) );
  NAND2X1 U1083 ( .A(\mem<27><13> ), .B(n1245), .Y(n1479) );
  OAI21X1 U1084 ( .A(n1243), .B(n1380), .C(n1479), .Y(n2360) );
  NAND2X1 U1085 ( .A(\mem<27><14> ), .B(n1245), .Y(n1480) );
  OAI21X1 U1086 ( .A(n1243), .B(n1382), .C(n1480), .Y(n2359) );
  NAND2X1 U1087 ( .A(\mem<27><15> ), .B(n1245), .Y(n1481) );
  OAI21X1 U1088 ( .A(n1243), .B(n1385), .C(n1481), .Y(n2358) );
  NAND3X1 U1089 ( .A(n1393), .B(n1390), .C(n1389), .Y(n1482) );
  NAND2X1 U1090 ( .A(\mem<26><0> ), .B(n1248), .Y(n1483) );
  OAI21X1 U1091 ( .A(n1246), .B(n1354), .C(n1483), .Y(n2357) );
  NAND2X1 U1092 ( .A(\mem<26><1> ), .B(n1248), .Y(n1484) );
  OAI21X1 U1093 ( .A(n1246), .B(n1356), .C(n1484), .Y(n2356) );
  NAND2X1 U1094 ( .A(\mem<26><2> ), .B(n1248), .Y(n1485) );
  OAI21X1 U1095 ( .A(n1246), .B(n1358), .C(n1485), .Y(n2355) );
  NAND2X1 U1096 ( .A(\mem<26><3> ), .B(n1248), .Y(n1486) );
  OAI21X1 U1097 ( .A(n1246), .B(n1360), .C(n1486), .Y(n2354) );
  NAND2X1 U1098 ( .A(\mem<26><4> ), .B(n1248), .Y(n1487) );
  OAI21X1 U1099 ( .A(n1246), .B(n1362), .C(n1487), .Y(n2353) );
  NAND2X1 U1100 ( .A(\mem<26><5> ), .B(n1248), .Y(n1488) );
  OAI21X1 U1101 ( .A(n1246), .B(n1365), .C(n1488), .Y(n2352) );
  NAND2X1 U1102 ( .A(\mem<26><6> ), .B(n1248), .Y(n1489) );
  OAI21X1 U1103 ( .A(n1246), .B(n1366), .C(n1489), .Y(n2351) );
  NAND2X1 U1104 ( .A(\mem<26><7> ), .B(n1248), .Y(n1490) );
  OAI21X1 U1105 ( .A(n1246), .B(n1367), .C(n1490), .Y(n2350) );
  NAND2X1 U1106 ( .A(\mem<26><8> ), .B(n1249), .Y(n1491) );
  OAI21X1 U1107 ( .A(n1247), .B(n1370), .C(n1491), .Y(n2349) );
  NAND2X1 U1108 ( .A(\mem<26><9> ), .B(n1249), .Y(n1492) );
  OAI21X1 U1109 ( .A(n1247), .B(n1372), .C(n1492), .Y(n2348) );
  NAND2X1 U1110 ( .A(\mem<26><10> ), .B(n1249), .Y(n1493) );
  OAI21X1 U1111 ( .A(n1247), .B(n1375), .C(n1493), .Y(n2347) );
  NAND2X1 U1112 ( .A(\mem<26><11> ), .B(n1249), .Y(n1494) );
  OAI21X1 U1113 ( .A(n1247), .B(n1376), .C(n1494), .Y(n2346) );
  NAND2X1 U1114 ( .A(\mem<26><12> ), .B(n1249), .Y(n1495) );
  OAI21X1 U1115 ( .A(n1247), .B(n1378), .C(n1495), .Y(n2345) );
  NAND2X1 U1116 ( .A(\mem<26><13> ), .B(n1249), .Y(n1496) );
  OAI21X1 U1117 ( .A(n1247), .B(n1381), .C(n1496), .Y(n2344) );
  NAND2X1 U1118 ( .A(\mem<26><14> ), .B(n1249), .Y(n1497) );
  OAI21X1 U1119 ( .A(n1247), .B(n1383), .C(n1497), .Y(n2343) );
  NAND2X1 U1120 ( .A(\mem<26><15> ), .B(n1249), .Y(n1498) );
  OAI21X1 U1121 ( .A(n1247), .B(n1385), .C(n1498), .Y(n2342) );
  NAND3X1 U1122 ( .A(n1388), .B(n1393), .C(n1391), .Y(n1499) );
  NAND2X1 U1123 ( .A(\mem<25><0> ), .B(n1252), .Y(n1500) );
  OAI21X1 U1124 ( .A(n1250), .B(n1354), .C(n1500), .Y(n2341) );
  NAND2X1 U1125 ( .A(\mem<25><1> ), .B(n1252), .Y(n1501) );
  OAI21X1 U1126 ( .A(n1250), .B(n1357), .C(n1501), .Y(n2340) );
  NAND2X1 U1127 ( .A(\mem<25><2> ), .B(n1252), .Y(n1502) );
  OAI21X1 U1128 ( .A(n1250), .B(n1358), .C(n1502), .Y(n2339) );
  NAND2X1 U1129 ( .A(\mem<25><3> ), .B(n1252), .Y(n1503) );
  OAI21X1 U1130 ( .A(n1250), .B(n1360), .C(n1503), .Y(n2338) );
  NAND2X1 U1131 ( .A(\mem<25><4> ), .B(n1252), .Y(n1504) );
  OAI21X1 U1132 ( .A(n1250), .B(n1362), .C(n1504), .Y(n2337) );
  NAND2X1 U1133 ( .A(\mem<25><5> ), .B(n1252), .Y(n1505) );
  OAI21X1 U1134 ( .A(n1250), .B(n1365), .C(n1505), .Y(n2336) );
  NAND2X1 U1135 ( .A(\mem<25><6> ), .B(n1252), .Y(n1506) );
  OAI21X1 U1136 ( .A(n1250), .B(n1366), .C(n1506), .Y(n2335) );
  NAND2X1 U1137 ( .A(\mem<25><7> ), .B(n1252), .Y(n1507) );
  OAI21X1 U1138 ( .A(n1250), .B(n1368), .C(n1507), .Y(n2334) );
  NAND2X1 U1139 ( .A(\mem<25><8> ), .B(n1253), .Y(n1508) );
  OAI21X1 U1140 ( .A(n1251), .B(n1370), .C(n1508), .Y(n2333) );
  NAND2X1 U1141 ( .A(\mem<25><9> ), .B(n1253), .Y(n1509) );
  OAI21X1 U1142 ( .A(n1251), .B(n1372), .C(n1509), .Y(n2332) );
  NAND2X1 U1143 ( .A(\mem<25><10> ), .B(n1253), .Y(n1510) );
  OAI21X1 U1144 ( .A(n1251), .B(n1375), .C(n1510), .Y(n2331) );
  NAND2X1 U1145 ( .A(\mem<25><11> ), .B(n1253), .Y(n1511) );
  OAI21X1 U1146 ( .A(n1251), .B(n1377), .C(n1511), .Y(n2330) );
  NAND2X1 U1147 ( .A(\mem<25><12> ), .B(n1253), .Y(n1512) );
  OAI21X1 U1148 ( .A(n1251), .B(n1379), .C(n1512), .Y(n2329) );
  NAND2X1 U1149 ( .A(\mem<25><13> ), .B(n1253), .Y(n1513) );
  OAI21X1 U1150 ( .A(n1251), .B(n1380), .C(n1513), .Y(n2328) );
  NAND2X1 U1151 ( .A(\mem<25><14> ), .B(n1253), .Y(n1514) );
  OAI21X1 U1152 ( .A(n1251), .B(n1382), .C(n1514), .Y(n2327) );
  NAND2X1 U1153 ( .A(\mem<25><15> ), .B(n1253), .Y(n1515) );
  OAI21X1 U1154 ( .A(n1251), .B(n1385), .C(n1515), .Y(n2326) );
  NOR3X1 U1155 ( .A(n1388), .B(n1390), .C(n1392), .Y(n1909) );
  NAND2X1 U1156 ( .A(\mem<24><0> ), .B(n1255), .Y(n1516) );
  OAI21X1 U1157 ( .A(n1254), .B(n1354), .C(n1516), .Y(n2325) );
  NAND2X1 U1158 ( .A(\mem<24><1> ), .B(n1256), .Y(n1517) );
  OAI21X1 U1159 ( .A(n1254), .B(n1357), .C(n1517), .Y(n2324) );
  NAND2X1 U1160 ( .A(\mem<24><2> ), .B(n1255), .Y(n1518) );
  OAI21X1 U1161 ( .A(n1254), .B(n1358), .C(n1518), .Y(n2323) );
  NAND2X1 U1162 ( .A(\mem<24><3> ), .B(n1), .Y(n1519) );
  OAI21X1 U1163 ( .A(n1254), .B(n1360), .C(n1519), .Y(n2322) );
  NAND2X1 U1164 ( .A(\mem<24><4> ), .B(n1256), .Y(n1520) );
  OAI21X1 U1165 ( .A(n1254), .B(n1362), .C(n1520), .Y(n2321) );
  NAND2X1 U1166 ( .A(\mem<24><5> ), .B(n1255), .Y(n1521) );
  OAI21X1 U1167 ( .A(n1254), .B(n1365), .C(n1521), .Y(n2320) );
  NAND2X1 U1168 ( .A(\mem<24><6> ), .B(n1), .Y(n1522) );
  OAI21X1 U1169 ( .A(n1254), .B(n1366), .C(n1522), .Y(n2319) );
  NAND2X1 U1170 ( .A(\mem<24><7> ), .B(n1256), .Y(n1523) );
  OAI21X1 U1171 ( .A(n1254), .B(n1368), .C(n1523), .Y(n2318) );
  NAND2X1 U1172 ( .A(\mem<24><8> ), .B(n1255), .Y(n1524) );
  OAI21X1 U1173 ( .A(n1254), .B(n1370), .C(n1524), .Y(n2317) );
  NAND2X1 U1174 ( .A(\mem<24><9> ), .B(n1), .Y(n1525) );
  OAI21X1 U1175 ( .A(n1254), .B(n1372), .C(n1525), .Y(n2316) );
  NAND2X1 U1177 ( .A(\mem<24><10> ), .B(n1256), .Y(n1526) );
  OAI21X1 U1178 ( .A(n1254), .B(n1375), .C(n1526), .Y(n2315) );
  NAND2X1 U1179 ( .A(\mem<24><11> ), .B(n1255), .Y(n1527) );
  OAI21X1 U1180 ( .A(n1254), .B(n1377), .C(n1527), .Y(n2314) );
  NAND2X1 U1181 ( .A(\mem<24><12> ), .B(n1), .Y(n1528) );
  OAI21X1 U1182 ( .A(n1254), .B(n1379), .C(n1528), .Y(n2313) );
  NAND2X1 U1183 ( .A(\mem<24><13> ), .B(n1256), .Y(n1529) );
  OAI21X1 U1184 ( .A(n1254), .B(n1381), .C(n1529), .Y(n2312) );
  NAND2X1 U1185 ( .A(\mem<24><14> ), .B(n1255), .Y(n1530) );
  OAI21X1 U1186 ( .A(n1254), .B(n1382), .C(n1530), .Y(n2311) );
  NAND2X1 U1187 ( .A(\mem<24><15> ), .B(n1), .Y(n1531) );
  OAI21X1 U1188 ( .A(n1254), .B(n1385), .C(n1531), .Y(n2310) );
  NAND2X1 U1189 ( .A(\mem<23><0> ), .B(n1259), .Y(n1532) );
  OAI21X1 U1190 ( .A(n1257), .B(n1354), .C(n1532), .Y(n2309) );
  NAND2X1 U1191 ( .A(\mem<23><1> ), .B(n1259), .Y(n1533) );
  OAI21X1 U1192 ( .A(n1257), .B(n1357), .C(n1533), .Y(n2308) );
  NAND2X1 U1193 ( .A(\mem<23><2> ), .B(n1259), .Y(n1534) );
  OAI21X1 U1194 ( .A(n1257), .B(n1358), .C(n1534), .Y(n2307) );
  NAND2X1 U1195 ( .A(\mem<23><3> ), .B(n1259), .Y(n1535) );
  OAI21X1 U1196 ( .A(n1257), .B(n1360), .C(n1535), .Y(n2306) );
  NAND2X1 U1197 ( .A(\mem<23><4> ), .B(n1259), .Y(n1536) );
  OAI21X1 U1198 ( .A(n1257), .B(n1361), .C(n1536), .Y(n2305) );
  NAND2X1 U1199 ( .A(\mem<23><5> ), .B(n1259), .Y(n1537) );
  OAI21X1 U1200 ( .A(n1257), .B(n1364), .C(n1537), .Y(n2304) );
  NAND2X1 U1201 ( .A(\mem<23><6> ), .B(n1259), .Y(n1538) );
  OAI21X1 U1202 ( .A(n1257), .B(n1366), .C(n1538), .Y(n2303) );
  NAND2X1 U1203 ( .A(\mem<23><7> ), .B(n1259), .Y(n1539) );
  OAI21X1 U1204 ( .A(n1257), .B(n1368), .C(n1539), .Y(n2302) );
  NAND2X1 U1205 ( .A(\mem<23><8> ), .B(n1260), .Y(n1540) );
  OAI21X1 U1206 ( .A(n1258), .B(n1370), .C(n1540), .Y(n2301) );
  NAND2X1 U1207 ( .A(\mem<23><9> ), .B(n1260), .Y(n1541) );
  OAI21X1 U1208 ( .A(n1258), .B(n1372), .C(n1541), .Y(n2300) );
  NAND2X1 U1209 ( .A(\mem<23><10> ), .B(n1260), .Y(n1542) );
  OAI21X1 U1210 ( .A(n1258), .B(n1375), .C(n1542), .Y(n2299) );
  NAND2X1 U1211 ( .A(\mem<23><11> ), .B(n1260), .Y(n1543) );
  OAI21X1 U1212 ( .A(n1258), .B(n1377), .C(n1543), .Y(n2298) );
  NAND2X1 U1213 ( .A(\mem<23><12> ), .B(n1260), .Y(n1544) );
  OAI21X1 U1214 ( .A(n1258), .B(n1379), .C(n1544), .Y(n2297) );
  NAND2X1 U1215 ( .A(\mem<23><13> ), .B(n1260), .Y(n1545) );
  OAI21X1 U1216 ( .A(n1258), .B(n1381), .C(n1545), .Y(n2296) );
  NAND2X1 U1217 ( .A(\mem<23><14> ), .B(n1260), .Y(n1546) );
  OAI21X1 U1218 ( .A(n1258), .B(n1383), .C(n1546), .Y(n2295) );
  NAND2X1 U1219 ( .A(\mem<23><15> ), .B(n1260), .Y(n1547) );
  OAI21X1 U1220 ( .A(n1258), .B(n1385), .C(n1547), .Y(n2294) );
  NAND2X1 U1221 ( .A(\mem<22><0> ), .B(n1263), .Y(n1548) );
  OAI21X1 U1222 ( .A(n1261), .B(n1354), .C(n1548), .Y(n2293) );
  NAND2X1 U1223 ( .A(\mem<22><1> ), .B(n1263), .Y(n1549) );
  OAI21X1 U1224 ( .A(n1261), .B(n1357), .C(n1549), .Y(n2292) );
  NAND2X1 U1225 ( .A(\mem<22><2> ), .B(n1263), .Y(n1550) );
  OAI21X1 U1226 ( .A(n1261), .B(n1358), .C(n1550), .Y(n2291) );
  NAND2X1 U1227 ( .A(\mem<22><3> ), .B(n1263), .Y(n1551) );
  OAI21X1 U1228 ( .A(n1261), .B(n1360), .C(n1551), .Y(n2290) );
  NAND2X1 U1229 ( .A(\mem<22><4> ), .B(n1263), .Y(n1552) );
  OAI21X1 U1230 ( .A(n1261), .B(n1361), .C(n1552), .Y(n2289) );
  NAND2X1 U1231 ( .A(\mem<22><5> ), .B(n1263), .Y(n1553) );
  OAI21X1 U1232 ( .A(n1261), .B(n1364), .C(n1553), .Y(n2288) );
  NAND2X1 U1233 ( .A(\mem<22><6> ), .B(n1263), .Y(n1554) );
  OAI21X1 U1234 ( .A(n1261), .B(n1366), .C(n1554), .Y(n2287) );
  NAND2X1 U1235 ( .A(\mem<22><7> ), .B(n1263), .Y(n1555) );
  OAI21X1 U1236 ( .A(n1261), .B(n1368), .C(n1555), .Y(n2286) );
  NAND2X1 U1237 ( .A(\mem<22><8> ), .B(n1264), .Y(n1556) );
  OAI21X1 U1238 ( .A(n1262), .B(n1370), .C(n1556), .Y(n2285) );
  NAND2X1 U1239 ( .A(\mem<22><9> ), .B(n1264), .Y(n1557) );
  OAI21X1 U1240 ( .A(n1262), .B(n1372), .C(n1557), .Y(n2284) );
  NAND2X1 U1241 ( .A(\mem<22><10> ), .B(n1264), .Y(n1558) );
  OAI21X1 U1242 ( .A(n1262), .B(n1375), .C(n1558), .Y(n2283) );
  NAND2X1 U1243 ( .A(\mem<22><11> ), .B(n1264), .Y(n1559) );
  OAI21X1 U1244 ( .A(n1262), .B(n1376), .C(n1559), .Y(n2282) );
  NAND2X1 U1245 ( .A(\mem<22><12> ), .B(n1264), .Y(n1560) );
  OAI21X1 U1246 ( .A(n1262), .B(n1378), .C(n1560), .Y(n2281) );
  NAND2X1 U1247 ( .A(\mem<22><13> ), .B(n1264), .Y(n1561) );
  OAI21X1 U1248 ( .A(n1262), .B(n1381), .C(n1561), .Y(n2280) );
  NAND2X1 U1249 ( .A(\mem<22><14> ), .B(n1264), .Y(n1562) );
  OAI21X1 U1250 ( .A(n1262), .B(n1383), .C(n1562), .Y(n2279) );
  NAND2X1 U1251 ( .A(\mem<22><15> ), .B(n1264), .Y(n1563) );
  OAI21X1 U1252 ( .A(n1262), .B(n1385), .C(n1563), .Y(n2278) );
  NAND2X1 U1253 ( .A(\mem<21><0> ), .B(n1267), .Y(n1564) );
  OAI21X1 U1254 ( .A(n1265), .B(n1354), .C(n1564), .Y(n2277) );
  NAND2X1 U1255 ( .A(\mem<21><1> ), .B(n1267), .Y(n1565) );
  OAI21X1 U1256 ( .A(n1265), .B(n1357), .C(n1565), .Y(n2276) );
  NAND2X1 U1257 ( .A(\mem<21><2> ), .B(n1267), .Y(n1566) );
  OAI21X1 U1258 ( .A(n1265), .B(n1358), .C(n1566), .Y(n2275) );
  NAND2X1 U1259 ( .A(\mem<21><3> ), .B(n1267), .Y(n1567) );
  OAI21X1 U1260 ( .A(n1265), .B(n1360), .C(n1567), .Y(n2274) );
  NAND2X1 U1261 ( .A(\mem<21><4> ), .B(n1267), .Y(n1568) );
  OAI21X1 U1262 ( .A(n1265), .B(n1361), .C(n1568), .Y(n2273) );
  NAND2X1 U1263 ( .A(\mem<21><5> ), .B(n1267), .Y(n1569) );
  OAI21X1 U1264 ( .A(n1265), .B(n1364), .C(n1569), .Y(n2272) );
  NAND2X1 U1265 ( .A(\mem<21><6> ), .B(n1267), .Y(n1570) );
  OAI21X1 U1266 ( .A(n1265), .B(n1366), .C(n1570), .Y(n2271) );
  NAND2X1 U1267 ( .A(\mem<21><7> ), .B(n1267), .Y(n1571) );
  OAI21X1 U1268 ( .A(n1265), .B(n1368), .C(n1571), .Y(n2270) );
  NAND2X1 U1269 ( .A(\mem<21><8> ), .B(n1268), .Y(n1572) );
  OAI21X1 U1270 ( .A(n1266), .B(n1370), .C(n1572), .Y(n2269) );
  NAND2X1 U1271 ( .A(\mem<21><9> ), .B(n1268), .Y(n1573) );
  OAI21X1 U1272 ( .A(n1266), .B(n1372), .C(n1573), .Y(n2268) );
  NAND2X1 U1273 ( .A(\mem<21><10> ), .B(n1268), .Y(n1574) );
  OAI21X1 U1274 ( .A(n1266), .B(n1375), .C(n1574), .Y(n2267) );
  NAND2X1 U1275 ( .A(\mem<21><11> ), .B(n1268), .Y(n1575) );
  OAI21X1 U1276 ( .A(n1266), .B(n1377), .C(n1575), .Y(n2266) );
  NAND2X1 U1277 ( .A(\mem<21><12> ), .B(n1268), .Y(n1576) );
  OAI21X1 U1278 ( .A(n1266), .B(n1379), .C(n1576), .Y(n2265) );
  NAND2X1 U1279 ( .A(\mem<21><13> ), .B(n1268), .Y(n1577) );
  OAI21X1 U1280 ( .A(n1266), .B(n1381), .C(n1577), .Y(n2264) );
  NAND2X1 U1281 ( .A(\mem<21><14> ), .B(n1268), .Y(n1578) );
  OAI21X1 U1282 ( .A(n1266), .B(n1383), .C(n1578), .Y(n2263) );
  NAND2X1 U1283 ( .A(\mem<21><15> ), .B(n1268), .Y(n1579) );
  OAI21X1 U1284 ( .A(n1266), .B(n1385), .C(n1579), .Y(n2262) );
  NAND2X1 U1285 ( .A(\mem<20><0> ), .B(n1271), .Y(n1580) );
  OAI21X1 U1286 ( .A(n1269), .B(n1354), .C(n1580), .Y(n2261) );
  NAND2X1 U1287 ( .A(\mem<20><1> ), .B(n1271), .Y(n1581) );
  OAI21X1 U1288 ( .A(n1269), .B(n1357), .C(n1581), .Y(n2260) );
  NAND2X1 U1289 ( .A(\mem<20><2> ), .B(n1271), .Y(n1582) );
  OAI21X1 U1290 ( .A(n1269), .B(n1358), .C(n1582), .Y(n2259) );
  NAND2X1 U1291 ( .A(\mem<20><3> ), .B(n1271), .Y(n1583) );
  OAI21X1 U1292 ( .A(n1269), .B(n1360), .C(n1583), .Y(n2258) );
  NAND2X1 U1293 ( .A(\mem<20><4> ), .B(n1271), .Y(n1584) );
  OAI21X1 U1294 ( .A(n1269), .B(n1361), .C(n1584), .Y(n2257) );
  NAND2X1 U1295 ( .A(\mem<20><5> ), .B(n1271), .Y(n1585) );
  OAI21X1 U1296 ( .A(n1269), .B(n1364), .C(n1585), .Y(n2256) );
  NAND2X1 U1297 ( .A(\mem<20><6> ), .B(n1271), .Y(n1586) );
  OAI21X1 U1298 ( .A(n1269), .B(n1366), .C(n1586), .Y(n2255) );
  NAND2X1 U1299 ( .A(\mem<20><7> ), .B(n1271), .Y(n1587) );
  OAI21X1 U1300 ( .A(n1269), .B(n1368), .C(n1587), .Y(n2254) );
  NAND2X1 U1301 ( .A(\mem<20><8> ), .B(n1272), .Y(n1588) );
  OAI21X1 U1302 ( .A(n1270), .B(n1370), .C(n1588), .Y(n2253) );
  NAND2X1 U1303 ( .A(\mem<20><9> ), .B(n1272), .Y(n1589) );
  OAI21X1 U1304 ( .A(n1270), .B(n1372), .C(n1589), .Y(n2252) );
  NAND2X1 U1305 ( .A(\mem<20><10> ), .B(n1272), .Y(n1590) );
  OAI21X1 U1306 ( .A(n1270), .B(n1375), .C(n1590), .Y(n2251) );
  NAND2X1 U1307 ( .A(\mem<20><11> ), .B(n1272), .Y(n1591) );
  OAI21X1 U1308 ( .A(n1270), .B(n1377), .C(n1591), .Y(n2250) );
  NAND2X1 U1309 ( .A(\mem<20><12> ), .B(n1272), .Y(n1592) );
  OAI21X1 U1310 ( .A(n1270), .B(n1379), .C(n1592), .Y(n2249) );
  NAND2X1 U1311 ( .A(\mem<20><13> ), .B(n1272), .Y(n1593) );
  OAI21X1 U1312 ( .A(n1270), .B(n1381), .C(n1593), .Y(n2248) );
  NAND2X1 U1313 ( .A(\mem<20><14> ), .B(n1272), .Y(n1594) );
  OAI21X1 U1314 ( .A(n1270), .B(n1383), .C(n1594), .Y(n2247) );
  NAND2X1 U1315 ( .A(\mem<20><15> ), .B(n1272), .Y(n1595) );
  OAI21X1 U1316 ( .A(n1270), .B(n1385), .C(n1595), .Y(n2246) );
  NAND2X1 U1317 ( .A(\mem<19><0> ), .B(n1275), .Y(n1596) );
  OAI21X1 U1318 ( .A(n1273), .B(n1355), .C(n1596), .Y(n2245) );
  NAND2X1 U1319 ( .A(\mem<19><1> ), .B(n1275), .Y(n1597) );
  OAI21X1 U1320 ( .A(n1273), .B(n1357), .C(n1597), .Y(n2244) );
  NAND2X1 U1321 ( .A(\mem<19><2> ), .B(n1275), .Y(n1598) );
  OAI21X1 U1322 ( .A(n1273), .B(n1358), .C(n1598), .Y(n2243) );
  NAND2X1 U1323 ( .A(\mem<19><3> ), .B(n1275), .Y(n1599) );
  OAI21X1 U1324 ( .A(n1273), .B(n1360), .C(n1599), .Y(n2242) );
  NAND2X1 U1325 ( .A(\mem<19><4> ), .B(n1275), .Y(n1600) );
  OAI21X1 U1326 ( .A(n1273), .B(n1361), .C(n1600), .Y(n2241) );
  NAND2X1 U1327 ( .A(\mem<19><5> ), .B(n1275), .Y(n1601) );
  OAI21X1 U1328 ( .A(n1273), .B(n1364), .C(n1601), .Y(n2240) );
  NAND2X1 U1329 ( .A(\mem<19><6> ), .B(n1275), .Y(n1602) );
  OAI21X1 U1330 ( .A(n1273), .B(n1366), .C(n1602), .Y(n2239) );
  NAND2X1 U1331 ( .A(\mem<19><7> ), .B(n1275), .Y(n1603) );
  OAI21X1 U1332 ( .A(n1273), .B(n1368), .C(n1603), .Y(n2238) );
  NAND2X1 U1333 ( .A(\mem<19><8> ), .B(n1276), .Y(n1604) );
  OAI21X1 U1334 ( .A(n1274), .B(n1370), .C(n1604), .Y(n2237) );
  NAND2X1 U1335 ( .A(\mem<19><9> ), .B(n1276), .Y(n1605) );
  OAI21X1 U1336 ( .A(n1274), .B(n1372), .C(n1605), .Y(n2236) );
  NAND2X1 U1337 ( .A(\mem<19><10> ), .B(n1276), .Y(n1606) );
  OAI21X1 U1338 ( .A(n1274), .B(n1375), .C(n1606), .Y(n2235) );
  NAND2X1 U1339 ( .A(\mem<19><11> ), .B(n1276), .Y(n1607) );
  OAI21X1 U1340 ( .A(n1274), .B(n1376), .C(n1607), .Y(n2234) );
  NAND2X1 U1341 ( .A(\mem<19><12> ), .B(n1276), .Y(n1608) );
  OAI21X1 U1342 ( .A(n1274), .B(n1378), .C(n1608), .Y(n2233) );
  NAND2X1 U1343 ( .A(\mem<19><13> ), .B(n1276), .Y(n1609) );
  OAI21X1 U1344 ( .A(n1274), .B(n1381), .C(n1609), .Y(n2232) );
  NAND2X1 U1345 ( .A(\mem<19><14> ), .B(n1276), .Y(n1610) );
  OAI21X1 U1346 ( .A(n1274), .B(n1383), .C(n1610), .Y(n2231) );
  NAND2X1 U1347 ( .A(\mem<19><15> ), .B(n1276), .Y(n1611) );
  OAI21X1 U1348 ( .A(n1274), .B(n1385), .C(n1611), .Y(n2230) );
  NAND2X1 U1349 ( .A(\mem<18><0> ), .B(n1279), .Y(n1612) );
  OAI21X1 U1350 ( .A(n1277), .B(n1355), .C(n1612), .Y(n2229) );
  NAND2X1 U1351 ( .A(\mem<18><1> ), .B(n1279), .Y(n1613) );
  OAI21X1 U1352 ( .A(n1277), .B(n1357), .C(n1613), .Y(n2228) );
  NAND2X1 U1353 ( .A(\mem<18><2> ), .B(n1279), .Y(n1614) );
  OAI21X1 U1354 ( .A(n1277), .B(n1358), .C(n1614), .Y(n2227) );
  NAND2X1 U1355 ( .A(\mem<18><3> ), .B(n1279), .Y(n1615) );
  OAI21X1 U1356 ( .A(n1277), .B(n1359), .C(n1615), .Y(n2226) );
  NAND2X1 U1357 ( .A(\mem<18><4> ), .B(n1279), .Y(n1616) );
  OAI21X1 U1358 ( .A(n1277), .B(n1361), .C(n1616), .Y(n2225) );
  NAND2X1 U1359 ( .A(\mem<18><5> ), .B(n1279), .Y(n1617) );
  OAI21X1 U1360 ( .A(n1277), .B(n1364), .C(n1617), .Y(n2224) );
  NAND2X1 U1361 ( .A(\mem<18><6> ), .B(n1279), .Y(n1618) );
  OAI21X1 U1362 ( .A(n1277), .B(n1366), .C(n1618), .Y(n2223) );
  NAND2X1 U1363 ( .A(\mem<18><7> ), .B(n1279), .Y(n1619) );
  OAI21X1 U1364 ( .A(n1277), .B(n1368), .C(n1619), .Y(n2222) );
  NAND2X1 U1365 ( .A(\mem<18><8> ), .B(n1280), .Y(n1620) );
  OAI21X1 U1366 ( .A(n1278), .B(n1369), .C(n1620), .Y(n2221) );
  NAND2X1 U1367 ( .A(\mem<18><9> ), .B(n1280), .Y(n1621) );
  OAI21X1 U1368 ( .A(n1278), .B(n1371), .C(n1621), .Y(n2220) );
  NAND2X1 U1369 ( .A(\mem<18><10> ), .B(n1280), .Y(n1622) );
  OAI21X1 U1370 ( .A(n1278), .B(n1374), .C(n1622), .Y(n2219) );
  NAND2X1 U1371 ( .A(\mem<18><11> ), .B(n1280), .Y(n1623) );
  OAI21X1 U1372 ( .A(n1278), .B(n1376), .C(n1623), .Y(n2218) );
  NAND2X1 U1373 ( .A(\mem<18><12> ), .B(n1280), .Y(n1624) );
  OAI21X1 U1374 ( .A(n1278), .B(n1378), .C(n1624), .Y(n2217) );
  NAND2X1 U1375 ( .A(\mem<18><13> ), .B(n1280), .Y(n1625) );
  OAI21X1 U1376 ( .A(n1278), .B(n1381), .C(n1625), .Y(n2216) );
  NAND2X1 U1377 ( .A(\mem<18><14> ), .B(n1280), .Y(n1626) );
  OAI21X1 U1378 ( .A(n1278), .B(n1383), .C(n1626), .Y(n2215) );
  NAND2X1 U1379 ( .A(\mem<18><15> ), .B(n1280), .Y(n1627) );
  OAI21X1 U1380 ( .A(n1278), .B(n1384), .C(n1627), .Y(n2214) );
  NAND2X1 U1381 ( .A(\mem<17><0> ), .B(n1283), .Y(n1628) );
  OAI21X1 U1382 ( .A(n1281), .B(n1355), .C(n1628), .Y(n2213) );
  NAND2X1 U1383 ( .A(\mem<17><1> ), .B(n1283), .Y(n1629) );
  OAI21X1 U1384 ( .A(n1281), .B(n1357), .C(n1629), .Y(n2212) );
  NAND2X1 U1385 ( .A(\mem<17><2> ), .B(n1283), .Y(n1630) );
  OAI21X1 U1386 ( .A(n1281), .B(n1358), .C(n1630), .Y(n2211) );
  NAND2X1 U1387 ( .A(\mem<17><3> ), .B(n1283), .Y(n1631) );
  OAI21X1 U1388 ( .A(n1281), .B(n1360), .C(n1631), .Y(n2210) );
  NAND2X1 U1389 ( .A(\mem<17><4> ), .B(n1283), .Y(n1632) );
  OAI21X1 U1390 ( .A(n1281), .B(n1361), .C(n1632), .Y(n2209) );
  NAND2X1 U1391 ( .A(\mem<17><5> ), .B(n1283), .Y(n1633) );
  OAI21X1 U1392 ( .A(n1281), .B(n1364), .C(n1633), .Y(n2208) );
  NAND2X1 U1393 ( .A(\mem<17><6> ), .B(n1283), .Y(n1634) );
  OAI21X1 U1394 ( .A(n1281), .B(n1366), .C(n1634), .Y(n2207) );
  NAND2X1 U1395 ( .A(\mem<17><7> ), .B(n1283), .Y(n1635) );
  OAI21X1 U1396 ( .A(n1281), .B(n1368), .C(n1635), .Y(n2206) );
  NAND2X1 U1397 ( .A(\mem<17><8> ), .B(n1284), .Y(n1636) );
  OAI21X1 U1398 ( .A(n1282), .B(n1370), .C(n1636), .Y(n2205) );
  NAND2X1 U1399 ( .A(\mem<17><9> ), .B(n1284), .Y(n1637) );
  OAI21X1 U1400 ( .A(n1282), .B(n1372), .C(n1637), .Y(n2204) );
  NAND2X1 U1401 ( .A(\mem<17><10> ), .B(n1284), .Y(n1638) );
  OAI21X1 U1402 ( .A(n1282), .B(n1375), .C(n1638), .Y(n2203) );
  NAND2X1 U1403 ( .A(\mem<17><11> ), .B(n1284), .Y(n1639) );
  OAI21X1 U1404 ( .A(n1282), .B(n1377), .C(n1639), .Y(n2202) );
  NAND2X1 U1405 ( .A(\mem<17><12> ), .B(n1284), .Y(n1640) );
  OAI21X1 U1406 ( .A(n1282), .B(n1379), .C(n1640), .Y(n2201) );
  NAND2X1 U1407 ( .A(\mem<17><13> ), .B(n1284), .Y(n1641) );
  OAI21X1 U1408 ( .A(n1282), .B(n1381), .C(n1641), .Y(n2200) );
  NAND2X1 U1409 ( .A(\mem<17><14> ), .B(n1284), .Y(n1642) );
  OAI21X1 U1410 ( .A(n1282), .B(n1383), .C(n1642), .Y(n2199) );
  NAND2X1 U1411 ( .A(\mem<17><15> ), .B(n1284), .Y(n1643) );
  OAI21X1 U1412 ( .A(n1282), .B(n1385), .C(n1643), .Y(n2198) );
  NAND2X1 U1413 ( .A(\mem<16><0> ), .B(n1286), .Y(n1644) );
  OAI21X1 U1414 ( .A(n1285), .B(n1355), .C(n1644), .Y(n2197) );
  NAND2X1 U1415 ( .A(\mem<16><1> ), .B(n1286), .Y(n1645) );
  OAI21X1 U1416 ( .A(n1285), .B(n1357), .C(n1645), .Y(n2196) );
  NAND2X1 U1417 ( .A(\mem<16><2> ), .B(n1286), .Y(n1646) );
  OAI21X1 U1418 ( .A(n1285), .B(n1358), .C(n1646), .Y(n2195) );
  NAND2X1 U1419 ( .A(\mem<16><3> ), .B(n1286), .Y(n1647) );
  OAI21X1 U1420 ( .A(n1285), .B(n1359), .C(n1647), .Y(n2194) );
  NAND2X1 U1421 ( .A(\mem<16><4> ), .B(n1286), .Y(n1648) );
  OAI21X1 U1422 ( .A(n1285), .B(n1361), .C(n1648), .Y(n2193) );
  NAND2X1 U1423 ( .A(\mem<16><5> ), .B(n1286), .Y(n1649) );
  OAI21X1 U1424 ( .A(n1285), .B(n1364), .C(n1649), .Y(n2192) );
  NAND2X1 U1425 ( .A(\mem<16><6> ), .B(n1286), .Y(n1650) );
  OAI21X1 U1426 ( .A(n1285), .B(n1366), .C(n1650), .Y(n2191) );
  NAND2X1 U1427 ( .A(\mem<16><7> ), .B(n1286), .Y(n1651) );
  OAI21X1 U1428 ( .A(n1285), .B(n1368), .C(n1651), .Y(n2190) );
  NAND2X1 U1429 ( .A(\mem<16><8> ), .B(n1287), .Y(n1652) );
  OAI21X1 U1430 ( .A(n1285), .B(n1369), .C(n1652), .Y(n2189) );
  NAND2X1 U1431 ( .A(\mem<16><9> ), .B(n1287), .Y(n1653) );
  OAI21X1 U1432 ( .A(n1285), .B(n1371), .C(n1653), .Y(n2188) );
  NAND2X1 U1433 ( .A(\mem<16><10> ), .B(n1287), .Y(n1654) );
  OAI21X1 U1434 ( .A(n1285), .B(n1374), .C(n1654), .Y(n2187) );
  NAND2X1 U1435 ( .A(\mem<16><11> ), .B(n1287), .Y(n1655) );
  OAI21X1 U1436 ( .A(n1285), .B(n1377), .C(n1655), .Y(n2186) );
  NAND2X1 U1437 ( .A(\mem<16><12> ), .B(n1287), .Y(n1656) );
  OAI21X1 U1438 ( .A(n1285), .B(n1379), .C(n1656), .Y(n2185) );
  NAND2X1 U1439 ( .A(\mem<16><13> ), .B(n1287), .Y(n1657) );
  OAI21X1 U1440 ( .A(n1285), .B(n1381), .C(n1657), .Y(n2184) );
  NAND2X1 U1441 ( .A(\mem<16><14> ), .B(n1287), .Y(n1658) );
  OAI21X1 U1442 ( .A(n1285), .B(n1383), .C(n1658), .Y(n2183) );
  NAND2X1 U1443 ( .A(\mem<16><15> ), .B(n1287), .Y(n1659) );
  OAI21X1 U1444 ( .A(n1285), .B(n1384), .C(n1659), .Y(n2182) );
  NAND3X1 U1445 ( .A(n1394), .B(n2438), .C(n1397), .Y(n1660) );
  NAND2X1 U1446 ( .A(\mem<15><0> ), .B(n1290), .Y(n1661) );
  OAI21X1 U1447 ( .A(n1288), .B(n1354), .C(n1661), .Y(n2181) );
  NAND2X1 U1448 ( .A(\mem<15><1> ), .B(n1290), .Y(n1662) );
  OAI21X1 U1449 ( .A(n1288), .B(n1357), .C(n1662), .Y(n2180) );
  NAND2X1 U1450 ( .A(\mem<15><2> ), .B(n1290), .Y(n1663) );
  OAI21X1 U1451 ( .A(n1288), .B(n1358), .C(n1663), .Y(n2179) );
  NAND2X1 U1452 ( .A(\mem<15><3> ), .B(n1290), .Y(n1664) );
  OAI21X1 U1453 ( .A(n1288), .B(n1359), .C(n1664), .Y(n2178) );
  NAND2X1 U1454 ( .A(\mem<15><4> ), .B(n1290), .Y(n1665) );
  OAI21X1 U1455 ( .A(n1288), .B(n1361), .C(n1665), .Y(n2177) );
  NAND2X1 U1456 ( .A(\mem<15><5> ), .B(n1290), .Y(n1666) );
  OAI21X1 U1457 ( .A(n1288), .B(n1364), .C(n1666), .Y(n2176) );
  NAND2X1 U1458 ( .A(\mem<15><6> ), .B(n1290), .Y(n1667) );
  OAI21X1 U1459 ( .A(n1288), .B(n1366), .C(n1667), .Y(n2175) );
  NAND2X1 U1460 ( .A(\mem<15><7> ), .B(n1290), .Y(n1668) );
  OAI21X1 U1461 ( .A(n1288), .B(n1368), .C(n1668), .Y(n2174) );
  NAND2X1 U1462 ( .A(\mem<15><8> ), .B(n1291), .Y(n1669) );
  OAI21X1 U1463 ( .A(n1289), .B(n1369), .C(n1669), .Y(n2173) );
  NAND2X1 U1464 ( .A(\mem<15><9> ), .B(n1291), .Y(n1670) );
  OAI21X1 U1465 ( .A(n1289), .B(n1371), .C(n1670), .Y(n2172) );
  NAND2X1 U1466 ( .A(\mem<15><10> ), .B(n1291), .Y(n1671) );
  OAI21X1 U1467 ( .A(n1289), .B(n1374), .C(n1671), .Y(n2171) );
  NAND2X1 U1468 ( .A(\mem<15><11> ), .B(n1291), .Y(n1672) );
  OAI21X1 U1469 ( .A(n1289), .B(n1376), .C(n1672), .Y(n2170) );
  NAND2X1 U1470 ( .A(\mem<15><12> ), .B(n1291), .Y(n1673) );
  OAI21X1 U1471 ( .A(n1289), .B(n1378), .C(n1673), .Y(n2169) );
  NAND2X1 U1472 ( .A(\mem<15><13> ), .B(n1291), .Y(n1674) );
  OAI21X1 U1473 ( .A(n1289), .B(n1381), .C(n1674), .Y(n2168) );
  NAND2X1 U1474 ( .A(\mem<15><14> ), .B(n1291), .Y(n1675) );
  OAI21X1 U1475 ( .A(n1289), .B(n1383), .C(n1675), .Y(n2167) );
  NAND2X1 U1476 ( .A(\mem<15><15> ), .B(n1291), .Y(n1676) );
  OAI21X1 U1477 ( .A(n1289), .B(n1384), .C(n1676), .Y(n2166) );
  NAND2X1 U1478 ( .A(\mem<14><0> ), .B(n1294), .Y(n1677) );
  OAI21X1 U1479 ( .A(n1292), .B(n1355), .C(n1677), .Y(n2165) );
  NAND2X1 U1480 ( .A(\mem<14><1> ), .B(n1294), .Y(n1678) );
  OAI21X1 U1481 ( .A(n1292), .B(n1357), .C(n1678), .Y(n2164) );
  NAND2X1 U1482 ( .A(\mem<14><2> ), .B(n1294), .Y(n1679) );
  OAI21X1 U1483 ( .A(n1292), .B(n1358), .C(n1679), .Y(n2163) );
  NAND2X1 U1484 ( .A(\mem<14><3> ), .B(n1294), .Y(n1680) );
  OAI21X1 U1485 ( .A(n1292), .B(n1360), .C(n1680), .Y(n2162) );
  NAND2X1 U1486 ( .A(\mem<14><4> ), .B(n1294), .Y(n1681) );
  OAI21X1 U1487 ( .A(n1292), .B(n1361), .C(n1681), .Y(n2161) );
  NAND2X1 U1488 ( .A(\mem<14><5> ), .B(n1294), .Y(n1682) );
  OAI21X1 U1489 ( .A(n1292), .B(n1364), .C(n1682), .Y(n2160) );
  NAND2X1 U1490 ( .A(\mem<14><6> ), .B(n1294), .Y(n1683) );
  OAI21X1 U1491 ( .A(n1292), .B(n1366), .C(n1683), .Y(n2159) );
  NAND2X1 U1492 ( .A(\mem<14><7> ), .B(n1294), .Y(n1684) );
  OAI21X1 U1493 ( .A(n1292), .B(n1368), .C(n1684), .Y(n2158) );
  NAND2X1 U1494 ( .A(\mem<14><8> ), .B(n1295), .Y(n1685) );
  OAI21X1 U1495 ( .A(n1293), .B(n1370), .C(n1685), .Y(n2157) );
  NAND2X1 U1496 ( .A(\mem<14><9> ), .B(n1295), .Y(n1686) );
  OAI21X1 U1497 ( .A(n1293), .B(n1372), .C(n1686), .Y(n2156) );
  NAND2X1 U1498 ( .A(\mem<14><10> ), .B(n1295), .Y(n1687) );
  OAI21X1 U1499 ( .A(n1293), .B(n1375), .C(n1687), .Y(n2155) );
  NAND2X1 U1500 ( .A(\mem<14><11> ), .B(n1295), .Y(n1688) );
  OAI21X1 U1501 ( .A(n1293), .B(n1377), .C(n1688), .Y(n2154) );
  NAND2X1 U1502 ( .A(\mem<14><12> ), .B(n1295), .Y(n1689) );
  OAI21X1 U1503 ( .A(n1293), .B(n1379), .C(n1689), .Y(n2153) );
  NAND2X1 U1504 ( .A(\mem<14><13> ), .B(n1295), .Y(n1690) );
  OAI21X1 U1505 ( .A(n1293), .B(n1381), .C(n1690), .Y(n2152) );
  NAND2X1 U1506 ( .A(\mem<14><14> ), .B(n1295), .Y(n1691) );
  OAI21X1 U1507 ( .A(n1293), .B(n1383), .C(n1691), .Y(n2151) );
  NAND2X1 U1508 ( .A(\mem<14><15> ), .B(n1295), .Y(n1692) );
  OAI21X1 U1509 ( .A(n1293), .B(n1385), .C(n1692), .Y(n2150) );
  NAND2X1 U1510 ( .A(\mem<13><0> ), .B(n1298), .Y(n1693) );
  OAI21X1 U1511 ( .A(n1296), .B(n1354), .C(n1693), .Y(n2149) );
  NAND2X1 U1512 ( .A(\mem<13><1> ), .B(n1298), .Y(n1694) );
  OAI21X1 U1513 ( .A(n1296), .B(n1357), .C(n1694), .Y(n2148) );
  NAND2X1 U1514 ( .A(\mem<13><2> ), .B(n1298), .Y(n1695) );
  OAI21X1 U1515 ( .A(n1296), .B(n1358), .C(n1695), .Y(n2147) );
  NAND2X1 U1516 ( .A(\mem<13><3> ), .B(n1298), .Y(n1696) );
  OAI21X1 U1517 ( .A(n1296), .B(n1359), .C(n1696), .Y(n2146) );
  NAND2X1 U1518 ( .A(\mem<13><4> ), .B(n1298), .Y(n1697) );
  OAI21X1 U1519 ( .A(n1296), .B(n1361), .C(n1697), .Y(n2145) );
  NAND2X1 U1520 ( .A(\mem<13><5> ), .B(n1298), .Y(n1698) );
  OAI21X1 U1521 ( .A(n1296), .B(n1364), .C(n1698), .Y(n2144) );
  NAND2X1 U1522 ( .A(\mem<13><6> ), .B(n1298), .Y(n1699) );
  OAI21X1 U1523 ( .A(n1296), .B(n1366), .C(n1699), .Y(n2143) );
  NAND2X1 U1524 ( .A(\mem<13><7> ), .B(n1298), .Y(n1700) );
  OAI21X1 U1525 ( .A(n1296), .B(n1368), .C(n1700), .Y(n2142) );
  NAND2X1 U1526 ( .A(\mem<13><8> ), .B(n1299), .Y(n1701) );
  OAI21X1 U1527 ( .A(n1297), .B(n1369), .C(n1701), .Y(n2141) );
  NAND2X1 U1528 ( .A(\mem<13><9> ), .B(n1299), .Y(n1702) );
  OAI21X1 U1529 ( .A(n1297), .B(n1371), .C(n1702), .Y(n2140) );
  NAND2X1 U1530 ( .A(\mem<13><10> ), .B(n1299), .Y(n1703) );
  OAI21X1 U1531 ( .A(n1297), .B(n1374), .C(n1703), .Y(n2139) );
  NAND2X1 U1532 ( .A(\mem<13><11> ), .B(n1299), .Y(n1704) );
  OAI21X1 U1533 ( .A(n1297), .B(n1377), .C(n1704), .Y(n2138) );
  NAND2X1 U1534 ( .A(\mem<13><12> ), .B(n1299), .Y(n1705) );
  OAI21X1 U1535 ( .A(n1297), .B(n1379), .C(n1705), .Y(n2137) );
  NAND2X1 U1536 ( .A(\mem<13><13> ), .B(n1299), .Y(n1706) );
  OAI21X1 U1537 ( .A(n1297), .B(n1381), .C(n1706), .Y(n2136) );
  NAND2X1 U1538 ( .A(\mem<13><14> ), .B(n1299), .Y(n1707) );
  OAI21X1 U1539 ( .A(n1297), .B(n1383), .C(n1707), .Y(n2135) );
  NAND2X1 U1540 ( .A(\mem<13><15> ), .B(n1299), .Y(n1708) );
  OAI21X1 U1541 ( .A(n1297), .B(n1384), .C(n1708), .Y(n2134) );
  NAND2X1 U1542 ( .A(\mem<12><0> ), .B(n1302), .Y(n1709) );
  OAI21X1 U1543 ( .A(n1300), .B(n1355), .C(n1709), .Y(n2133) );
  NAND2X1 U1544 ( .A(\mem<12><1> ), .B(n1302), .Y(n1710) );
  OAI21X1 U1545 ( .A(n1300), .B(n1357), .C(n1710), .Y(n2132) );
  NAND2X1 U1546 ( .A(\mem<12><2> ), .B(n1302), .Y(n1711) );
  OAI21X1 U1547 ( .A(n1300), .B(n1358), .C(n1711), .Y(n2131) );
  NAND2X1 U1548 ( .A(\mem<12><3> ), .B(n1302), .Y(n1712) );
  OAI21X1 U1549 ( .A(n1300), .B(n1360), .C(n1712), .Y(n2130) );
  NAND2X1 U1550 ( .A(\mem<12><4> ), .B(n1302), .Y(n1713) );
  OAI21X1 U1551 ( .A(n1300), .B(n1361), .C(n1713), .Y(n2129) );
  NAND2X1 U1552 ( .A(\mem<12><5> ), .B(n1302), .Y(n1714) );
  OAI21X1 U1553 ( .A(n1300), .B(n1364), .C(n1714), .Y(n2128) );
  NAND2X1 U1554 ( .A(\mem<12><6> ), .B(n1302), .Y(n1715) );
  OAI21X1 U1555 ( .A(n1300), .B(n1366), .C(n1715), .Y(n2127) );
  NAND2X1 U1556 ( .A(\mem<12><7> ), .B(n1302), .Y(n1716) );
  OAI21X1 U1557 ( .A(n1300), .B(n1368), .C(n1716), .Y(n2126) );
  NAND2X1 U1558 ( .A(\mem<12><8> ), .B(n1303), .Y(n1717) );
  OAI21X1 U1559 ( .A(n1301), .B(n1370), .C(n1717), .Y(n2125) );
  NAND2X1 U1560 ( .A(\mem<12><9> ), .B(n1303), .Y(n1718) );
  OAI21X1 U1561 ( .A(n1301), .B(n1372), .C(n1718), .Y(n2124) );
  NAND2X1 U1562 ( .A(\mem<12><10> ), .B(n1303), .Y(n1719) );
  OAI21X1 U1563 ( .A(n1301), .B(n1375), .C(n1719), .Y(n2123) );
  NAND2X1 U1564 ( .A(\mem<12><11> ), .B(n1303), .Y(n1720) );
  OAI21X1 U1565 ( .A(n1301), .B(n1376), .C(n1720), .Y(n2122) );
  NAND2X1 U1566 ( .A(\mem<12><12> ), .B(n1303), .Y(n1721) );
  OAI21X1 U1567 ( .A(n1301), .B(n1378), .C(n1721), .Y(n2121) );
  NAND2X1 U1568 ( .A(\mem<12><13> ), .B(n1303), .Y(n1722) );
  OAI21X1 U1569 ( .A(n1301), .B(n1381), .C(n1722), .Y(n2120) );
  NAND2X1 U1570 ( .A(\mem<12><14> ), .B(n1303), .Y(n1723) );
  OAI21X1 U1571 ( .A(n1301), .B(n1383), .C(n1723), .Y(n2119) );
  NAND2X1 U1572 ( .A(\mem<12><15> ), .B(n1303), .Y(n1724) );
  OAI21X1 U1573 ( .A(n1301), .B(n1385), .C(n1724), .Y(n2118) );
  NAND2X1 U1574 ( .A(\mem<11><0> ), .B(n1306), .Y(n1725) );
  OAI21X1 U1575 ( .A(n1304), .B(n1354), .C(n1725), .Y(n2117) );
  NAND2X1 U1576 ( .A(\mem<11><1> ), .B(n1306), .Y(n1726) );
  OAI21X1 U1577 ( .A(n1304), .B(n1356), .C(n1726), .Y(n2116) );
  NAND2X1 U1578 ( .A(\mem<11><2> ), .B(n1306), .Y(n1727) );
  OAI21X1 U1579 ( .A(n1304), .B(n1358), .C(n1727), .Y(n2115) );
  NAND2X1 U1580 ( .A(\mem<11><3> ), .B(n1306), .Y(n1728) );
  OAI21X1 U1581 ( .A(n1304), .B(n1359), .C(n1728), .Y(n2114) );
  NAND2X1 U1582 ( .A(\mem<11><4> ), .B(n1306), .Y(n1729) );
  OAI21X1 U1583 ( .A(n1304), .B(n1362), .C(n1729), .Y(n2113) );
  NAND2X1 U1584 ( .A(\mem<11><5> ), .B(n1306), .Y(n1730) );
  OAI21X1 U1585 ( .A(n1304), .B(n1365), .C(n1730), .Y(n2112) );
  NAND2X1 U1586 ( .A(\mem<11><6> ), .B(n1306), .Y(n1731) );
  OAI21X1 U1587 ( .A(n1304), .B(n1366), .C(n1731), .Y(n2111) );
  NAND2X1 U1588 ( .A(\mem<11><7> ), .B(n1306), .Y(n1732) );
  OAI21X1 U1589 ( .A(n1304), .B(n1367), .C(n1732), .Y(n2110) );
  NAND2X1 U1590 ( .A(\mem<11><8> ), .B(n1307), .Y(n1733) );
  OAI21X1 U1591 ( .A(n1305), .B(n1369), .C(n1733), .Y(n2109) );
  NAND2X1 U1592 ( .A(\mem<11><9> ), .B(n1307), .Y(n1734) );
  OAI21X1 U1593 ( .A(n1305), .B(n1371), .C(n1734), .Y(n2108) );
  NAND2X1 U1594 ( .A(\mem<11><10> ), .B(n1307), .Y(n1735) );
  OAI21X1 U1595 ( .A(n1305), .B(n1374), .C(n1735), .Y(n2107) );
  NAND2X1 U1596 ( .A(\mem<11><11> ), .B(n1307), .Y(n1736) );
  OAI21X1 U1597 ( .A(n1305), .B(n1376), .C(n1736), .Y(n2106) );
  NAND2X1 U1598 ( .A(\mem<11><12> ), .B(n1307), .Y(n1737) );
  OAI21X1 U1599 ( .A(n1305), .B(n1378), .C(n1737), .Y(n2105) );
  NAND2X1 U1600 ( .A(\mem<11><13> ), .B(n1307), .Y(n1738) );
  OAI21X1 U1601 ( .A(n1305), .B(n1380), .C(n1738), .Y(n2104) );
  NAND2X1 U1602 ( .A(\mem<11><14> ), .B(n1307), .Y(n1739) );
  OAI21X1 U1603 ( .A(n1305), .B(n1382), .C(n1739), .Y(n2103) );
  NAND2X1 U1604 ( .A(\mem<11><15> ), .B(n1307), .Y(n1740) );
  OAI21X1 U1605 ( .A(n1305), .B(n1384), .C(n1740), .Y(n2102) );
  NAND2X1 U1606 ( .A(\mem<10><0> ), .B(n1310), .Y(n1741) );
  OAI21X1 U1607 ( .A(n1308), .B(n1355), .C(n1741), .Y(n2101) );
  NAND2X1 U1608 ( .A(\mem<10><1> ), .B(n1310), .Y(n1742) );
  OAI21X1 U1609 ( .A(n1308), .B(n1356), .C(n1742), .Y(n2100) );
  NAND2X1 U1610 ( .A(\mem<10><2> ), .B(n1310), .Y(n1743) );
  OAI21X1 U1611 ( .A(n1308), .B(n1358), .C(n1743), .Y(n2099) );
  NAND2X1 U1612 ( .A(\mem<10><3> ), .B(n1310), .Y(n1744) );
  OAI21X1 U1613 ( .A(n1308), .B(n1359), .C(n1744), .Y(n2098) );
  NAND2X1 U1614 ( .A(\mem<10><4> ), .B(n1310), .Y(n1745) );
  OAI21X1 U1615 ( .A(n1308), .B(n1362), .C(n1745), .Y(n2097) );
  NAND2X1 U1616 ( .A(\mem<10><5> ), .B(n1310), .Y(n1746) );
  OAI21X1 U1617 ( .A(n1308), .B(n1365), .C(n1746), .Y(n2096) );
  NAND2X1 U1618 ( .A(\mem<10><6> ), .B(n1310), .Y(n1747) );
  OAI21X1 U1619 ( .A(n1308), .B(n1366), .C(n1747), .Y(n2095) );
  NAND2X1 U1620 ( .A(\mem<10><7> ), .B(n1310), .Y(n1748) );
  OAI21X1 U1621 ( .A(n1308), .B(n1367), .C(n1748), .Y(n2094) );
  NAND2X1 U1622 ( .A(\mem<10><8> ), .B(n1311), .Y(n1749) );
  OAI21X1 U1623 ( .A(n1309), .B(n1369), .C(n1749), .Y(n2093) );
  NAND2X1 U1624 ( .A(\mem<10><9> ), .B(n1311), .Y(n1750) );
  OAI21X1 U1625 ( .A(n1309), .B(n1371), .C(n1750), .Y(n2092) );
  NAND2X1 U1626 ( .A(\mem<10><10> ), .B(n1311), .Y(n1751) );
  OAI21X1 U1627 ( .A(n1309), .B(n1374), .C(n1751), .Y(n2091) );
  NAND2X1 U1628 ( .A(\mem<10><11> ), .B(n1311), .Y(n1752) );
  OAI21X1 U1629 ( .A(n1309), .B(n1377), .C(n1752), .Y(n2090) );
  NAND2X1 U1630 ( .A(\mem<10><12> ), .B(n1311), .Y(n1753) );
  OAI21X1 U1631 ( .A(n1309), .B(n1379), .C(n1753), .Y(n2089) );
  NAND2X1 U1632 ( .A(\mem<10><13> ), .B(n1311), .Y(n1754) );
  OAI21X1 U1633 ( .A(n1309), .B(n1380), .C(n1754), .Y(n2088) );
  NAND2X1 U1634 ( .A(\mem<10><14> ), .B(n1311), .Y(n1755) );
  OAI21X1 U1635 ( .A(n1309), .B(n1382), .C(n1755), .Y(n2087) );
  NAND2X1 U1636 ( .A(\mem<10><15> ), .B(n1311), .Y(n1756) );
  OAI21X1 U1637 ( .A(n1309), .B(n1384), .C(n1756), .Y(n2086) );
  NAND2X1 U1638 ( .A(\mem<9><0> ), .B(n1314), .Y(n1757) );
  OAI21X1 U1639 ( .A(n1312), .B(n1355), .C(n1757), .Y(n2085) );
  NAND2X1 U1640 ( .A(\mem<9><1> ), .B(n1314), .Y(n1758) );
  OAI21X1 U1641 ( .A(n1312), .B(n1356), .C(n1758), .Y(n2084) );
  NAND2X1 U1642 ( .A(\mem<9><2> ), .B(n1314), .Y(n1759) );
  OAI21X1 U1643 ( .A(n1312), .B(n1358), .C(n1759), .Y(n2083) );
  NAND2X1 U1644 ( .A(\mem<9><3> ), .B(n1314), .Y(n1760) );
  OAI21X1 U1645 ( .A(n1312), .B(n1359), .C(n1760), .Y(n2082) );
  NAND2X1 U1646 ( .A(\mem<9><4> ), .B(n1314), .Y(n1761) );
  OAI21X1 U1647 ( .A(n1312), .B(n1362), .C(n1761), .Y(n2081) );
  NAND2X1 U1648 ( .A(\mem<9><5> ), .B(n1314), .Y(n1762) );
  OAI21X1 U1649 ( .A(n1312), .B(n1365), .C(n1762), .Y(n2080) );
  NAND2X1 U1650 ( .A(\mem<9><6> ), .B(n1314), .Y(n1763) );
  OAI21X1 U1651 ( .A(n1312), .B(n1366), .C(n1763), .Y(n2079) );
  NAND2X1 U1652 ( .A(\mem<9><7> ), .B(n1314), .Y(n1764) );
  OAI21X1 U1653 ( .A(n1312), .B(n1367), .C(n1764), .Y(n2078) );
  NAND2X1 U1654 ( .A(\mem<9><8> ), .B(n1315), .Y(n1765) );
  OAI21X1 U1655 ( .A(n1313), .B(n1369), .C(n1765), .Y(n2077) );
  NAND2X1 U1656 ( .A(\mem<9><9> ), .B(n1315), .Y(n1766) );
  OAI21X1 U1657 ( .A(n1313), .B(n1371), .C(n1766), .Y(n2076) );
  NAND2X1 U1658 ( .A(\mem<9><10> ), .B(n1315), .Y(n1767) );
  OAI21X1 U1659 ( .A(n1313), .B(n1374), .C(n1767), .Y(n2075) );
  NAND2X1 U1660 ( .A(\mem<9><11> ), .B(n1315), .Y(n1768) );
  OAI21X1 U1661 ( .A(n1313), .B(n1376), .C(n1768), .Y(n2074) );
  NAND2X1 U1662 ( .A(\mem<9><12> ), .B(n1315), .Y(n1769) );
  OAI21X1 U1663 ( .A(n1313), .B(n1378), .C(n1769), .Y(n2073) );
  NAND2X1 U1664 ( .A(\mem<9><13> ), .B(n1315), .Y(n1770) );
  OAI21X1 U1665 ( .A(n1313), .B(n1380), .C(n1770), .Y(n2072) );
  NAND2X1 U1666 ( .A(\mem<9><14> ), .B(n1315), .Y(n1771) );
  OAI21X1 U1667 ( .A(n1313), .B(n1382), .C(n1771), .Y(n2071) );
  NAND2X1 U1668 ( .A(\mem<9><15> ), .B(n1315), .Y(n1772) );
  OAI21X1 U1669 ( .A(n1313), .B(n1384), .C(n1772), .Y(n2070) );
  NAND2X1 U1670 ( .A(\mem<8><0> ), .B(n1317), .Y(n1774) );
  OAI21X1 U1671 ( .A(n1316), .B(n1354), .C(n1774), .Y(n2069) );
  NAND2X1 U1672 ( .A(\mem<8><1> ), .B(n1317), .Y(n1775) );
  OAI21X1 U1673 ( .A(n1316), .B(n1356), .C(n1775), .Y(n2068) );
  NAND2X1 U1674 ( .A(\mem<8><2> ), .B(n1317), .Y(n1776) );
  OAI21X1 U1675 ( .A(n1316), .B(n1358), .C(n1776), .Y(n2067) );
  NAND2X1 U1676 ( .A(\mem<8><3> ), .B(n1317), .Y(n1777) );
  OAI21X1 U1677 ( .A(n1316), .B(n1359), .C(n1777), .Y(n2066) );
  NAND2X1 U1678 ( .A(\mem<8><4> ), .B(n1317), .Y(n1778) );
  OAI21X1 U1679 ( .A(n1316), .B(n1362), .C(n1778), .Y(n2065) );
  NAND2X1 U1680 ( .A(\mem<8><5> ), .B(n1317), .Y(n1779) );
  OAI21X1 U1681 ( .A(n1316), .B(n1365), .C(n1779), .Y(n2064) );
  NAND2X1 U1682 ( .A(\mem<8><6> ), .B(n1317), .Y(n1780) );
  OAI21X1 U1683 ( .A(n1316), .B(n1366), .C(n1780), .Y(n2063) );
  NAND2X1 U1684 ( .A(\mem<8><7> ), .B(n1317), .Y(n1781) );
  OAI21X1 U1685 ( .A(n1316), .B(n1367), .C(n1781), .Y(n2062) );
  NAND2X1 U1686 ( .A(\mem<8><8> ), .B(n1318), .Y(n1782) );
  OAI21X1 U1687 ( .A(n1316), .B(n1369), .C(n1782), .Y(n2061) );
  NAND2X1 U1688 ( .A(\mem<8><9> ), .B(n1318), .Y(n1783) );
  OAI21X1 U1689 ( .A(n1316), .B(n1371), .C(n1783), .Y(n2060) );
  NAND2X1 U1690 ( .A(\mem<8><10> ), .B(n1318), .Y(n1784) );
  OAI21X1 U1691 ( .A(n1316), .B(n1374), .C(n1784), .Y(n2059) );
  NAND2X1 U1692 ( .A(\mem<8><11> ), .B(n1318), .Y(n1785) );
  OAI21X1 U1693 ( .A(n1316), .B(n1376), .C(n1785), .Y(n2058) );
  NAND2X1 U1694 ( .A(\mem<8><12> ), .B(n1318), .Y(n1786) );
  OAI21X1 U1695 ( .A(n1316), .B(n1378), .C(n1786), .Y(n2057) );
  NAND2X1 U1696 ( .A(\mem<8><13> ), .B(n1318), .Y(n1787) );
  OAI21X1 U1697 ( .A(n1316), .B(n1380), .C(n1787), .Y(n2056) );
  NAND2X1 U1698 ( .A(\mem<8><14> ), .B(n1318), .Y(n1788) );
  OAI21X1 U1699 ( .A(n1316), .B(n1382), .C(n1788), .Y(n2055) );
  NAND2X1 U1700 ( .A(\mem<8><15> ), .B(n1318), .Y(n1789) );
  OAI21X1 U1701 ( .A(n1316), .B(n1384), .C(n1789), .Y(n2054) );
  NAND3X1 U1702 ( .A(n1395), .B(n2438), .C(n1397), .Y(n1790) );
  NAND2X1 U1703 ( .A(\mem<7><0> ), .B(n1321), .Y(n1791) );
  OAI21X1 U1704 ( .A(n1319), .B(n1355), .C(n1791), .Y(n2053) );
  NAND2X1 U1705 ( .A(\mem<7><1> ), .B(n1321), .Y(n1792) );
  OAI21X1 U1706 ( .A(n1319), .B(n1356), .C(n1792), .Y(n2052) );
  NAND2X1 U1707 ( .A(\mem<7><2> ), .B(n1321), .Y(n1793) );
  OAI21X1 U1708 ( .A(n1319), .B(n1358), .C(n1793), .Y(n2051) );
  NAND2X1 U1709 ( .A(\mem<7><3> ), .B(n1321), .Y(n1794) );
  OAI21X1 U1710 ( .A(n1319), .B(n1359), .C(n1794), .Y(n2050) );
  NAND2X1 U1711 ( .A(\mem<7><4> ), .B(n1321), .Y(n1795) );
  OAI21X1 U1712 ( .A(n1319), .B(n1362), .C(n1795), .Y(n2049) );
  NAND2X1 U1713 ( .A(\mem<7><5> ), .B(n1321), .Y(n1796) );
  OAI21X1 U1714 ( .A(n1319), .B(n1364), .C(n1796), .Y(n2048) );
  NAND2X1 U1715 ( .A(\mem<7><6> ), .B(n1321), .Y(n1797) );
  OAI21X1 U1716 ( .A(n1319), .B(n1366), .C(n1797), .Y(n2047) );
  NAND2X1 U1717 ( .A(\mem<7><7> ), .B(n1321), .Y(n1798) );
  OAI21X1 U1718 ( .A(n1319), .B(n1367), .C(n1798), .Y(n2046) );
  NAND2X1 U1719 ( .A(\mem<7><8> ), .B(n1322), .Y(n1799) );
  OAI21X1 U1720 ( .A(n1320), .B(n1369), .C(n1799), .Y(n2045) );
  NAND2X1 U1721 ( .A(\mem<7><9> ), .B(n1322), .Y(n1800) );
  OAI21X1 U1722 ( .A(n1320), .B(n1371), .C(n1800), .Y(n2044) );
  NAND2X1 U1723 ( .A(\mem<7><10> ), .B(n1322), .Y(n1801) );
  OAI21X1 U1724 ( .A(n1320), .B(n1374), .C(n1801), .Y(n2043) );
  NAND2X1 U1725 ( .A(\mem<7><11> ), .B(n1322), .Y(n1802) );
  OAI21X1 U1726 ( .A(n1320), .B(n1377), .C(n1802), .Y(n2042) );
  NAND2X1 U1727 ( .A(\mem<7><12> ), .B(n1322), .Y(n1803) );
  OAI21X1 U1728 ( .A(n1320), .B(n1379), .C(n1803), .Y(n2041) );
  NAND2X1 U1729 ( .A(\mem<7><13> ), .B(n1322), .Y(n1804) );
  OAI21X1 U1730 ( .A(n1320), .B(n1380), .C(n1804), .Y(n2040) );
  NAND2X1 U1731 ( .A(\mem<7><14> ), .B(n1322), .Y(n1805) );
  OAI21X1 U1732 ( .A(n1320), .B(n1382), .C(n1805), .Y(n2039) );
  NAND2X1 U1733 ( .A(\mem<7><15> ), .B(n1322), .Y(n1806) );
  OAI21X1 U1734 ( .A(n1320), .B(n1384), .C(n1806), .Y(n2038) );
  NAND2X1 U1735 ( .A(\mem<6><0> ), .B(n1325), .Y(n1807) );
  OAI21X1 U1736 ( .A(n1323), .B(n1355), .C(n1807), .Y(n2037) );
  NAND2X1 U1737 ( .A(\mem<6><1> ), .B(n1325), .Y(n1808) );
  OAI21X1 U1738 ( .A(n1323), .B(n1356), .C(n1808), .Y(n2036) );
  NAND2X1 U1739 ( .A(\mem<6><2> ), .B(n1325), .Y(n1809) );
  OAI21X1 U1740 ( .A(n1323), .B(n1358), .C(n1809), .Y(n2035) );
  NAND2X1 U1741 ( .A(\mem<6><3> ), .B(n1325), .Y(n1810) );
  OAI21X1 U1742 ( .A(n1323), .B(n1359), .C(n1810), .Y(n2034) );
  NAND2X1 U1743 ( .A(\mem<6><4> ), .B(n1325), .Y(n1811) );
  OAI21X1 U1744 ( .A(n1323), .B(n1362), .C(n1811), .Y(n2033) );
  NAND2X1 U1745 ( .A(\mem<6><5> ), .B(n1325), .Y(n1812) );
  OAI21X1 U1746 ( .A(n1323), .B(n1365), .C(n1812), .Y(n2032) );
  NAND2X1 U1747 ( .A(\mem<6><6> ), .B(n1325), .Y(n1813) );
  OAI21X1 U1748 ( .A(n1323), .B(n1366), .C(n1813), .Y(n2031) );
  NAND2X1 U1749 ( .A(\mem<6><7> ), .B(n1325), .Y(n1814) );
  OAI21X1 U1750 ( .A(n1323), .B(n1367), .C(n1814), .Y(n2030) );
  NAND2X1 U1751 ( .A(\mem<6><8> ), .B(n1326), .Y(n1815) );
  OAI21X1 U1752 ( .A(n1324), .B(n1369), .C(n1815), .Y(n2029) );
  NAND2X1 U1753 ( .A(\mem<6><9> ), .B(n1326), .Y(n1816) );
  OAI21X1 U1754 ( .A(n1324), .B(n1371), .C(n1816), .Y(n2028) );
  NAND2X1 U1755 ( .A(\mem<6><10> ), .B(n1326), .Y(n1817) );
  OAI21X1 U1756 ( .A(n1324), .B(n1374), .C(n1817), .Y(n2027) );
  NAND2X1 U1757 ( .A(\mem<6><11> ), .B(n1326), .Y(n1818) );
  OAI21X1 U1758 ( .A(n1324), .B(n1377), .C(n1818), .Y(n2026) );
  NAND2X1 U1759 ( .A(\mem<6><12> ), .B(n1326), .Y(n1819) );
  OAI21X1 U1760 ( .A(n1324), .B(n1379), .C(n1819), .Y(n2025) );
  NAND2X1 U1761 ( .A(\mem<6><13> ), .B(n1326), .Y(n1820) );
  OAI21X1 U1762 ( .A(n1324), .B(n1380), .C(n1820), .Y(n2024) );
  NAND2X1 U1763 ( .A(\mem<6><14> ), .B(n1326), .Y(n1821) );
  OAI21X1 U1764 ( .A(n1324), .B(n1382), .C(n1821), .Y(n2023) );
  NAND2X1 U1765 ( .A(\mem<6><15> ), .B(n1326), .Y(n1822) );
  OAI21X1 U1766 ( .A(n1324), .B(n1384), .C(n1822), .Y(n2022) );
  NAND2X1 U1767 ( .A(\mem<5><0> ), .B(n1329), .Y(n1824) );
  OAI21X1 U1768 ( .A(n1327), .B(n1355), .C(n1824), .Y(n2021) );
  NAND2X1 U1769 ( .A(\mem<5><1> ), .B(n1329), .Y(n1825) );
  OAI21X1 U1770 ( .A(n1327), .B(n1356), .C(n1825), .Y(n2020) );
  NAND2X1 U1771 ( .A(\mem<5><2> ), .B(n1329), .Y(n1826) );
  OAI21X1 U1772 ( .A(n1327), .B(n1358), .C(n1826), .Y(n2019) );
  NAND2X1 U1773 ( .A(\mem<5><3> ), .B(n1329), .Y(n1827) );
  OAI21X1 U1774 ( .A(n1327), .B(n1359), .C(n1827), .Y(n2018) );
  NAND2X1 U1775 ( .A(\mem<5><4> ), .B(n1329), .Y(n1828) );
  OAI21X1 U1776 ( .A(n1327), .B(n1361), .C(n1828), .Y(n2017) );
  NAND2X1 U1777 ( .A(\mem<5><5> ), .B(n1329), .Y(n1829) );
  OAI21X1 U1778 ( .A(n1327), .B(n1364), .C(n1829), .Y(n2016) );
  NAND2X1 U1779 ( .A(\mem<5><6> ), .B(n1329), .Y(n1830) );
  OAI21X1 U1780 ( .A(n1327), .B(n1366), .C(n1830), .Y(n2015) );
  NAND2X1 U1781 ( .A(\mem<5><7> ), .B(n1329), .Y(n1831) );
  OAI21X1 U1782 ( .A(n1327), .B(n1367), .C(n1831), .Y(n2014) );
  NAND2X1 U1783 ( .A(\mem<5><8> ), .B(n1330), .Y(n1832) );
  OAI21X1 U1784 ( .A(n1328), .B(n1369), .C(n1832), .Y(n2013) );
  NAND2X1 U1785 ( .A(\mem<5><9> ), .B(n1330), .Y(n1833) );
  OAI21X1 U1786 ( .A(n1328), .B(n1371), .C(n1833), .Y(n2012) );
  NAND2X1 U1787 ( .A(\mem<5><10> ), .B(n1330), .Y(n1834) );
  OAI21X1 U1788 ( .A(n1328), .B(n1374), .C(n1834), .Y(n2011) );
  NAND2X1 U1789 ( .A(\mem<5><11> ), .B(n1330), .Y(n1835) );
  OAI21X1 U1790 ( .A(n1328), .B(n1376), .C(n1835), .Y(n2010) );
  NAND2X1 U1791 ( .A(\mem<5><12> ), .B(n1330), .Y(n1836) );
  OAI21X1 U1792 ( .A(n1328), .B(n1378), .C(n1836), .Y(n2009) );
  NAND2X1 U1793 ( .A(\mem<5><13> ), .B(n1330), .Y(n1837) );
  OAI21X1 U1794 ( .A(n1328), .B(n1380), .C(n1837), .Y(n2008) );
  NAND2X1 U1795 ( .A(\mem<5><14> ), .B(n1330), .Y(n1838) );
  OAI21X1 U1796 ( .A(n1328), .B(n1382), .C(n1838), .Y(n2007) );
  NAND2X1 U1797 ( .A(\mem<5><15> ), .B(n1330), .Y(n1839) );
  OAI21X1 U1798 ( .A(n1328), .B(n1384), .C(n1839), .Y(n2006) );
  NAND2X1 U1799 ( .A(\mem<4><0> ), .B(n1333), .Y(n1841) );
  OAI21X1 U1800 ( .A(n1331), .B(n1355), .C(n1841), .Y(n2005) );
  NAND2X1 U1801 ( .A(\mem<4><1> ), .B(n1333), .Y(n1842) );
  OAI21X1 U1802 ( .A(n1331), .B(n1356), .C(n1842), .Y(n2004) );
  NAND2X1 U1803 ( .A(\mem<4><2> ), .B(n1333), .Y(n1843) );
  OAI21X1 U1804 ( .A(n1331), .B(n1358), .C(n1843), .Y(n2003) );
  NAND2X1 U1805 ( .A(\mem<4><3> ), .B(n1333), .Y(n1844) );
  OAI21X1 U1806 ( .A(n1331), .B(n1359), .C(n1844), .Y(n2002) );
  NAND2X1 U1807 ( .A(\mem<4><4> ), .B(n1333), .Y(n1845) );
  OAI21X1 U1808 ( .A(n1331), .B(n1362), .C(n1845), .Y(n2001) );
  NAND2X1 U1809 ( .A(\mem<4><5> ), .B(n1333), .Y(n1846) );
  OAI21X1 U1810 ( .A(n1331), .B(n1365), .C(n1846), .Y(n2000) );
  NAND2X1 U1811 ( .A(\mem<4><6> ), .B(n1333), .Y(n1847) );
  OAI21X1 U1812 ( .A(n1331), .B(n1366), .C(n1847), .Y(n1999) );
  NAND2X1 U1813 ( .A(\mem<4><7> ), .B(n1333), .Y(n1848) );
  OAI21X1 U1814 ( .A(n1331), .B(n1367), .C(n1848), .Y(n1998) );
  NAND2X1 U1815 ( .A(\mem<4><8> ), .B(n1334), .Y(n1849) );
  OAI21X1 U1816 ( .A(n1332), .B(n1369), .C(n1849), .Y(n1997) );
  NAND2X1 U1817 ( .A(\mem<4><9> ), .B(n1334), .Y(n1850) );
  OAI21X1 U1818 ( .A(n1332), .B(n1371), .C(n1850), .Y(n1996) );
  NAND2X1 U1819 ( .A(\mem<4><10> ), .B(n1334), .Y(n1851) );
  OAI21X1 U1820 ( .A(n1332), .B(n1374), .C(n1851), .Y(n1995) );
  NAND2X1 U1821 ( .A(\mem<4><11> ), .B(n1334), .Y(n1852) );
  OAI21X1 U1822 ( .A(n1332), .B(n1376), .C(n1852), .Y(n1994) );
  NAND2X1 U1823 ( .A(\mem<4><12> ), .B(n1334), .Y(n1853) );
  OAI21X1 U1824 ( .A(n1332), .B(n1378), .C(n1853), .Y(n1993) );
  NAND2X1 U1825 ( .A(\mem<4><13> ), .B(n1334), .Y(n1854) );
  OAI21X1 U1826 ( .A(n1332), .B(n1380), .C(n1854), .Y(n1992) );
  NAND2X1 U1827 ( .A(\mem<4><14> ), .B(n1334), .Y(n1855) );
  OAI21X1 U1828 ( .A(n1332), .B(n1382), .C(n1855), .Y(n1991) );
  NAND2X1 U1829 ( .A(\mem<4><15> ), .B(n1334), .Y(n1856) );
  OAI21X1 U1830 ( .A(n1332), .B(n1384), .C(n1856), .Y(n1990) );
  NAND2X1 U1831 ( .A(\mem<3><0> ), .B(n1337), .Y(n1858) );
  OAI21X1 U1832 ( .A(n1335), .B(n1355), .C(n1858), .Y(n1989) );
  NAND2X1 U1833 ( .A(\mem<3><1> ), .B(n1337), .Y(n1859) );
  OAI21X1 U1834 ( .A(n1335), .B(n1356), .C(n1859), .Y(n1988) );
  NAND2X1 U1835 ( .A(\mem<3><2> ), .B(n1337), .Y(n1860) );
  OAI21X1 U1836 ( .A(n1335), .B(n1358), .C(n1860), .Y(n1987) );
  NAND2X1 U1837 ( .A(\mem<3><3> ), .B(n1337), .Y(n1861) );
  OAI21X1 U1838 ( .A(n1335), .B(n1359), .C(n1861), .Y(n1986) );
  NAND2X1 U1839 ( .A(\mem<3><4> ), .B(n1337), .Y(n1862) );
  OAI21X1 U1840 ( .A(n1335), .B(n1361), .C(n1862), .Y(n1985) );
  NAND2X1 U1841 ( .A(\mem<3><5> ), .B(n1337), .Y(n1863) );
  OAI21X1 U1842 ( .A(n1335), .B(n1364), .C(n1863), .Y(n1984) );
  NAND2X1 U1843 ( .A(\mem<3><6> ), .B(n1337), .Y(n1864) );
  OAI21X1 U1844 ( .A(n1335), .B(n1366), .C(n1864), .Y(n1983) );
  NAND2X1 U1845 ( .A(\mem<3><7> ), .B(n1337), .Y(n1865) );
  OAI21X1 U1846 ( .A(n1335), .B(n1367), .C(n1865), .Y(n1982) );
  NAND2X1 U1847 ( .A(\mem<3><8> ), .B(n1338), .Y(n1866) );
  OAI21X1 U1848 ( .A(n1336), .B(n1369), .C(n1866), .Y(n1981) );
  NAND2X1 U1849 ( .A(\mem<3><9> ), .B(n1338), .Y(n1867) );
  OAI21X1 U1850 ( .A(n1336), .B(n1371), .C(n1867), .Y(n1980) );
  NAND2X1 U1851 ( .A(\mem<3><10> ), .B(n1338), .Y(n1868) );
  OAI21X1 U1852 ( .A(n1336), .B(n1374), .C(n1868), .Y(n1979) );
  NAND2X1 U1853 ( .A(\mem<3><11> ), .B(n1338), .Y(n1869) );
  OAI21X1 U1854 ( .A(n1336), .B(n1377), .C(n1869), .Y(n1978) );
  NAND2X1 U1855 ( .A(\mem<3><12> ), .B(n1338), .Y(n1870) );
  OAI21X1 U1856 ( .A(n1336), .B(n1379), .C(n1870), .Y(n1977) );
  NAND2X1 U1857 ( .A(\mem<3><13> ), .B(n1338), .Y(n1871) );
  OAI21X1 U1858 ( .A(n1336), .B(n1380), .C(n1871), .Y(n1976) );
  NAND2X1 U1859 ( .A(\mem<3><14> ), .B(n1338), .Y(n1872) );
  OAI21X1 U1860 ( .A(n1336), .B(n1382), .C(n1872), .Y(n1975) );
  NAND2X1 U1861 ( .A(\mem<3><15> ), .B(n1338), .Y(n1873) );
  OAI21X1 U1862 ( .A(n1336), .B(n1384), .C(n1873), .Y(n1974) );
  NAND2X1 U1863 ( .A(\mem<2><0> ), .B(n1341), .Y(n1875) );
  OAI21X1 U1864 ( .A(n1339), .B(n1355), .C(n1875), .Y(n1973) );
  NAND2X1 U1865 ( .A(\mem<2><1> ), .B(n1341), .Y(n1876) );
  OAI21X1 U1866 ( .A(n1339), .B(n1356), .C(n1876), .Y(n1972) );
  NAND2X1 U1867 ( .A(\mem<2><2> ), .B(n1341), .Y(n1877) );
  OAI21X1 U1868 ( .A(n1339), .B(n1358), .C(n1877), .Y(n1971) );
  NAND2X1 U1869 ( .A(\mem<2><3> ), .B(n1341), .Y(n1878) );
  OAI21X1 U1870 ( .A(n1339), .B(n1359), .C(n1878), .Y(n1970) );
  NAND2X1 U1871 ( .A(\mem<2><4> ), .B(n1341), .Y(n1879) );
  OAI21X1 U1872 ( .A(n1339), .B(n1362), .C(n1879), .Y(n1969) );
  NAND2X1 U1873 ( .A(\mem<2><5> ), .B(n1341), .Y(n1880) );
  OAI21X1 U1874 ( .A(n1339), .B(n1365), .C(n1880), .Y(n1968) );
  NAND2X1 U1875 ( .A(\mem<2><6> ), .B(n1341), .Y(n1881) );
  OAI21X1 U1876 ( .A(n1339), .B(n1366), .C(n1881), .Y(n1967) );
  NAND2X1 U1877 ( .A(\mem<2><7> ), .B(n1341), .Y(n1882) );
  OAI21X1 U1878 ( .A(n1339), .B(n1367), .C(n1882), .Y(n1966) );
  NAND2X1 U1879 ( .A(\mem<2><8> ), .B(n1342), .Y(n1883) );
  OAI21X1 U1880 ( .A(n1340), .B(n1369), .C(n1883), .Y(n1965) );
  NAND2X1 U1881 ( .A(\mem<2><9> ), .B(n1342), .Y(n1884) );
  OAI21X1 U1882 ( .A(n1340), .B(n1371), .C(n1884), .Y(n1964) );
  NAND2X1 U1883 ( .A(\mem<2><10> ), .B(n1342), .Y(n1885) );
  OAI21X1 U1884 ( .A(n1340), .B(n1374), .C(n1885), .Y(n1963) );
  NAND2X1 U1885 ( .A(\mem<2><11> ), .B(n1342), .Y(n1886) );
  OAI21X1 U1886 ( .A(n1340), .B(n1376), .C(n1886), .Y(n1962) );
  NAND2X1 U1887 ( .A(\mem<2><12> ), .B(n1342), .Y(n1887) );
  OAI21X1 U1888 ( .A(n1340), .B(n1378), .C(n1887), .Y(n1961) );
  NAND2X1 U1889 ( .A(\mem<2><13> ), .B(n1342), .Y(n1888) );
  OAI21X1 U1890 ( .A(n1340), .B(n1380), .C(n1888), .Y(n1960) );
  NAND2X1 U1891 ( .A(\mem<2><14> ), .B(n1342), .Y(n1889) );
  OAI21X1 U1892 ( .A(n1340), .B(n1382), .C(n1889), .Y(n1959) );
  NAND2X1 U1893 ( .A(\mem<2><15> ), .B(n1342), .Y(n1890) );
  OAI21X1 U1894 ( .A(n1340), .B(n1384), .C(n1890), .Y(n1958) );
  NAND2X1 U1895 ( .A(\mem<1><0> ), .B(n1345), .Y(n1892) );
  OAI21X1 U1896 ( .A(n1343), .B(n1355), .C(n1892), .Y(n1957) );
  NAND2X1 U1897 ( .A(\mem<1><1> ), .B(n1345), .Y(n1893) );
  OAI21X1 U1898 ( .A(n1343), .B(n1356), .C(n1893), .Y(n1956) );
  NAND2X1 U1899 ( .A(\mem<1><2> ), .B(n1345), .Y(n1894) );
  OAI21X1 U1900 ( .A(n1343), .B(n1358), .C(n1894), .Y(n1955) );
  NAND2X1 U1901 ( .A(\mem<1><3> ), .B(n1345), .Y(n1895) );
  OAI21X1 U1902 ( .A(n1343), .B(n1359), .C(n1895), .Y(n1954) );
  NAND2X1 U1903 ( .A(\mem<1><4> ), .B(n1345), .Y(n1896) );
  OAI21X1 U1904 ( .A(n1343), .B(n1361), .C(n1896), .Y(n1953) );
  NAND2X1 U1905 ( .A(\mem<1><5> ), .B(n1345), .Y(n1897) );
  OAI21X1 U1906 ( .A(n1343), .B(n1364), .C(n1897), .Y(n1952) );
  NAND2X1 U1907 ( .A(\mem<1><6> ), .B(n1345), .Y(n1898) );
  OAI21X1 U1908 ( .A(n1343), .B(n1366), .C(n1898), .Y(n1951) );
  NAND2X1 U1909 ( .A(\mem<1><7> ), .B(n1345), .Y(n1899) );
  OAI21X1 U1910 ( .A(n1343), .B(n1367), .C(n1899), .Y(n1950) );
  NAND2X1 U1911 ( .A(\mem<1><8> ), .B(n1346), .Y(n1900) );
  OAI21X1 U1912 ( .A(n1344), .B(n1369), .C(n1900), .Y(n1949) );
  NAND2X1 U1913 ( .A(\mem<1><9> ), .B(n1346), .Y(n1901) );
  OAI21X1 U1914 ( .A(n1344), .B(n1371), .C(n1901), .Y(n1948) );
  NAND2X1 U1915 ( .A(\mem<1><10> ), .B(n1346), .Y(n1902) );
  OAI21X1 U1916 ( .A(n1344), .B(n1374), .C(n1902), .Y(n1947) );
  NAND2X1 U1917 ( .A(\mem<1><11> ), .B(n1346), .Y(n1903) );
  OAI21X1 U1918 ( .A(n1344), .B(n1377), .C(n1903), .Y(n1946) );
  NAND2X1 U1919 ( .A(\mem<1><12> ), .B(n1346), .Y(n1904) );
  OAI21X1 U1920 ( .A(n1344), .B(n1379), .C(n1904), .Y(n1945) );
  NAND2X1 U1921 ( .A(\mem<1><13> ), .B(n1346), .Y(n1905) );
  OAI21X1 U1922 ( .A(n1344), .B(n1380), .C(n1905), .Y(n1944) );
  NAND2X1 U1923 ( .A(\mem<1><14> ), .B(n1346), .Y(n1906) );
  OAI21X1 U1924 ( .A(n1344), .B(n1382), .C(n1906), .Y(n1943) );
  NAND2X1 U1925 ( .A(\mem<1><15> ), .B(n1346), .Y(n1907) );
  OAI21X1 U1926 ( .A(n1344), .B(n1384), .C(n1907), .Y(n1942) );
  NAND2X1 U1927 ( .A(\mem<0><0> ), .B(n1348), .Y(n1910) );
  OAI21X1 U1928 ( .A(n1347), .B(n1355), .C(n1910), .Y(n1941) );
  NAND2X1 U1929 ( .A(\mem<0><1> ), .B(n1348), .Y(n1911) );
  OAI21X1 U1930 ( .A(n1347), .B(n1356), .C(n1911), .Y(n1940) );
  NAND2X1 U1931 ( .A(\mem<0><2> ), .B(n1348), .Y(n1912) );
  OAI21X1 U1932 ( .A(n1347), .B(n1358), .C(n1912), .Y(n1939) );
  NAND2X1 U1933 ( .A(\mem<0><3> ), .B(n1348), .Y(n1913) );
  OAI21X1 U1934 ( .A(n1347), .B(n1359), .C(n1913), .Y(n1938) );
  NAND2X1 U1935 ( .A(\mem<0><4> ), .B(n1348), .Y(n1914) );
  OAI21X1 U1936 ( .A(n1347), .B(n1361), .C(n1914), .Y(n1937) );
  NAND2X1 U1937 ( .A(\mem<0><5> ), .B(n1348), .Y(n1915) );
  OAI21X1 U1938 ( .A(n1347), .B(n1365), .C(n1915), .Y(n1936) );
  NAND2X1 U1939 ( .A(\mem<0><6> ), .B(n1348), .Y(n1916) );
  OAI21X1 U1940 ( .A(n1347), .B(n1366), .C(n1916), .Y(n1935) );
  NAND2X1 U1941 ( .A(\mem<0><7> ), .B(n1348), .Y(n1917) );
  OAI21X1 U1942 ( .A(n1347), .B(n1367), .C(n1917), .Y(n1934) );
  NAND2X1 U1943 ( .A(\mem<0><8> ), .B(n1349), .Y(n1918) );
  OAI21X1 U1944 ( .A(n1347), .B(n1369), .C(n1918), .Y(n1933) );
  NAND2X1 U1945 ( .A(\mem<0><9> ), .B(n1349), .Y(n1919) );
  OAI21X1 U1946 ( .A(n1347), .B(n1371), .C(n1919), .Y(n1932) );
  NAND2X1 U1947 ( .A(\mem<0><10> ), .B(n1349), .Y(n1920) );
  OAI21X1 U1948 ( .A(n1347), .B(n1374), .C(n1920), .Y(n1931) );
  NAND2X1 U1949 ( .A(\mem<0><11> ), .B(n1349), .Y(n1921) );
  OAI21X1 U1950 ( .A(n1347), .B(n1376), .C(n1921), .Y(n1930) );
  NAND2X1 U1951 ( .A(\mem<0><12> ), .B(n1349), .Y(n1922) );
  OAI21X1 U1952 ( .A(n1347), .B(n1378), .C(n1922), .Y(n1929) );
  NAND2X1 U1953 ( .A(\mem<0><13> ), .B(n1349), .Y(n1923) );
  OAI21X1 U1954 ( .A(n1347), .B(n1380), .C(n1923), .Y(n1928) );
  NAND2X1 U1955 ( .A(\mem<0><14> ), .B(n1349), .Y(n1924) );
  OAI21X1 U1956 ( .A(n1347), .B(n1382), .C(n1924), .Y(n1927) );
  NAND2X1 U1957 ( .A(\mem<0><15> ), .B(n1349), .Y(n1925) );
  OAI21X1 U1958 ( .A(n1347), .B(n1384), .C(n1925), .Y(n1926) );
endmodule


module memc_Size16_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1896), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1897), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1898), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1899), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1900), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1901), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1902), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1903), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1904), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1905), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1906), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1907), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1908), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1909), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1910), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1911), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1912), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1913), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1914), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1915), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1916), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1917), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1918), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1919), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1920), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1921), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1922), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1923), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1924), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1925), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1926), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1927), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1928), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1929), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1930), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1931), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1932), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1933), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1934), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1935), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1936), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1937), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1938), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1939), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1940), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1941), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1942), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1943), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1944), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1945), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1946), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1947), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1948), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1949), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1950), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1951), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1952), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1953), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1954), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1955), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1956), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1957), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1958), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1959), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1960), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1961), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1962), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1963), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1964), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1965), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1966), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1967), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1968), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1969), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1970), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1971), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1972), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1973), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1974), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1975), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1976), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1977), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1978), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1979), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1980), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1981), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1982), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1983), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1984), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1985), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1986), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1987), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1988), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1989), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1990), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1991), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1992), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1993), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1994), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1995), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1996), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1997), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1998), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1999), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2000), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2001), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2002), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2003), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2004), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2005), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2006), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2007), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2008), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2009), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2010), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2011), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2012), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2013), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2014), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2015), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2016), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2017), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2018), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2019), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2020), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2021), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2022), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2023), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2024), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2025), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2026), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2027), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2028), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2029), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2030), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2031), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2032), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2033), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2034), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2035), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2036), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2037), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2038), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2039), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2040), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2041), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2042), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2043), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2044), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2045), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2046), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2047), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2048), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2049), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2050), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2051), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2052), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2053), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2054), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2055), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2056), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2057), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2058), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2059), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2060), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2061), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2062), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2063), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2064), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2065), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2066), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2067), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2068), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2069), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2070), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2071), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2072), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2073), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2074), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2075), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2076), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2077), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2078), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2079), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2080), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2081), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2082), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2083), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2084), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2085), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2086), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2087), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2088), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2089), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2090), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2091), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2092), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2093), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2094), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2095), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2096), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2097), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2098), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2099), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2100), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2101), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2102), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2103), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2104), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2105), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2106), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2107), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2108), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2109), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2110), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2111), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2112), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2113), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2114), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2115), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2116), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2117), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2118), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2119), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2120), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2121), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2122), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2123), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2124), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2125), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2126), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2127), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2128), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2129), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2130), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2131), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2132), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2133), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2134), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2135), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2136), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2137), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2138), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2139), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2140), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2141), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2142), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2143), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2144), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2145), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2146), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2147), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2148), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2149), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2150), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2151), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2152), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2153), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2154), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2155), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2156), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2157), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2158), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2159), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2160), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2161), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2162), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2163), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2164), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2165), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2166), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2167), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2168), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2169), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2170), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2171), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2172), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2173), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2174), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2175), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2176), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2177), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2178), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2179), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2180), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2181), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2182), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2183), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2184), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2185), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2186), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2187), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2188), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2189), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2190), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2191), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2192), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2193), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2194), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2195), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2196), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2197), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2198), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2199), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2200), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2201), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2202), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2203), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2204), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2205), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2206), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2207), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2208), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2209), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2210), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2211), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2212), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2213), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2214), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2215), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2216), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2217), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2218), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2219), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2220), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2221), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2222), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2223), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2224), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2225), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2226), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2227), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2228), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2229), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2230), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2231), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2232), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2233), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2234), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2235), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2236), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2237), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2238), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2239), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2240), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2241), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2242), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2243), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2244), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2245), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2246), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2247), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2248), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2249), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2250), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2251), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2252), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2253), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2254), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2255), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2256), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2257), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2258), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2259), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2260), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2261), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2262), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2263), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2264), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2265), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2266), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2267), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2268), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2269), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2270), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2271), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2272), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2273), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2274), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2275), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2276), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2277), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2278), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2279), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2280), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2281), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2282), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2283), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2284), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2285), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2286), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2287), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2288), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2289), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2290), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2291), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2292), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2293), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2294), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2295), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2296), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2297), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2298), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2299), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2300), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2301), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2302), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2303), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2304), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2305), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2306), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2307), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2308), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2309), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2310), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2311), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2312), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2313), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2314), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2315), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2316), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2317), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2318), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2319), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2320), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2321), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2322), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2323), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2324), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2325), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2326), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2327), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2328), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2329), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2330), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2331), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2332), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2333), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2334), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2335), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2336), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2337), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2338), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2339), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2340), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2341), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2342), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2343), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2344), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2345), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2346), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2347), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2348), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2349), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2350), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2351), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2352), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2353), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2354), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2355), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2356), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2357), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2358), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2359), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2360), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2361), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2362), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2363), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2364), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2365), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2366), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2367), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2368), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2369), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2370), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2371), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2372), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2373), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2374), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2375), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2376), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2377), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2378), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2379), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2380), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2381), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2382), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2383), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2384), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2385), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2386), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2387), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2388), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2389), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2390), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2391), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2392), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2393), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2394), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2395), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2396), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2397), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2398), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2399), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2400), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2401), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2402), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2403), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2404), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2405), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2406), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2407), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2408) );
  INVX1 U2 ( .A(n1355), .Y(n1191) );
  INVX1 U3 ( .A(n1355), .Y(n1190) );
  INVX1 U4 ( .A(n1232), .Y(n1209) );
  INVX1 U5 ( .A(n1232), .Y(n1208) );
  INVX1 U6 ( .A(n1211), .Y(n1212) );
  INVX1 U7 ( .A(n1194), .Y(n1195) );
  INVX1 U8 ( .A(n1211), .Y(n1213) );
  INVX1 U9 ( .A(n1194), .Y(n1196) );
  INVX2 U10 ( .A(n1210), .Y(n1215) );
  INVX2 U11 ( .A(n1210), .Y(n1216) );
  INVX1 U12 ( .A(n1194), .Y(n1197) );
  INVX1 U13 ( .A(n1206), .Y(n1198) );
  INVX1 U14 ( .A(n1206), .Y(n1199) );
  INVX1 U15 ( .A(n1209), .Y(n1221) );
  INVX1 U16 ( .A(n1209), .Y(n1222) );
  INVX1 U17 ( .A(n1206), .Y(n1200) );
  INVX1 U18 ( .A(n1208), .Y(n1223) );
  INVX1 U19 ( .A(n1208), .Y(n1224) );
  INVX1 U20 ( .A(n1193), .Y(n1201) );
  INVX1 U21 ( .A(n1207), .Y(n1226) );
  INVX1 U22 ( .A(n1193), .Y(n1202) );
  INVX2 U23 ( .A(n1207), .Y(n1227) );
  INVX2 U24 ( .A(n1207), .Y(n1228) );
  INVX1 U25 ( .A(n1193), .Y(n1203) );
  INVX2 U26 ( .A(n1211), .Y(n1229) );
  INVX2 U27 ( .A(n1211), .Y(n1230) );
  INVX1 U28 ( .A(n1194), .Y(n1204) );
  INVX1 U29 ( .A(n1209), .Y(n1220) );
  INVX1 U30 ( .A(n1208), .Y(n1225) );
  INVX2 U31 ( .A(n1207), .Y(n1231) );
  INVX1 U32 ( .A(n1193), .Y(n1205) );
  INVX1 U33 ( .A(n1170), .Y(N32) );
  INVX1 U34 ( .A(n1171), .Y(N31) );
  INVX1 U35 ( .A(n1172), .Y(N30) );
  INVX1 U36 ( .A(n1173), .Y(N29) );
  INVX1 U37 ( .A(n1174), .Y(N28) );
  INVX1 U38 ( .A(n1175), .Y(N27) );
  INVX1 U39 ( .A(n1176), .Y(N26) );
  INVX1 U40 ( .A(n1177), .Y(N25) );
  INVX1 U41 ( .A(n1178), .Y(N24) );
  INVX1 U42 ( .A(n1179), .Y(N23) );
  INVX1 U43 ( .A(n1180), .Y(N22) );
  INVX1 U44 ( .A(n1181), .Y(N21) );
  INVX1 U45 ( .A(n1182), .Y(N20) );
  INVX1 U46 ( .A(n1183), .Y(N19) );
  INVX1 U47 ( .A(n1184), .Y(N18) );
  INVX1 U48 ( .A(n1185), .Y(N17) );
  BUFX2 U49 ( .A(n105), .Y(n1233) );
  BUFX2 U50 ( .A(n107), .Y(n1235) );
  BUFX2 U51 ( .A(n109), .Y(n1237) );
  BUFX2 U52 ( .A(n111), .Y(n1239) );
  BUFX2 U53 ( .A(n113), .Y(n1241) );
  BUFX2 U54 ( .A(n115), .Y(n1243) );
  BUFX2 U55 ( .A(n117), .Y(n1245) );
  BUFX2 U56 ( .A(n119), .Y(n1247) );
  BUFX2 U57 ( .A(n121), .Y(n1249) );
  BUFX2 U58 ( .A(n123), .Y(n1253) );
  BUFX2 U59 ( .A(n125), .Y(n1257) );
  BUFX2 U60 ( .A(n127), .Y(n1261) );
  BUFX2 U61 ( .A(n130), .Y(n1263) );
  BUFX2 U62 ( .A(n133), .Y(n1265) );
  BUFX2 U63 ( .A(n137), .Y(n1268) );
  BUFX2 U64 ( .A(n140), .Y(n1270) );
  BUFX2 U65 ( .A(n142), .Y(n1274) );
  BUFX2 U66 ( .A(n144), .Y(n1278) );
  BUFX2 U67 ( .A(n146), .Y(n1282) );
  BUFX2 U68 ( .A(n148), .Y(n1286) );
  BUFX2 U69 ( .A(n150), .Y(n1290) );
  BUFX2 U70 ( .A(n152), .Y(n1297) );
  BUFX2 U71 ( .A(n154), .Y(n1301) );
  BUFX2 U72 ( .A(n156), .Y(n1305) );
  BUFX2 U73 ( .A(n158), .Y(n1309) );
  BUFX2 U74 ( .A(n160), .Y(n1311) );
  BUFX2 U75 ( .A(n162), .Y(n1313) );
  BUFX2 U76 ( .A(n165), .Y(n1315) );
  INVX1 U77 ( .A(n1232), .Y(n1207) );
  INVX1 U78 ( .A(n1355), .Y(n1192) );
  INVX1 U79 ( .A(n1357), .Y(n1187) );
  INVX1 U80 ( .A(n1359), .Y(n1358) );
  INVX1 U81 ( .A(N14), .Y(n1359) );
  INVX1 U82 ( .A(n1353), .Y(n1206) );
  INVX1 U83 ( .A(n1351), .Y(n1210) );
  INVX1 U84 ( .A(n1355), .Y(n1189) );
  INVX1 U85 ( .A(n1355), .Y(n1188) );
  INVX1 U86 ( .A(n1359), .Y(n1186) );
  INVX1 U87 ( .A(n1357), .Y(n1356) );
  INVX1 U88 ( .A(N13), .Y(n1357) );
  BUFX2 U89 ( .A(n115), .Y(n1244) );
  BUFX2 U90 ( .A(n113), .Y(n1242) );
  BUFX2 U91 ( .A(n109), .Y(n1238) );
  INVX1 U92 ( .A(n1353), .Y(n1194) );
  INVX1 U93 ( .A(n1353), .Y(n1193) );
  INVX1 U94 ( .A(n102), .Y(n1294) );
  INVX1 U95 ( .A(n103), .Y(n1317) );
  BUFX2 U96 ( .A(n123), .Y(n1254) );
  BUFX2 U97 ( .A(n125), .Y(n1258) );
  BUFX2 U98 ( .A(n142), .Y(n1275) );
  BUFX2 U99 ( .A(n146), .Y(n1283) );
  BUFX2 U100 ( .A(n148), .Y(n1287) );
  BUFX2 U101 ( .A(n150), .Y(n1291) );
  BUFX2 U102 ( .A(n156), .Y(n1306) );
  INVX1 U103 ( .A(n1352), .Y(n1232) );
  INVX1 U104 ( .A(rst), .Y(n1350) );
  BUFX2 U105 ( .A(n105), .Y(n1234) );
  BUFX2 U106 ( .A(n121), .Y(n1250) );
  BUFX2 U107 ( .A(n127), .Y(n1262) );
  BUFX2 U108 ( .A(n130), .Y(n1264) );
  BUFX2 U109 ( .A(n133), .Y(n1266) );
  BUFX2 U110 ( .A(n137), .Y(n1269) );
  BUFX2 U111 ( .A(n140), .Y(n1271) );
  BUFX2 U112 ( .A(n144), .Y(n1279) );
  BUFX2 U113 ( .A(n152), .Y(n1298) );
  BUFX2 U114 ( .A(n154), .Y(n1302) );
  BUFX2 U115 ( .A(n158), .Y(n1310) );
  BUFX2 U116 ( .A(n160), .Y(n1312) );
  BUFX2 U117 ( .A(n162), .Y(n1314) );
  BUFX2 U118 ( .A(n165), .Y(n1316) );
  BUFX2 U119 ( .A(n119), .Y(n1248) );
  BUFX2 U120 ( .A(n117), .Y(n1246) );
  BUFX2 U121 ( .A(n111), .Y(n1240) );
  BUFX2 U122 ( .A(n107), .Y(n1236) );
  INVX1 U123 ( .A(n101), .Y(n1267) );
  INVX1 U124 ( .A(n1232), .Y(n1211) );
  INVX4 U125 ( .A(n64), .Y(n65) );
  INVX4 U126 ( .A(n62), .Y(n63) );
  INVX4 U127 ( .A(n68), .Y(n167) );
  INVX4 U128 ( .A(n40), .Y(n135) );
  INVX4 U129 ( .A(n67), .Y(n166) );
  INVX4 U130 ( .A(n66), .Y(n163) );
  INVX4 U131 ( .A(n41), .Y(n138) );
  INVX4 U132 ( .A(n39), .Y(n134) );
  INVX4 U133 ( .A(n38), .Y(n131) );
  INVX4 U134 ( .A(n37), .Y(n128) );
  INVX1 U135 ( .A(n69), .Y(n1) );
  INVX1 U136 ( .A(n69), .Y(n2) );
  INVX1 U137 ( .A(n69), .Y(n3) );
  INVX1 U138 ( .A(n69), .Y(n4) );
  INVX1 U139 ( .A(n69), .Y(n5) );
  INVX1 U140 ( .A(n4), .Y(n6) );
  INVX1 U141 ( .A(n1), .Y(n7) );
  INVX1 U142 ( .A(n2), .Y(n8) );
  INVX1 U143 ( .A(n1), .Y(n9) );
  INVX1 U144 ( .A(n1), .Y(n10) );
  INVX1 U145 ( .A(n3), .Y(n11) );
  INVX1 U146 ( .A(n2), .Y(n12) );
  INVX1 U147 ( .A(n2), .Y(n13) );
  INVX1 U148 ( .A(n2), .Y(n14) );
  INVX1 U149 ( .A(n3), .Y(n15) );
  INVX1 U150 ( .A(n3), .Y(n16) );
  INVX1 U151 ( .A(n3), .Y(n17) );
  INVX1 U152 ( .A(n4), .Y(n18) );
  INVX1 U153 ( .A(n4), .Y(n19) );
  INVX1 U154 ( .A(n4), .Y(n20) );
  INVX1 U155 ( .A(n5), .Y(n21) );
  INVX1 U156 ( .A(n5), .Y(n22) );
  INVX1 U157 ( .A(n5), .Y(n23) );
  BUFX2 U158 ( .A(n1), .Y(n24) );
  INVX1 U159 ( .A(n24), .Y(n25) );
  INVX1 U160 ( .A(n24), .Y(n26) );
  INVX1 U161 ( .A(n29), .Y(n27) );
  INVX2 U162 ( .A(n29), .Y(n28) );
  INVX2 U163 ( .A(n29), .Y(n30) );
  OR2X2 U164 ( .A(write), .B(rst), .Y(n29) );
  AND2X2 U165 ( .A(n18), .B(n120), .Y(n31) );
  INVX1 U166 ( .A(n31), .Y(n32) );
  AND2X2 U167 ( .A(n19), .B(n122), .Y(n33) );
  INVX1 U168 ( .A(n33), .Y(n34) );
  AND2X2 U169 ( .A(n20), .B(n124), .Y(n35) );
  INVX1 U170 ( .A(n35), .Y(n36) );
  AND2X2 U171 ( .A(n25), .B(n126), .Y(n37) );
  AND2X2 U172 ( .A(n26), .B(n129), .Y(n38) );
  AND2X2 U173 ( .A(n16), .B(n132), .Y(n39) );
  AND2X2 U174 ( .A(n17), .B(n101), .Y(n40) );
  AND2X2 U175 ( .A(n16), .B(n136), .Y(n41) );
  AND2X2 U176 ( .A(n6), .B(n139), .Y(n42) );
  INVX1 U177 ( .A(n42), .Y(n43) );
  AND2X2 U178 ( .A(n6), .B(n141), .Y(n44) );
  INVX1 U179 ( .A(n44), .Y(n45) );
  AND2X2 U180 ( .A(n7), .B(n143), .Y(n46) );
  INVX1 U181 ( .A(n46), .Y(n47) );
  AND2X2 U182 ( .A(n8), .B(n145), .Y(n48) );
  INVX1 U183 ( .A(n48), .Y(n49) );
  AND2X2 U184 ( .A(n9), .B(n147), .Y(n50) );
  INVX1 U185 ( .A(n50), .Y(n51) );
  AND2X2 U186 ( .A(n10), .B(n149), .Y(n52) );
  INVX1 U187 ( .A(n52), .Y(n53) );
  AND2X2 U188 ( .A(n7), .B(n102), .Y(n54) );
  INVX1 U189 ( .A(n54), .Y(n55) );
  AND2X2 U190 ( .A(n21), .B(n151), .Y(n56) );
  INVX1 U191 ( .A(n56), .Y(n57) );
  AND2X2 U192 ( .A(n22), .B(n153), .Y(n58) );
  INVX1 U193 ( .A(n58), .Y(n59) );
  AND2X2 U194 ( .A(n23), .B(n155), .Y(n60) );
  INVX1 U195 ( .A(n60), .Y(n61) );
  AND2X2 U196 ( .A(n14), .B(n157), .Y(n62) );
  AND2X2 U197 ( .A(n13), .B(n159), .Y(n64) );
  AND2X2 U198 ( .A(n17), .B(n161), .Y(n66) );
  AND2X2 U199 ( .A(n12), .B(n164), .Y(n67) );
  AND2X2 U200 ( .A(n11), .B(n103), .Y(n68) );
  BUFX2 U201 ( .A(n43), .Y(n1272) );
  BUFX2 U202 ( .A(n43), .Y(n1273) );
  BUFX2 U203 ( .A(n45), .Y(n1276) );
  BUFX2 U204 ( .A(n45), .Y(n1277) );
  BUFX2 U205 ( .A(n47), .Y(n1280) );
  BUFX2 U206 ( .A(n47), .Y(n1281) );
  BUFX2 U207 ( .A(n49), .Y(n1284) );
  BUFX2 U208 ( .A(n49), .Y(n1285) );
  BUFX2 U209 ( .A(n51), .Y(n1288) );
  BUFX2 U210 ( .A(n51), .Y(n1289) );
  BUFX2 U211 ( .A(n53), .Y(n1292) );
  BUFX2 U212 ( .A(n53), .Y(n1293) );
  BUFX2 U213 ( .A(n55), .Y(n1295) );
  BUFX2 U214 ( .A(n55), .Y(n1296) );
  BUFX2 U215 ( .A(n57), .Y(n1299) );
  BUFX2 U216 ( .A(n57), .Y(n1300) );
  BUFX2 U217 ( .A(n59), .Y(n1303) );
  BUFX2 U218 ( .A(n59), .Y(n1304) );
  BUFX2 U219 ( .A(n61), .Y(n1307) );
  BUFX2 U220 ( .A(n61), .Y(n1308) );
  AND2X2 U221 ( .A(write), .B(n1350), .Y(n69) );
  AND2X2 U222 ( .A(\data_in<0> ), .B(n20), .Y(n70) );
  AND2X2 U223 ( .A(\data_in<1> ), .B(n17), .Y(n71) );
  AND2X2 U224 ( .A(\data_in<2> ), .B(n23), .Y(n72) );
  AND2X2 U225 ( .A(\data_in<3> ), .B(n17), .Y(n73) );
  AND2X2 U226 ( .A(\data_in<4> ), .B(n15), .Y(n74) );
  AND2X2 U227 ( .A(\data_in<5> ), .B(n18), .Y(n75) );
  AND2X2 U228 ( .A(\data_in<6> ), .B(n16), .Y(n76) );
  AND2X2 U229 ( .A(\data_in<7> ), .B(n19), .Y(n77) );
  AND2X2 U230 ( .A(\data_in<8> ), .B(n21), .Y(n78) );
  AND2X2 U231 ( .A(\data_in<9> ), .B(n22), .Y(n79) );
  AND2X2 U232 ( .A(\data_in<10> ), .B(n16), .Y(n80) );
  AND2X2 U233 ( .A(\data_in<11> ), .B(n13), .Y(n81) );
  AND2X2 U234 ( .A(\data_in<12> ), .B(n12), .Y(n82) );
  AND2X2 U235 ( .A(\data_in<13> ), .B(n14), .Y(n83) );
  AND2X2 U236 ( .A(\data_in<14> ), .B(n15), .Y(n84) );
  AND2X2 U237 ( .A(\data_in<15> ), .B(n16), .Y(n85) );
  INVX1 U238 ( .A(n1352), .Y(n1351) );
  INVX1 U239 ( .A(N12), .Y(n1355) );
  AND2X1 U240 ( .A(n1192), .B(n1353), .Y(n86) );
  INVX1 U241 ( .A(n1354), .Y(n1353) );
  AND2X1 U242 ( .A(n2408), .B(n1358), .Y(n87) );
  INVX2 U243 ( .A(n176), .Y(n1375) );
  INVX2 U244 ( .A(n175), .Y(n1392) );
  INVX2 U245 ( .A(n173), .Y(n1410) );
  INVX2 U246 ( .A(n174), .Y(n1428) );
  INVX2 U247 ( .A(n172), .Y(n1446) );
  INVX2 U248 ( .A(n171), .Y(n1464) );
  INVX2 U249 ( .A(n170), .Y(n1482) );
  INVX2 U250 ( .A(n168), .Y(n1499) );
  INVX2 U251 ( .A(n169), .Y(n1516) );
  BUFX2 U252 ( .A(n1394), .Y(n88) );
  INVX1 U253 ( .A(n88), .Y(n1793) );
  BUFX2 U254 ( .A(n1412), .Y(n89) );
  INVX1 U255 ( .A(n89), .Y(n1810) );
  BUFX2 U256 ( .A(n1430), .Y(n90) );
  INVX1 U257 ( .A(n90), .Y(n1827) );
  BUFX2 U258 ( .A(n1448), .Y(n91) );
  INVX1 U259 ( .A(n91), .Y(n1844) );
  BUFX2 U260 ( .A(n1466), .Y(n92) );
  INVX1 U261 ( .A(n92), .Y(n1861) );
  BUFX2 U262 ( .A(n1630), .Y(n93) );
  INVX1 U263 ( .A(n93), .Y(n1743) );
  BUFX2 U264 ( .A(n1760), .Y(n94) );
  INVX1 U265 ( .A(n94), .Y(n1878) );
  AND2X1 U266 ( .A(n1351), .B(n86), .Y(n95) );
  AND2X1 U267 ( .A(n1356), .B(n87), .Y(n96) );
  AND2X1 U268 ( .A(n1352), .B(n86), .Y(n97) );
  AND2X1 U269 ( .A(n1357), .B(n87), .Y(n98) );
  AND2X1 U270 ( .A(n96), .B(n1879), .Y(n99) );
  INVX1 U271 ( .A(n99), .Y(n100) );
  AND2X1 U272 ( .A(n1879), .B(n98), .Y(n101) );
  AND2X1 U273 ( .A(n1879), .B(n1743), .Y(n102) );
  AND2X1 U274 ( .A(n1879), .B(n1878), .Y(n103) );
  AND2X1 U275 ( .A(n95), .B(n96), .Y(n104) );
  INVX1 U276 ( .A(n104), .Y(n105) );
  AND2X1 U277 ( .A(n96), .B(n97), .Y(n106) );
  INVX1 U278 ( .A(n106), .Y(n107) );
  AND2X1 U279 ( .A(n96), .B(n1793), .Y(n108) );
  INVX1 U280 ( .A(n108), .Y(n109) );
  AND2X1 U281 ( .A(n96), .B(n1810), .Y(n110) );
  INVX1 U282 ( .A(n110), .Y(n111) );
  AND2X1 U283 ( .A(n96), .B(n1827), .Y(n112) );
  INVX1 U284 ( .A(n112), .Y(n113) );
  AND2X1 U285 ( .A(n96), .B(n1844), .Y(n114) );
  INVX1 U286 ( .A(n114), .Y(n115) );
  AND2X1 U287 ( .A(n96), .B(n1861), .Y(n116) );
  INVX1 U288 ( .A(n116), .Y(n117) );
  AND2X1 U289 ( .A(n95), .B(n98), .Y(n118) );
  INVX1 U290 ( .A(n118), .Y(n119) );
  AND2X1 U291 ( .A(n97), .B(n98), .Y(n120) );
  INVX1 U292 ( .A(n120), .Y(n121) );
  AND2X1 U293 ( .A(n1793), .B(n98), .Y(n122) );
  INVX1 U294 ( .A(n122), .Y(n123) );
  AND2X1 U295 ( .A(n1810), .B(n98), .Y(n124) );
  INVX1 U296 ( .A(n124), .Y(n125) );
  AND2X1 U297 ( .A(n1827), .B(n98), .Y(n126) );
  INVX1 U298 ( .A(n126), .Y(n127) );
  AND2X1 U299 ( .A(n1844), .B(n98), .Y(n129) );
  INVX1 U300 ( .A(n129), .Y(n130) );
  AND2X1 U301 ( .A(n1861), .B(n98), .Y(n132) );
  INVX1 U302 ( .A(n132), .Y(n133) );
  AND2X1 U303 ( .A(n95), .B(n1743), .Y(n136) );
  INVX1 U304 ( .A(n136), .Y(n137) );
  AND2X1 U305 ( .A(n97), .B(n1743), .Y(n139) );
  INVX1 U306 ( .A(n139), .Y(n140) );
  AND2X1 U307 ( .A(n1793), .B(n1743), .Y(n141) );
  INVX1 U308 ( .A(n141), .Y(n142) );
  AND2X1 U309 ( .A(n1810), .B(n1743), .Y(n143) );
  INVX1 U310 ( .A(n143), .Y(n144) );
  AND2X1 U311 ( .A(n1827), .B(n1743), .Y(n145) );
  INVX1 U312 ( .A(n145), .Y(n146) );
  AND2X1 U313 ( .A(n1844), .B(n1743), .Y(n147) );
  INVX1 U314 ( .A(n147), .Y(n148) );
  AND2X1 U315 ( .A(n1861), .B(n1743), .Y(n149) );
  INVX1 U316 ( .A(n149), .Y(n150) );
  AND2X1 U317 ( .A(n95), .B(n1878), .Y(n151) );
  INVX1 U318 ( .A(n151), .Y(n152) );
  AND2X1 U319 ( .A(n97), .B(n1878), .Y(n153) );
  INVX1 U320 ( .A(n153), .Y(n154) );
  AND2X1 U321 ( .A(n1793), .B(n1878), .Y(n155) );
  INVX1 U322 ( .A(n155), .Y(n156) );
  AND2X1 U323 ( .A(n1810), .B(n1878), .Y(n157) );
  INVX1 U324 ( .A(n157), .Y(n158) );
  AND2X1 U325 ( .A(n1827), .B(n1878), .Y(n159) );
  INVX1 U326 ( .A(n159), .Y(n160) );
  AND2X1 U327 ( .A(n1844), .B(n1878), .Y(n161) );
  INVX1 U328 ( .A(n161), .Y(n162) );
  AND2X1 U329 ( .A(n1861), .B(n1878), .Y(n164) );
  INVX1 U330 ( .A(n164), .Y(n165) );
  AND2X2 U331 ( .A(n11), .B(n99), .Y(n168) );
  BUFX2 U332 ( .A(n36), .Y(n1259) );
  BUFX2 U333 ( .A(n36), .Y(n1260) );
  BUFX2 U334 ( .A(n34), .Y(n1255) );
  BUFX2 U335 ( .A(n34), .Y(n1256) );
  BUFX2 U336 ( .A(n32), .Y(n1251) );
  BUFX2 U337 ( .A(n32), .Y(n1252) );
  AND2X2 U338 ( .A(n13), .B(n118), .Y(n169) );
  AND2X2 U339 ( .A(n14), .B(n116), .Y(n170) );
  AND2X2 U340 ( .A(n15), .B(n114), .Y(n171) );
  AND2X2 U341 ( .A(n8), .B(n112), .Y(n172) );
  AND2X2 U342 ( .A(n9), .B(n108), .Y(n173) );
  AND2X2 U343 ( .A(n10), .B(n110), .Y(n174) );
  AND2X2 U344 ( .A(n11), .B(n106), .Y(n175) );
  AND2X2 U345 ( .A(n12), .B(n104), .Y(n176) );
  INVX1 U346 ( .A(N11), .Y(n1354) );
  MUX2X1 U347 ( .B(n178), .A(n179), .S(n1195), .Y(n177) );
  MUX2X1 U348 ( .B(n181), .A(n182), .S(n1195), .Y(n180) );
  MUX2X1 U349 ( .B(n184), .A(n185), .S(n1195), .Y(n183) );
  MUX2X1 U350 ( .B(n187), .A(n188), .S(n1195), .Y(n186) );
  MUX2X1 U351 ( .B(n190), .A(n191), .S(n1187), .Y(n189) );
  MUX2X1 U352 ( .B(n193), .A(n194), .S(n1195), .Y(n192) );
  MUX2X1 U353 ( .B(n196), .A(n197), .S(n1195), .Y(n195) );
  MUX2X1 U354 ( .B(n199), .A(n200), .S(n1195), .Y(n198) );
  MUX2X1 U355 ( .B(n202), .A(n203), .S(n1195), .Y(n201) );
  MUX2X1 U356 ( .B(n205), .A(n206), .S(n1187), .Y(n204) );
  MUX2X1 U357 ( .B(n208), .A(n209), .S(n1196), .Y(n207) );
  MUX2X1 U358 ( .B(n211), .A(n212), .S(n1196), .Y(n210) );
  MUX2X1 U359 ( .B(n215), .A(n216), .S(n1196), .Y(n213) );
  MUX2X1 U360 ( .B(n218), .A(n219), .S(n1196), .Y(n217) );
  MUX2X1 U361 ( .B(n221), .A(n222), .S(n1187), .Y(n220) );
  MUX2X1 U362 ( .B(n224), .A(n225), .S(n1196), .Y(n223) );
  MUX2X1 U363 ( .B(n227), .A(n228), .S(n1196), .Y(n226) );
  MUX2X1 U364 ( .B(n230), .A(n231), .S(n1196), .Y(n229) );
  MUX2X1 U365 ( .B(n233), .A(n234), .S(n1196), .Y(n232) );
  MUX2X1 U366 ( .B(n236), .A(n237), .S(n1187), .Y(n235) );
  MUX2X1 U367 ( .B(n239), .A(n240), .S(n1196), .Y(n238) );
  MUX2X1 U368 ( .B(n242), .A(n243), .S(n1196), .Y(n241) );
  MUX2X1 U369 ( .B(n245), .A(n246), .S(n1196), .Y(n244) );
  MUX2X1 U370 ( .B(n248), .A(n249), .S(n1196), .Y(n247) );
  MUX2X1 U371 ( .B(n251), .A(n252), .S(n1187), .Y(n250) );
  MUX2X1 U372 ( .B(n254), .A(n255), .S(n1197), .Y(n253) );
  MUX2X1 U373 ( .B(n257), .A(n258), .S(n1197), .Y(n256) );
  MUX2X1 U374 ( .B(n260), .A(n261), .S(n1197), .Y(n259) );
  MUX2X1 U375 ( .B(n263), .A(n264), .S(n1197), .Y(n262) );
  MUX2X1 U376 ( .B(n266), .A(n267), .S(n1187), .Y(n265) );
  MUX2X1 U377 ( .B(n269), .A(n270), .S(n1197), .Y(n268) );
  MUX2X1 U378 ( .B(n272), .A(n273), .S(n1197), .Y(n271) );
  MUX2X1 U379 ( .B(n275), .A(n276), .S(n1197), .Y(n274) );
  MUX2X1 U380 ( .B(n278), .A(n279), .S(n1197), .Y(n277) );
  MUX2X1 U381 ( .B(n281), .A(n282), .S(n1187), .Y(n280) );
  MUX2X1 U382 ( .B(n284), .A(n285), .S(n1197), .Y(n283) );
  MUX2X1 U383 ( .B(n287), .A(n288), .S(n1197), .Y(n286) );
  MUX2X1 U384 ( .B(n290), .A(n291), .S(n1197), .Y(n289) );
  MUX2X1 U385 ( .B(n293), .A(n294), .S(n1197), .Y(n292) );
  MUX2X1 U386 ( .B(n296), .A(n297), .S(n1187), .Y(n295) );
  MUX2X1 U387 ( .B(n299), .A(n300), .S(n1198), .Y(n298) );
  MUX2X1 U388 ( .B(n302), .A(n303), .S(n1198), .Y(n301) );
  MUX2X1 U389 ( .B(n305), .A(n306), .S(n1198), .Y(n304) );
  MUX2X1 U390 ( .B(n308), .A(n309), .S(n1198), .Y(n307) );
  MUX2X1 U391 ( .B(n311), .A(n312), .S(n1187), .Y(n310) );
  MUX2X1 U392 ( .B(n314), .A(n315), .S(n1198), .Y(n313) );
  MUX2X1 U393 ( .B(n317), .A(n318), .S(n1198), .Y(n316) );
  MUX2X1 U394 ( .B(n320), .A(n321), .S(n1198), .Y(n319) );
  MUX2X1 U395 ( .B(n323), .A(n324), .S(n1198), .Y(n322) );
  MUX2X1 U396 ( .B(n326), .A(n327), .S(n1187), .Y(n325) );
  MUX2X1 U397 ( .B(n329), .A(n330), .S(n1198), .Y(n328) );
  MUX2X1 U398 ( .B(n332), .A(n333), .S(n1198), .Y(n331) );
  MUX2X1 U399 ( .B(n335), .A(n336), .S(n1198), .Y(n334) );
  MUX2X1 U400 ( .B(n338), .A(n339), .S(n1198), .Y(n337) );
  MUX2X1 U401 ( .B(n341), .A(n342), .S(n1187), .Y(n340) );
  MUX2X1 U402 ( .B(n344), .A(n345), .S(n1199), .Y(n343) );
  MUX2X1 U403 ( .B(n347), .A(n348), .S(n1199), .Y(n346) );
  MUX2X1 U404 ( .B(n350), .A(n351), .S(n1199), .Y(n349) );
  MUX2X1 U405 ( .B(n353), .A(n354), .S(n1199), .Y(n352) );
  MUX2X1 U406 ( .B(n356), .A(n357), .S(n1187), .Y(n355) );
  MUX2X1 U407 ( .B(n359), .A(n360), .S(n1199), .Y(n358) );
  MUX2X1 U408 ( .B(n362), .A(n363), .S(n1199), .Y(n361) );
  MUX2X1 U409 ( .B(n365), .A(n366), .S(n1199), .Y(n364) );
  MUX2X1 U410 ( .B(n368), .A(n369), .S(n1199), .Y(n367) );
  MUX2X1 U411 ( .B(n371), .A(n372), .S(n1356), .Y(n370) );
  MUX2X1 U412 ( .B(n374), .A(n375), .S(n1199), .Y(n373) );
  MUX2X1 U413 ( .B(n377), .A(n378), .S(n1199), .Y(n376) );
  MUX2X1 U414 ( .B(n380), .A(n381), .S(n1199), .Y(n379) );
  MUX2X1 U415 ( .B(n383), .A(n384), .S(n1199), .Y(n382) );
  MUX2X1 U416 ( .B(n386), .A(n387), .S(n1356), .Y(n385) );
  MUX2X1 U417 ( .B(n389), .A(n390), .S(n1200), .Y(n388) );
  MUX2X1 U418 ( .B(n392), .A(n393), .S(n1200), .Y(n391) );
  MUX2X1 U419 ( .B(n395), .A(n396), .S(n1200), .Y(n394) );
  MUX2X1 U420 ( .B(n398), .A(n399), .S(n1200), .Y(n397) );
  MUX2X1 U421 ( .B(n401), .A(n402), .S(n1356), .Y(n400) );
  MUX2X1 U422 ( .B(n404), .A(n405), .S(n1200), .Y(n403) );
  MUX2X1 U423 ( .B(n407), .A(n408), .S(n1200), .Y(n406) );
  MUX2X1 U424 ( .B(n410), .A(n411), .S(n1200), .Y(n409) );
  MUX2X1 U425 ( .B(n413), .A(n414), .S(n1200), .Y(n412) );
  MUX2X1 U426 ( .B(n416), .A(n417), .S(n1356), .Y(n415) );
  MUX2X1 U427 ( .B(n419), .A(n420), .S(n1200), .Y(n418) );
  MUX2X1 U428 ( .B(n422), .A(n423), .S(n1200), .Y(n421) );
  MUX2X1 U429 ( .B(n425), .A(n426), .S(n1200), .Y(n424) );
  MUX2X1 U430 ( .B(n428), .A(n429), .S(n1200), .Y(n427) );
  MUX2X1 U431 ( .B(n431), .A(n432), .S(n1356), .Y(n430) );
  MUX2X1 U432 ( .B(n434), .A(n435), .S(n1201), .Y(n433) );
  MUX2X1 U433 ( .B(n437), .A(n438), .S(n1201), .Y(n436) );
  MUX2X1 U434 ( .B(n440), .A(n441), .S(n1201), .Y(n439) );
  MUX2X1 U435 ( .B(n443), .A(n444), .S(n1201), .Y(n442) );
  MUX2X1 U436 ( .B(n446), .A(n447), .S(n1356), .Y(n445) );
  MUX2X1 U437 ( .B(n449), .A(n450), .S(n1201), .Y(n448) );
  MUX2X1 U438 ( .B(n452), .A(n453), .S(n1201), .Y(n451) );
  MUX2X1 U439 ( .B(n455), .A(n456), .S(n1201), .Y(n454) );
  MUX2X1 U440 ( .B(n458), .A(n459), .S(n1201), .Y(n457) );
  MUX2X1 U441 ( .B(n461), .A(n462), .S(n1356), .Y(n460) );
  MUX2X1 U442 ( .B(n464), .A(n465), .S(n1201), .Y(n463) );
  MUX2X1 U443 ( .B(n467), .A(n468), .S(n1201), .Y(n466) );
  MUX2X1 U444 ( .B(n470), .A(n471), .S(n1201), .Y(n469) );
  MUX2X1 U445 ( .B(n473), .A(n474), .S(n1201), .Y(n472) );
  MUX2X1 U446 ( .B(n476), .A(n477), .S(n1356), .Y(n475) );
  MUX2X1 U447 ( .B(n479), .A(n480), .S(n1202), .Y(n478) );
  MUX2X1 U448 ( .B(n482), .A(n483), .S(n1202), .Y(n481) );
  MUX2X1 U449 ( .B(n485), .A(n486), .S(n1202), .Y(n484) );
  MUX2X1 U450 ( .B(n488), .A(n489), .S(n1202), .Y(n487) );
  MUX2X1 U451 ( .B(n491), .A(n492), .S(n1356), .Y(n490) );
  MUX2X1 U452 ( .B(n494), .A(n495), .S(n1202), .Y(n493) );
  MUX2X1 U453 ( .B(n497), .A(n498), .S(n1202), .Y(n496) );
  MUX2X1 U454 ( .B(n500), .A(n501), .S(n1202), .Y(n499) );
  MUX2X1 U455 ( .B(n503), .A(n504), .S(n1202), .Y(n502) );
  MUX2X1 U456 ( .B(n506), .A(n507), .S(n1356), .Y(n505) );
  MUX2X1 U457 ( .B(n509), .A(n510), .S(n1202), .Y(n508) );
  MUX2X1 U458 ( .B(n512), .A(n513), .S(n1202), .Y(n511) );
  MUX2X1 U459 ( .B(n515), .A(n516), .S(n1202), .Y(n514) );
  MUX2X1 U460 ( .B(n518), .A(n519), .S(n1202), .Y(n517) );
  MUX2X1 U461 ( .B(n521), .A(n522), .S(n1356), .Y(n520) );
  MUX2X1 U462 ( .B(n524), .A(n525), .S(n1203), .Y(n523) );
  MUX2X1 U463 ( .B(n527), .A(n528), .S(n1203), .Y(n526) );
  MUX2X1 U464 ( .B(n530), .A(n531), .S(n1203), .Y(n529) );
  MUX2X1 U465 ( .B(n533), .A(n534), .S(n1203), .Y(n532) );
  MUX2X1 U466 ( .B(n536), .A(n537), .S(n1356), .Y(n535) );
  MUX2X1 U467 ( .B(n539), .A(n540), .S(n1203), .Y(n538) );
  MUX2X1 U468 ( .B(n542), .A(n543), .S(n1203), .Y(n541) );
  MUX2X1 U469 ( .B(n545), .A(n546), .S(n1203), .Y(n544) );
  MUX2X1 U470 ( .B(n548), .A(n549), .S(n1203), .Y(n547) );
  MUX2X1 U471 ( .B(n551), .A(n552), .S(n1356), .Y(n550) );
  MUX2X1 U472 ( .B(n554), .A(n555), .S(n1203), .Y(n553) );
  MUX2X1 U473 ( .B(n557), .A(n558), .S(n1203), .Y(n556) );
  MUX2X1 U474 ( .B(n560), .A(n561), .S(n1203), .Y(n559) );
  MUX2X1 U475 ( .B(n563), .A(n564), .S(n1203), .Y(n562) );
  MUX2X1 U476 ( .B(n566), .A(n567), .S(n1356), .Y(n565) );
  MUX2X1 U477 ( .B(n569), .A(n570), .S(n1204), .Y(n568) );
  MUX2X1 U478 ( .B(n572), .A(n573), .S(n1204), .Y(n571) );
  MUX2X1 U479 ( .B(n575), .A(n576), .S(n1204), .Y(n574) );
  MUX2X1 U480 ( .B(n578), .A(n579), .S(n1204), .Y(n577) );
  MUX2X1 U481 ( .B(n581), .A(n582), .S(n1187), .Y(n580) );
  MUX2X1 U482 ( .B(n584), .A(n585), .S(n1204), .Y(n583) );
  MUX2X1 U483 ( .B(n587), .A(n588), .S(n1204), .Y(n586) );
  MUX2X1 U484 ( .B(n590), .A(n591), .S(n1204), .Y(n589) );
  MUX2X1 U485 ( .B(n593), .A(n594), .S(n1204), .Y(n592) );
  MUX2X1 U486 ( .B(n596), .A(n597), .S(n1187), .Y(n595) );
  MUX2X1 U487 ( .B(n599), .A(n600), .S(n1204), .Y(n598) );
  MUX2X1 U488 ( .B(n602), .A(n603), .S(n1204), .Y(n601) );
  MUX2X1 U489 ( .B(n605), .A(n606), .S(n1204), .Y(n604) );
  MUX2X1 U490 ( .B(n608), .A(n609), .S(n1204), .Y(n607) );
  MUX2X1 U491 ( .B(n611), .A(n612), .S(n1356), .Y(n610) );
  MUX2X1 U492 ( .B(n614), .A(n615), .S(n1205), .Y(n613) );
  MUX2X1 U493 ( .B(n617), .A(n618), .S(n1205), .Y(n616) );
  MUX2X1 U494 ( .B(n620), .A(n621), .S(n1205), .Y(n619) );
  MUX2X1 U495 ( .B(n623), .A(n624), .S(n1205), .Y(n622) );
  MUX2X1 U496 ( .B(n626), .A(n627), .S(n1187), .Y(n625) );
  MUX2X1 U497 ( .B(n629), .A(n630), .S(n1205), .Y(n628) );
  MUX2X1 U498 ( .B(n632), .A(n633), .S(n1205), .Y(n631) );
  MUX2X1 U499 ( .B(n635), .A(n636), .S(n1205), .Y(n634) );
  MUX2X1 U500 ( .B(n638), .A(n639), .S(n1205), .Y(n637) );
  MUX2X1 U501 ( .B(n641), .A(n642), .S(n1187), .Y(n640) );
  MUX2X1 U502 ( .B(n644), .A(n645), .S(n1205), .Y(n643) );
  MUX2X1 U503 ( .B(n647), .A(n648), .S(n1205), .Y(n646) );
  MUX2X1 U504 ( .B(n650), .A(n1163), .S(n1205), .Y(n649) );
  MUX2X1 U505 ( .B(n1165), .A(n1166), .S(n1205), .Y(n1164) );
  MUX2X1 U506 ( .B(n1168), .A(n1169), .S(n1187), .Y(n1167) );
  MUX2X1 U507 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1223), .Y(n179) );
  MUX2X1 U508 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1224), .Y(n178) );
  MUX2X1 U509 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1215), .Y(n182) );
  MUX2X1 U510 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1214), .Y(n181) );
  MUX2X1 U511 ( .B(n180), .A(n177), .S(n1192), .Y(n191) );
  MUX2X1 U512 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1212), .Y(n185) );
  MUX2X1 U513 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1212), .Y(n184) );
  MUX2X1 U514 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1212), .Y(n188) );
  MUX2X1 U515 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1212), .Y(n187) );
  MUX2X1 U516 ( .B(n186), .A(n183), .S(n1192), .Y(n190) );
  MUX2X1 U517 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1212), .Y(n194) );
  MUX2X1 U518 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1212), .Y(n193) );
  MUX2X1 U519 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1212), .Y(n197) );
  MUX2X1 U520 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1212), .Y(n196) );
  MUX2X1 U521 ( .B(n195), .A(n192), .S(n1192), .Y(n206) );
  MUX2X1 U522 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1212), .Y(n200) );
  MUX2X1 U523 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1212), .Y(n199) );
  MUX2X1 U524 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1212), .Y(n203) );
  MUX2X1 U525 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1212), .Y(n202) );
  MUX2X1 U526 ( .B(n201), .A(n198), .S(n1192), .Y(n205) );
  MUX2X1 U527 ( .B(n204), .A(n189), .S(n1186), .Y(n1170) );
  MUX2X1 U528 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1213), .Y(n209) );
  MUX2X1 U529 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1213), .Y(n208) );
  MUX2X1 U530 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1213), .Y(n212) );
  MUX2X1 U531 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1213), .Y(n211) );
  MUX2X1 U532 ( .B(n210), .A(n207), .S(n1192), .Y(n222) );
  MUX2X1 U533 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1213), .Y(n216) );
  MUX2X1 U534 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1213), .Y(n215) );
  MUX2X1 U535 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1213), .Y(n219) );
  MUX2X1 U536 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1213), .Y(n218) );
  MUX2X1 U537 ( .B(n217), .A(n213), .S(n1192), .Y(n221) );
  MUX2X1 U538 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1213), .Y(n225) );
  MUX2X1 U539 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1213), .Y(n224) );
  MUX2X1 U540 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1213), .Y(n228) );
  MUX2X1 U541 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1213), .Y(n227) );
  MUX2X1 U542 ( .B(n226), .A(n223), .S(n1192), .Y(n237) );
  MUX2X1 U543 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1214), .Y(n231) );
  MUX2X1 U544 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1214), .Y(n230) );
  MUX2X1 U545 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1214), .Y(n234) );
  MUX2X1 U546 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1214), .Y(n233) );
  MUX2X1 U547 ( .B(n232), .A(n229), .S(n1192), .Y(n236) );
  MUX2X1 U548 ( .B(n235), .A(n220), .S(n1186), .Y(n1171) );
  MUX2X1 U549 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1214), .Y(n240) );
  MUX2X1 U550 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1214), .Y(n239) );
  MUX2X1 U551 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1214), .Y(n243) );
  MUX2X1 U552 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1214), .Y(n242) );
  MUX2X1 U553 ( .B(n241), .A(n238), .S(n1192), .Y(n252) );
  MUX2X1 U554 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1214), .Y(n246) );
  MUX2X1 U555 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1214), .Y(n245) );
  MUX2X1 U556 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1214), .Y(n249) );
  MUX2X1 U557 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1214), .Y(n248) );
  MUX2X1 U558 ( .B(n247), .A(n244), .S(n1192), .Y(n251) );
  MUX2X1 U559 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1215), .Y(n255) );
  MUX2X1 U560 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1215), .Y(n254) );
  MUX2X1 U561 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1215), .Y(n258) );
  MUX2X1 U562 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1215), .Y(n257) );
  MUX2X1 U563 ( .B(n256), .A(n253), .S(n1192), .Y(n267) );
  MUX2X1 U564 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1215), .Y(n261) );
  MUX2X1 U565 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1215), .Y(n260) );
  MUX2X1 U566 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1215), .Y(n264) );
  MUX2X1 U567 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1215), .Y(n263) );
  MUX2X1 U568 ( .B(n262), .A(n259), .S(n1192), .Y(n266) );
  MUX2X1 U569 ( .B(n265), .A(n250), .S(n1186), .Y(n1172) );
  MUX2X1 U570 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1215), .Y(n270) );
  MUX2X1 U571 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1215), .Y(n269) );
  MUX2X1 U572 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1215), .Y(n273) );
  MUX2X1 U573 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1215), .Y(n272) );
  MUX2X1 U574 ( .B(n271), .A(n268), .S(n1191), .Y(n282) );
  MUX2X1 U575 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1216), .Y(n276) );
  MUX2X1 U576 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1216), .Y(n275) );
  MUX2X1 U577 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1216), .Y(n279) );
  MUX2X1 U578 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1216), .Y(n278) );
  MUX2X1 U579 ( .B(n277), .A(n274), .S(n1191), .Y(n281) );
  MUX2X1 U580 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1216), .Y(n285) );
  MUX2X1 U581 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1216), .Y(n284) );
  MUX2X1 U582 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1216), .Y(n288) );
  MUX2X1 U583 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1216), .Y(n287) );
  MUX2X1 U584 ( .B(n286), .A(n283), .S(n1191), .Y(n297) );
  MUX2X1 U585 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1216), .Y(n291) );
  MUX2X1 U586 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1216), .Y(n290) );
  MUX2X1 U587 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1216), .Y(n294) );
  MUX2X1 U588 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1216), .Y(n293) );
  MUX2X1 U589 ( .B(n292), .A(n289), .S(n1191), .Y(n296) );
  MUX2X1 U590 ( .B(n295), .A(n280), .S(n1186), .Y(n1173) );
  MUX2X1 U591 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1217), .Y(n300) );
  MUX2X1 U592 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1217), .Y(n299) );
  MUX2X1 U593 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1217), .Y(n303) );
  MUX2X1 U594 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1217), .Y(n302) );
  MUX2X1 U595 ( .B(n301), .A(n298), .S(n1191), .Y(n312) );
  MUX2X1 U596 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1217), .Y(n306) );
  MUX2X1 U597 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1217), .Y(n305) );
  MUX2X1 U598 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1217), .Y(n309) );
  MUX2X1 U599 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1217), .Y(n308) );
  MUX2X1 U600 ( .B(n307), .A(n304), .S(n1191), .Y(n311) );
  MUX2X1 U601 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1217), .Y(n315) );
  MUX2X1 U602 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1217), .Y(n314) );
  MUX2X1 U603 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1217), .Y(n318) );
  MUX2X1 U604 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1217), .Y(n317) );
  MUX2X1 U605 ( .B(n316), .A(n313), .S(n1191), .Y(n327) );
  MUX2X1 U606 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1218), .Y(n321) );
  MUX2X1 U607 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1218), .Y(n320) );
  MUX2X1 U608 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1218), .Y(n324) );
  MUX2X1 U609 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1218), .Y(n323) );
  MUX2X1 U610 ( .B(n322), .A(n319), .S(n1191), .Y(n326) );
  MUX2X1 U611 ( .B(n325), .A(n310), .S(n1186), .Y(n1174) );
  MUX2X1 U612 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1218), .Y(n330) );
  MUX2X1 U613 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1218), .Y(n329) );
  MUX2X1 U614 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1218), .Y(n333) );
  MUX2X1 U615 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1218), .Y(n332) );
  MUX2X1 U616 ( .B(n331), .A(n328), .S(n1191), .Y(n342) );
  MUX2X1 U617 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1218), .Y(n336) );
  MUX2X1 U618 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1218), .Y(n335) );
  MUX2X1 U619 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1218), .Y(n339) );
  MUX2X1 U620 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1218), .Y(n338) );
  MUX2X1 U621 ( .B(n337), .A(n334), .S(n1191), .Y(n341) );
  MUX2X1 U622 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1219), .Y(n345) );
  MUX2X1 U623 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1219), .Y(n344) );
  MUX2X1 U624 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1219), .Y(n348) );
  MUX2X1 U625 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1219), .Y(n347) );
  MUX2X1 U626 ( .B(n346), .A(n343), .S(n1191), .Y(n357) );
  MUX2X1 U627 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1219), .Y(n351) );
  MUX2X1 U628 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1219), .Y(n350) );
  MUX2X1 U629 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1219), .Y(n354) );
  MUX2X1 U630 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1219), .Y(n353) );
  MUX2X1 U631 ( .B(n352), .A(n349), .S(n1191), .Y(n356) );
  MUX2X1 U632 ( .B(n355), .A(n340), .S(n1186), .Y(n1175) );
  MUX2X1 U633 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1219), .Y(n360) );
  MUX2X1 U634 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1219), .Y(n359) );
  MUX2X1 U635 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1219), .Y(n363) );
  MUX2X1 U636 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1219), .Y(n362) );
  MUX2X1 U637 ( .B(n361), .A(n358), .S(n1190), .Y(n372) );
  MUX2X1 U638 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1220), .Y(n366) );
  MUX2X1 U639 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1220), .Y(n365) );
  MUX2X1 U640 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1220), .Y(n369) );
  MUX2X1 U641 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1220), .Y(n368) );
  MUX2X1 U642 ( .B(n367), .A(n364), .S(n1190), .Y(n371) );
  MUX2X1 U643 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1220), .Y(n375) );
  MUX2X1 U644 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1220), .Y(n374) );
  MUX2X1 U645 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1220), .Y(n378) );
  MUX2X1 U646 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1220), .Y(n377) );
  MUX2X1 U647 ( .B(n376), .A(n373), .S(n1190), .Y(n387) );
  MUX2X1 U648 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1220), .Y(n381) );
  MUX2X1 U649 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1220), .Y(n380) );
  MUX2X1 U650 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1220), .Y(n384) );
  MUX2X1 U651 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1220), .Y(n383) );
  MUX2X1 U652 ( .B(n382), .A(n379), .S(n1190), .Y(n386) );
  MUX2X1 U653 ( .B(n385), .A(n370), .S(n1186), .Y(n1176) );
  MUX2X1 U654 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1221), .Y(n390) );
  MUX2X1 U655 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1221), .Y(n389) );
  MUX2X1 U656 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1221), .Y(n393) );
  MUX2X1 U657 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1221), .Y(n392) );
  MUX2X1 U658 ( .B(n391), .A(n388), .S(n1190), .Y(n402) );
  MUX2X1 U659 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1221), .Y(n396) );
  MUX2X1 U660 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1221), .Y(n395) );
  MUX2X1 U661 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1221), .Y(n399) );
  MUX2X1 U662 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1221), .Y(n398) );
  MUX2X1 U663 ( .B(n397), .A(n394), .S(n1190), .Y(n401) );
  MUX2X1 U664 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1221), .Y(n405) );
  MUX2X1 U665 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1221), .Y(n404) );
  MUX2X1 U666 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1221), .Y(n408) );
  MUX2X1 U667 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1221), .Y(n407) );
  MUX2X1 U668 ( .B(n406), .A(n403), .S(n1190), .Y(n417) );
  MUX2X1 U669 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1222), .Y(n411) );
  MUX2X1 U670 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1222), .Y(n410) );
  MUX2X1 U671 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1222), .Y(n414) );
  MUX2X1 U672 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1222), .Y(n413) );
  MUX2X1 U673 ( .B(n412), .A(n409), .S(n1190), .Y(n416) );
  MUX2X1 U674 ( .B(n415), .A(n400), .S(n1186), .Y(n1177) );
  MUX2X1 U675 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1222), .Y(n420) );
  MUX2X1 U676 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1222), .Y(n419) );
  MUX2X1 U677 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1222), .Y(n423) );
  MUX2X1 U678 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1222), .Y(n422) );
  MUX2X1 U679 ( .B(n421), .A(n418), .S(n1190), .Y(n432) );
  MUX2X1 U680 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1222), .Y(n426) );
  MUX2X1 U681 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1222), .Y(n425) );
  MUX2X1 U682 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1222), .Y(n429) );
  MUX2X1 U683 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1222), .Y(n428) );
  MUX2X1 U684 ( .B(n427), .A(n424), .S(n1190), .Y(n431) );
  MUX2X1 U685 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1223), .Y(n435) );
  MUX2X1 U686 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1223), .Y(n434) );
  MUX2X1 U687 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1223), .Y(n438) );
  MUX2X1 U688 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1223), .Y(n437) );
  MUX2X1 U689 ( .B(n436), .A(n433), .S(n1190), .Y(n447) );
  MUX2X1 U690 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1223), .Y(n441) );
  MUX2X1 U691 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1223), .Y(n440) );
  MUX2X1 U692 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1223), .Y(n444) );
  MUX2X1 U693 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1223), .Y(n443) );
  MUX2X1 U694 ( .B(n442), .A(n439), .S(n1190), .Y(n446) );
  MUX2X1 U695 ( .B(n445), .A(n430), .S(n1186), .Y(n1178) );
  MUX2X1 U696 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1223), .Y(n450) );
  MUX2X1 U697 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1223), .Y(n449) );
  MUX2X1 U698 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1223), .Y(n453) );
  MUX2X1 U699 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1223), .Y(n452) );
  MUX2X1 U700 ( .B(n451), .A(n448), .S(n1189), .Y(n462) );
  MUX2X1 U701 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1224), .Y(n456) );
  MUX2X1 U702 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1224), .Y(n455) );
  MUX2X1 U703 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1224), .Y(n459) );
  MUX2X1 U704 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1224), .Y(n458) );
  MUX2X1 U705 ( .B(n457), .A(n454), .S(n1189), .Y(n461) );
  MUX2X1 U706 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1224), .Y(n465) );
  MUX2X1 U707 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1224), .Y(n464) );
  MUX2X1 U708 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1224), .Y(n468) );
  MUX2X1 U709 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1224), .Y(n467) );
  MUX2X1 U710 ( .B(n466), .A(n463), .S(n1189), .Y(n477) );
  MUX2X1 U711 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1224), .Y(n471) );
  MUX2X1 U712 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1224), .Y(n470) );
  MUX2X1 U713 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1224), .Y(n474) );
  MUX2X1 U714 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1224), .Y(n473) );
  MUX2X1 U715 ( .B(n472), .A(n469), .S(n1189), .Y(n476) );
  MUX2X1 U716 ( .B(n475), .A(n460), .S(n1186), .Y(n1179) );
  MUX2X1 U717 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1225), .Y(n480) );
  MUX2X1 U718 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1225), .Y(n479) );
  MUX2X1 U719 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1225), .Y(n483) );
  MUX2X1 U720 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1225), .Y(n482) );
  MUX2X1 U721 ( .B(n481), .A(n478), .S(n1189), .Y(n492) );
  MUX2X1 U722 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1225), .Y(n486) );
  MUX2X1 U723 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1225), .Y(n485) );
  MUX2X1 U724 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1225), .Y(n489) );
  MUX2X1 U725 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1225), .Y(n488) );
  MUX2X1 U726 ( .B(n487), .A(n484), .S(n1189), .Y(n491) );
  MUX2X1 U727 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1225), .Y(n495) );
  MUX2X1 U728 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1225), .Y(n494) );
  MUX2X1 U729 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1225), .Y(n498) );
  MUX2X1 U730 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1225), .Y(n497) );
  MUX2X1 U731 ( .B(n496), .A(n493), .S(n1189), .Y(n507) );
  MUX2X1 U732 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1226), .Y(n501) );
  MUX2X1 U733 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1226), .Y(n500) );
  MUX2X1 U734 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1226), .Y(n504) );
  MUX2X1 U735 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1226), .Y(n503) );
  MUX2X1 U736 ( .B(n502), .A(n499), .S(n1189), .Y(n506) );
  MUX2X1 U737 ( .B(n505), .A(n490), .S(n1186), .Y(n1180) );
  MUX2X1 U738 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1226), .Y(n510) );
  MUX2X1 U739 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1226), .Y(n509) );
  MUX2X1 U740 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1226), .Y(n513) );
  MUX2X1 U741 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1226), .Y(n512) );
  MUX2X1 U742 ( .B(n511), .A(n508), .S(n1189), .Y(n522) );
  MUX2X1 U743 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1226), .Y(n516) );
  MUX2X1 U744 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1226), .Y(n515) );
  MUX2X1 U745 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1226), .Y(n519) );
  MUX2X1 U746 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1226), .Y(n518) );
  MUX2X1 U747 ( .B(n517), .A(n514), .S(n1189), .Y(n521) );
  MUX2X1 U748 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1227), .Y(n525) );
  MUX2X1 U749 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1227), .Y(n524) );
  MUX2X1 U750 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1227), .Y(n528) );
  MUX2X1 U751 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1227), .Y(n527) );
  MUX2X1 U752 ( .B(n526), .A(n523), .S(n1189), .Y(n537) );
  MUX2X1 U753 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1227), .Y(n531) );
  MUX2X1 U754 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1227), .Y(n530) );
  MUX2X1 U755 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1227), .Y(n534) );
  MUX2X1 U756 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1227), .Y(n533) );
  MUX2X1 U757 ( .B(n532), .A(n529), .S(n1189), .Y(n536) );
  MUX2X1 U758 ( .B(n535), .A(n520), .S(n1186), .Y(n1181) );
  MUX2X1 U759 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1227), .Y(n540) );
  MUX2X1 U760 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1227), .Y(n539) );
  MUX2X1 U761 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1227), .Y(n543) );
  MUX2X1 U762 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1227), .Y(n542) );
  MUX2X1 U763 ( .B(n541), .A(n538), .S(n1188), .Y(n552) );
  MUX2X1 U764 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1228), .Y(n546) );
  MUX2X1 U765 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1228), .Y(n545) );
  MUX2X1 U766 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1228), .Y(n549) );
  MUX2X1 U767 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1228), .Y(n548) );
  MUX2X1 U768 ( .B(n547), .A(n544), .S(n1188), .Y(n551) );
  MUX2X1 U769 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1228), .Y(n555) );
  MUX2X1 U770 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1228), .Y(n554) );
  MUX2X1 U771 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1228), .Y(n558) );
  MUX2X1 U772 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1228), .Y(n557) );
  MUX2X1 U773 ( .B(n556), .A(n553), .S(n1188), .Y(n567) );
  MUX2X1 U774 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1228), .Y(n561) );
  MUX2X1 U775 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1228), .Y(n560) );
  MUX2X1 U776 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1228), .Y(n564) );
  MUX2X1 U777 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1228), .Y(n563) );
  MUX2X1 U778 ( .B(n562), .A(n559), .S(n1188), .Y(n566) );
  MUX2X1 U779 ( .B(n565), .A(n550), .S(n1186), .Y(n1182) );
  MUX2X1 U780 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1229), .Y(n570) );
  MUX2X1 U781 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1229), .Y(n569) );
  MUX2X1 U782 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1229), .Y(n573) );
  MUX2X1 U783 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1229), .Y(n572) );
  MUX2X1 U784 ( .B(n571), .A(n568), .S(n1188), .Y(n582) );
  MUX2X1 U785 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1229), .Y(n576) );
  MUX2X1 U786 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1229), .Y(n575) );
  MUX2X1 U787 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1229), .Y(n579) );
  MUX2X1 U788 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1229), .Y(n578) );
  MUX2X1 U789 ( .B(n577), .A(n574), .S(n1188), .Y(n581) );
  MUX2X1 U790 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1229), .Y(n585) );
  MUX2X1 U791 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1229), .Y(n584) );
  MUX2X1 U792 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1229), .Y(n588) );
  MUX2X1 U793 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1229), .Y(n587) );
  MUX2X1 U794 ( .B(n586), .A(n583), .S(n1188), .Y(n597) );
  MUX2X1 U795 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1230), .Y(n591) );
  MUX2X1 U796 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1230), .Y(n590) );
  MUX2X1 U797 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1230), .Y(n594) );
  MUX2X1 U798 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1230), .Y(n593) );
  MUX2X1 U799 ( .B(n592), .A(n589), .S(n1188), .Y(n596) );
  MUX2X1 U800 ( .B(n595), .A(n580), .S(n1186), .Y(n1183) );
  MUX2X1 U801 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1230), .Y(n600) );
  MUX2X1 U802 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1230), .Y(n599) );
  MUX2X1 U803 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1230), .Y(n603) );
  MUX2X1 U804 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1230), .Y(n602) );
  MUX2X1 U805 ( .B(n601), .A(n598), .S(n1188), .Y(n612) );
  MUX2X1 U806 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1230), .Y(n606) );
  MUX2X1 U807 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1230), .Y(n605) );
  MUX2X1 U808 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1230), .Y(n609) );
  MUX2X1 U809 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1230), .Y(n608) );
  MUX2X1 U810 ( .B(n607), .A(n604), .S(n1188), .Y(n611) );
  MUX2X1 U811 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1231), .Y(n615) );
  MUX2X1 U812 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1231), .Y(n614) );
  MUX2X1 U813 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1231), .Y(n618) );
  MUX2X1 U814 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1231), .Y(n617) );
  MUX2X1 U815 ( .B(n616), .A(n613), .S(n1188), .Y(n627) );
  MUX2X1 U816 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1231), .Y(n621) );
  MUX2X1 U817 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1231), .Y(n620) );
  MUX2X1 U818 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1231), .Y(n624) );
  MUX2X1 U819 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1231), .Y(n623) );
  MUX2X1 U820 ( .B(n622), .A(n619), .S(n1188), .Y(n626) );
  MUX2X1 U821 ( .B(n625), .A(n610), .S(n1186), .Y(n1184) );
  MUX2X1 U822 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1231), .Y(n630) );
  MUX2X1 U823 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1231), .Y(n629) );
  MUX2X1 U824 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1231), .Y(n633) );
  MUX2X1 U825 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1231), .Y(n632) );
  MUX2X1 U826 ( .B(n631), .A(n628), .S(n1189), .Y(n642) );
  MUX2X1 U827 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1226), .Y(n636) );
  MUX2X1 U828 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1225), .Y(n635) );
  MUX2X1 U829 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1219), .Y(n639) );
  MUX2X1 U830 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1227), .Y(n638) );
  MUX2X1 U831 ( .B(n637), .A(n634), .S(n1188), .Y(n641) );
  MUX2X1 U832 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1219), .Y(n645) );
  MUX2X1 U833 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1214), .Y(n644) );
  MUX2X1 U834 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1232), .Y(n648) );
  MUX2X1 U835 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1218), .Y(n647) );
  MUX2X1 U836 ( .B(n646), .A(n643), .S(n1189), .Y(n1169) );
  MUX2X1 U837 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1219), .Y(n1163) );
  MUX2X1 U838 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1220), .Y(n650) );
  MUX2X1 U839 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1217), .Y(n1166) );
  MUX2X1 U840 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1216), .Y(n1165) );
  MUX2X1 U841 ( .B(n1164), .A(n649), .S(n1189), .Y(n1168) );
  MUX2X1 U842 ( .B(n1167), .A(n640), .S(n1186), .Y(n1185) );
  INVX8 U843 ( .A(n1210), .Y(n1214) );
  INVX8 U844 ( .A(n1210), .Y(n1217) );
  INVX8 U845 ( .A(n1210), .Y(n1218) );
  INVX8 U846 ( .A(n1210), .Y(n1219) );
  INVX1 U847 ( .A(N10), .Y(n1352) );
  INVX8 U848 ( .A(n70), .Y(n1318) );
  INVX8 U849 ( .A(n70), .Y(n1319) );
  INVX8 U850 ( .A(n71), .Y(n1320) );
  INVX8 U851 ( .A(n71), .Y(n1321) );
  INVX8 U852 ( .A(n72), .Y(n1322) );
  INVX8 U853 ( .A(n72), .Y(n1323) );
  INVX8 U854 ( .A(n73), .Y(n1324) );
  INVX8 U855 ( .A(n73), .Y(n1325) );
  INVX8 U856 ( .A(n74), .Y(n1326) );
  INVX8 U857 ( .A(n74), .Y(n1327) );
  INVX8 U858 ( .A(n75), .Y(n1328) );
  INVX8 U859 ( .A(n75), .Y(n1329) );
  INVX8 U860 ( .A(n76), .Y(n1330) );
  INVX8 U861 ( .A(n76), .Y(n1331) );
  INVX8 U862 ( .A(n77), .Y(n1332) );
  INVX8 U863 ( .A(n77), .Y(n1333) );
  INVX8 U864 ( .A(n78), .Y(n1334) );
  INVX8 U865 ( .A(n78), .Y(n1335) );
  INVX8 U866 ( .A(n79), .Y(n1336) );
  INVX8 U867 ( .A(n79), .Y(n1337) );
  INVX8 U868 ( .A(n80), .Y(n1338) );
  INVX8 U869 ( .A(n80), .Y(n1339) );
  INVX8 U870 ( .A(n81), .Y(n1340) );
  INVX8 U871 ( .A(n81), .Y(n1341) );
  INVX8 U872 ( .A(n82), .Y(n1342) );
  INVX8 U873 ( .A(n82), .Y(n1343) );
  INVX8 U874 ( .A(n83), .Y(n1344) );
  INVX8 U875 ( .A(n83), .Y(n1345) );
  INVX8 U876 ( .A(n84), .Y(n1346) );
  INVX8 U877 ( .A(n84), .Y(n1347) );
  INVX8 U878 ( .A(n85), .Y(n1348) );
  INVX8 U879 ( .A(n85), .Y(n1349) );
  AND2X2 U880 ( .A(n28), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U881 ( .A(n30), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U882 ( .A(n28), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U883 ( .A(n28), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U884 ( .A(n30), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U885 ( .A(n28), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U886 ( .A(n27), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U887 ( .A(n27), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U888 ( .A(n28), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U889 ( .A(N23), .B(n30), .Y(\data_out<9> ) );
  AND2X2 U890 ( .A(n27), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U891 ( .A(N21), .B(n30), .Y(\data_out<11> ) );
  AND2X2 U892 ( .A(N20), .B(n30), .Y(\data_out<12> ) );
  AND2X2 U893 ( .A(n28), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U894 ( .A(N18), .B(n30), .Y(\data_out<14> ) );
  AND2X2 U895 ( .A(n28), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U896 ( .A(\mem<31><0> ), .B(n1375), .Y(n1360) );
  OAI21X1 U897 ( .A(n1234), .B(n1318), .C(n1360), .Y(n2407) );
  NAND2X1 U898 ( .A(\mem<31><1> ), .B(n1375), .Y(n1361) );
  OAI21X1 U899 ( .A(n1321), .B(n1233), .C(n1361), .Y(n2406) );
  NAND2X1 U900 ( .A(\mem<31><2> ), .B(n1375), .Y(n1362) );
  OAI21X1 U901 ( .A(n1323), .B(n1233), .C(n1362), .Y(n2405) );
  NAND2X1 U902 ( .A(\mem<31><3> ), .B(n1375), .Y(n1363) );
  OAI21X1 U903 ( .A(n1325), .B(n1233), .C(n1363), .Y(n2404) );
  NAND2X1 U904 ( .A(\mem<31><4> ), .B(n1375), .Y(n1364) );
  OAI21X1 U905 ( .A(n1327), .B(n1233), .C(n1364), .Y(n2403) );
  NAND2X1 U906 ( .A(\mem<31><5> ), .B(n1375), .Y(n1365) );
  OAI21X1 U907 ( .A(n1329), .B(n1233), .C(n1365), .Y(n2402) );
  NAND2X1 U908 ( .A(\mem<31><6> ), .B(n1375), .Y(n1366) );
  OAI21X1 U909 ( .A(n1331), .B(n1233), .C(n1366), .Y(n2401) );
  NAND2X1 U910 ( .A(\mem<31><7> ), .B(n1375), .Y(n1367) );
  OAI21X1 U911 ( .A(n1333), .B(n1233), .C(n1367), .Y(n2400) );
  NAND2X1 U912 ( .A(\mem<31><8> ), .B(n1375), .Y(n1368) );
  OAI21X1 U913 ( .A(n1335), .B(n1233), .C(n1368), .Y(n2399) );
  NAND2X1 U914 ( .A(\mem<31><9> ), .B(n1375), .Y(n1369) );
  OAI21X1 U915 ( .A(n1337), .B(n1234), .C(n1369), .Y(n2398) );
  NAND2X1 U916 ( .A(\mem<31><10> ), .B(n1375), .Y(n1370) );
  OAI21X1 U917 ( .A(n1339), .B(n1234), .C(n1370), .Y(n2397) );
  NAND2X1 U918 ( .A(\mem<31><11> ), .B(n1375), .Y(n1371) );
  OAI21X1 U919 ( .A(n1341), .B(n1234), .C(n1371), .Y(n2396) );
  NAND2X1 U920 ( .A(\mem<31><12> ), .B(n1375), .Y(n1372) );
  OAI21X1 U921 ( .A(n1343), .B(n1234), .C(n1372), .Y(n2395) );
  NAND2X1 U922 ( .A(\mem<31><13> ), .B(n1375), .Y(n1373) );
  OAI21X1 U923 ( .A(n1345), .B(n1234), .C(n1373), .Y(n2394) );
  NAND2X1 U924 ( .A(\mem<31><14> ), .B(n1375), .Y(n1374) );
  OAI21X1 U925 ( .A(n1347), .B(n1234), .C(n1374), .Y(n2393) );
  NAND2X1 U926 ( .A(\mem<31><15> ), .B(n1375), .Y(n1376) );
  OAI21X1 U927 ( .A(n1349), .B(n1234), .C(n1376), .Y(n2392) );
  NAND2X1 U928 ( .A(\mem<30><0> ), .B(n1392), .Y(n1377) );
  OAI21X1 U929 ( .A(n1235), .B(n1318), .C(n1377), .Y(n2391) );
  NAND2X1 U930 ( .A(\mem<30><1> ), .B(n1392), .Y(n1378) );
  OAI21X1 U931 ( .A(n1235), .B(n1321), .C(n1378), .Y(n2390) );
  NAND2X1 U932 ( .A(\mem<30><2> ), .B(n1392), .Y(n1379) );
  OAI21X1 U933 ( .A(n1235), .B(n1323), .C(n1379), .Y(n2389) );
  NAND2X1 U934 ( .A(\mem<30><3> ), .B(n1392), .Y(n1380) );
  OAI21X1 U935 ( .A(n1235), .B(n1325), .C(n1380), .Y(n2388) );
  NAND2X1 U936 ( .A(\mem<30><4> ), .B(n1392), .Y(n1381) );
  OAI21X1 U937 ( .A(n1235), .B(n1327), .C(n1381), .Y(n2387) );
  NAND2X1 U938 ( .A(\mem<30><5> ), .B(n1392), .Y(n1382) );
  OAI21X1 U939 ( .A(n1235), .B(n1329), .C(n1382), .Y(n2386) );
  NAND2X1 U940 ( .A(\mem<30><6> ), .B(n1392), .Y(n1383) );
  OAI21X1 U941 ( .A(n1235), .B(n1331), .C(n1383), .Y(n2385) );
  NAND2X1 U942 ( .A(\mem<30><7> ), .B(n1392), .Y(n1384) );
  OAI21X1 U943 ( .A(n1235), .B(n1333), .C(n1384), .Y(n2384) );
  NAND2X1 U944 ( .A(\mem<30><8> ), .B(n1392), .Y(n1385) );
  OAI21X1 U945 ( .A(n1236), .B(n1335), .C(n1385), .Y(n2383) );
  NAND2X1 U946 ( .A(\mem<30><9> ), .B(n1392), .Y(n1386) );
  OAI21X1 U947 ( .A(n1236), .B(n1337), .C(n1386), .Y(n2382) );
  NAND2X1 U948 ( .A(\mem<30><10> ), .B(n1392), .Y(n1387) );
  OAI21X1 U949 ( .A(n1236), .B(n1339), .C(n1387), .Y(n2381) );
  NAND2X1 U950 ( .A(\mem<30><11> ), .B(n1392), .Y(n1388) );
  OAI21X1 U951 ( .A(n1236), .B(n1341), .C(n1388), .Y(n2380) );
  NAND2X1 U952 ( .A(\mem<30><12> ), .B(n1392), .Y(n1389) );
  OAI21X1 U953 ( .A(n1236), .B(n1343), .C(n1389), .Y(n2379) );
  NAND2X1 U954 ( .A(\mem<30><13> ), .B(n1392), .Y(n1390) );
  OAI21X1 U955 ( .A(n1236), .B(n1345), .C(n1390), .Y(n2378) );
  NAND2X1 U956 ( .A(\mem<30><14> ), .B(n1392), .Y(n1391) );
  OAI21X1 U957 ( .A(n1236), .B(n1347), .C(n1391), .Y(n2377) );
  NAND2X1 U958 ( .A(\mem<30><15> ), .B(n1392), .Y(n1393) );
  OAI21X1 U959 ( .A(n1236), .B(n1349), .C(n1393), .Y(n2376) );
  NAND3X1 U960 ( .A(n1351), .B(n1192), .C(n1354), .Y(n1394) );
  NAND2X1 U961 ( .A(\mem<29><0> ), .B(n1410), .Y(n1395) );
  OAI21X1 U962 ( .A(n1237), .B(n1318), .C(n1395), .Y(n2375) );
  NAND2X1 U963 ( .A(\mem<29><1> ), .B(n1410), .Y(n1396) );
  OAI21X1 U964 ( .A(n1237), .B(n1321), .C(n1396), .Y(n2374) );
  NAND2X1 U965 ( .A(\mem<29><2> ), .B(n1410), .Y(n1397) );
  OAI21X1 U966 ( .A(n1237), .B(n1323), .C(n1397), .Y(n2373) );
  NAND2X1 U967 ( .A(\mem<29><3> ), .B(n1410), .Y(n1398) );
  OAI21X1 U968 ( .A(n1237), .B(n1325), .C(n1398), .Y(n2372) );
  NAND2X1 U969 ( .A(\mem<29><4> ), .B(n1410), .Y(n1399) );
  OAI21X1 U970 ( .A(n1237), .B(n1327), .C(n1399), .Y(n2371) );
  NAND2X1 U971 ( .A(\mem<29><5> ), .B(n1410), .Y(n1400) );
  OAI21X1 U972 ( .A(n1237), .B(n1329), .C(n1400), .Y(n2370) );
  NAND2X1 U973 ( .A(\mem<29><6> ), .B(n1410), .Y(n1401) );
  OAI21X1 U974 ( .A(n1237), .B(n1331), .C(n1401), .Y(n2369) );
  NAND2X1 U975 ( .A(\mem<29><7> ), .B(n1410), .Y(n1402) );
  OAI21X1 U976 ( .A(n1237), .B(n1333), .C(n1402), .Y(n2368) );
  NAND2X1 U977 ( .A(\mem<29><8> ), .B(n1410), .Y(n1403) );
  OAI21X1 U978 ( .A(n1238), .B(n1335), .C(n1403), .Y(n2367) );
  NAND2X1 U979 ( .A(\mem<29><9> ), .B(n1410), .Y(n1404) );
  OAI21X1 U980 ( .A(n1238), .B(n1337), .C(n1404), .Y(n2366) );
  NAND2X1 U981 ( .A(\mem<29><10> ), .B(n1410), .Y(n1405) );
  OAI21X1 U982 ( .A(n1238), .B(n1339), .C(n1405), .Y(n2365) );
  NAND2X1 U983 ( .A(\mem<29><11> ), .B(n1410), .Y(n1406) );
  OAI21X1 U984 ( .A(n1238), .B(n1341), .C(n1406), .Y(n2364) );
  NAND2X1 U985 ( .A(\mem<29><12> ), .B(n1410), .Y(n1407) );
  OAI21X1 U986 ( .A(n1238), .B(n1343), .C(n1407), .Y(n2363) );
  NAND2X1 U987 ( .A(\mem<29><13> ), .B(n1410), .Y(n1408) );
  OAI21X1 U988 ( .A(n1238), .B(n1345), .C(n1408), .Y(n2362) );
  NAND2X1 U989 ( .A(\mem<29><14> ), .B(n1410), .Y(n1409) );
  OAI21X1 U990 ( .A(n1238), .B(n1347), .C(n1409), .Y(n2361) );
  NAND2X1 U991 ( .A(\mem<29><15> ), .B(n1410), .Y(n1411) );
  OAI21X1 U992 ( .A(n1238), .B(n1349), .C(n1411), .Y(n2360) );
  NAND3X1 U993 ( .A(n1192), .B(n1354), .C(n1352), .Y(n1412) );
  NAND2X1 U994 ( .A(\mem<28><0> ), .B(n1428), .Y(n1413) );
  OAI21X1 U995 ( .A(n1239), .B(n1318), .C(n1413), .Y(n2359) );
  NAND2X1 U996 ( .A(\mem<28><1> ), .B(n1428), .Y(n1414) );
  OAI21X1 U997 ( .A(n1239), .B(n1321), .C(n1414), .Y(n2358) );
  NAND2X1 U998 ( .A(\mem<28><2> ), .B(n1428), .Y(n1415) );
  OAI21X1 U999 ( .A(n1239), .B(n1323), .C(n1415), .Y(n2357) );
  NAND2X1 U1000 ( .A(\mem<28><3> ), .B(n1428), .Y(n1416) );
  OAI21X1 U1001 ( .A(n1239), .B(n1325), .C(n1416), .Y(n2356) );
  NAND2X1 U1002 ( .A(\mem<28><4> ), .B(n1428), .Y(n1417) );
  OAI21X1 U1003 ( .A(n1239), .B(n1327), .C(n1417), .Y(n2355) );
  NAND2X1 U1004 ( .A(\mem<28><5> ), .B(n1428), .Y(n1418) );
  OAI21X1 U1005 ( .A(n1239), .B(n1329), .C(n1418), .Y(n2354) );
  NAND2X1 U1006 ( .A(\mem<28><6> ), .B(n1428), .Y(n1419) );
  OAI21X1 U1007 ( .A(n1239), .B(n1331), .C(n1419), .Y(n2353) );
  NAND2X1 U1008 ( .A(\mem<28><7> ), .B(n1428), .Y(n1420) );
  OAI21X1 U1009 ( .A(n1239), .B(n1333), .C(n1420), .Y(n2352) );
  NAND2X1 U1010 ( .A(\mem<28><8> ), .B(n1428), .Y(n1421) );
  OAI21X1 U1011 ( .A(n1240), .B(n1335), .C(n1421), .Y(n2351) );
  NAND2X1 U1012 ( .A(\mem<28><9> ), .B(n1428), .Y(n1422) );
  OAI21X1 U1013 ( .A(n1240), .B(n1337), .C(n1422), .Y(n2350) );
  NAND2X1 U1014 ( .A(\mem<28><10> ), .B(n1428), .Y(n1423) );
  OAI21X1 U1015 ( .A(n1240), .B(n1339), .C(n1423), .Y(n2349) );
  NAND2X1 U1016 ( .A(\mem<28><11> ), .B(n1428), .Y(n1424) );
  OAI21X1 U1017 ( .A(n1240), .B(n1341), .C(n1424), .Y(n2348) );
  NAND2X1 U1018 ( .A(\mem<28><12> ), .B(n1428), .Y(n1425) );
  OAI21X1 U1019 ( .A(n1240), .B(n1343), .C(n1425), .Y(n2347) );
  NAND2X1 U1020 ( .A(\mem<28><13> ), .B(n1428), .Y(n1426) );
  OAI21X1 U1021 ( .A(n1240), .B(n1345), .C(n1426), .Y(n2346) );
  NAND2X1 U1022 ( .A(\mem<28><14> ), .B(n1428), .Y(n1427) );
  OAI21X1 U1023 ( .A(n1240), .B(n1347), .C(n1427), .Y(n2345) );
  NAND2X1 U1024 ( .A(\mem<28><15> ), .B(n1428), .Y(n1429) );
  OAI21X1 U1025 ( .A(n1240), .B(n1349), .C(n1429), .Y(n2344) );
  NAND3X1 U1026 ( .A(n1351), .B(n1353), .C(n1355), .Y(n1430) );
  NAND2X1 U1027 ( .A(\mem<27><0> ), .B(n1446), .Y(n1431) );
  OAI21X1 U1028 ( .A(n1241), .B(n1318), .C(n1431), .Y(n2343) );
  NAND2X1 U1029 ( .A(\mem<27><1> ), .B(n1446), .Y(n1432) );
  OAI21X1 U1030 ( .A(n1241), .B(n1321), .C(n1432), .Y(n2342) );
  NAND2X1 U1031 ( .A(\mem<27><2> ), .B(n1446), .Y(n1433) );
  OAI21X1 U1032 ( .A(n1241), .B(n1323), .C(n1433), .Y(n2341) );
  NAND2X1 U1033 ( .A(\mem<27><3> ), .B(n1446), .Y(n1434) );
  OAI21X1 U1034 ( .A(n1241), .B(n1325), .C(n1434), .Y(n2340) );
  NAND2X1 U1035 ( .A(\mem<27><4> ), .B(n1446), .Y(n1435) );
  OAI21X1 U1036 ( .A(n1241), .B(n1327), .C(n1435), .Y(n2339) );
  NAND2X1 U1037 ( .A(\mem<27><5> ), .B(n1446), .Y(n1436) );
  OAI21X1 U1038 ( .A(n1241), .B(n1329), .C(n1436), .Y(n2338) );
  NAND2X1 U1039 ( .A(\mem<27><6> ), .B(n1446), .Y(n1437) );
  OAI21X1 U1040 ( .A(n1241), .B(n1331), .C(n1437), .Y(n2337) );
  NAND2X1 U1041 ( .A(\mem<27><7> ), .B(n1446), .Y(n1438) );
  OAI21X1 U1042 ( .A(n1241), .B(n1333), .C(n1438), .Y(n2336) );
  NAND2X1 U1043 ( .A(\mem<27><8> ), .B(n1446), .Y(n1439) );
  OAI21X1 U1044 ( .A(n1242), .B(n1335), .C(n1439), .Y(n2335) );
  NAND2X1 U1045 ( .A(\mem<27><9> ), .B(n1446), .Y(n1440) );
  OAI21X1 U1046 ( .A(n1242), .B(n1337), .C(n1440), .Y(n2334) );
  NAND2X1 U1047 ( .A(\mem<27><10> ), .B(n1446), .Y(n1441) );
  OAI21X1 U1048 ( .A(n1242), .B(n1339), .C(n1441), .Y(n2333) );
  NAND2X1 U1049 ( .A(\mem<27><11> ), .B(n1446), .Y(n1442) );
  OAI21X1 U1050 ( .A(n1242), .B(n1341), .C(n1442), .Y(n2332) );
  NAND2X1 U1051 ( .A(\mem<27><12> ), .B(n1446), .Y(n1443) );
  OAI21X1 U1052 ( .A(n1242), .B(n1343), .C(n1443), .Y(n2331) );
  NAND2X1 U1053 ( .A(\mem<27><13> ), .B(n1446), .Y(n1444) );
  OAI21X1 U1054 ( .A(n1242), .B(n1345), .C(n1444), .Y(n2330) );
  NAND2X1 U1055 ( .A(\mem<27><14> ), .B(n1446), .Y(n1445) );
  OAI21X1 U1056 ( .A(n1242), .B(n1347), .C(n1445), .Y(n2329) );
  NAND2X1 U1057 ( .A(\mem<27><15> ), .B(n1446), .Y(n1447) );
  OAI21X1 U1058 ( .A(n1242), .B(n1349), .C(n1447), .Y(n2328) );
  NAND3X1 U1059 ( .A(n1355), .B(n1353), .C(n1352), .Y(n1448) );
  NAND2X1 U1060 ( .A(\mem<26><0> ), .B(n1464), .Y(n1449) );
  OAI21X1 U1061 ( .A(n1243), .B(n1318), .C(n1449), .Y(n2327) );
  NAND2X1 U1062 ( .A(\mem<26><1> ), .B(n1464), .Y(n1450) );
  OAI21X1 U1063 ( .A(n1243), .B(n1321), .C(n1450), .Y(n2326) );
  NAND2X1 U1064 ( .A(\mem<26><2> ), .B(n1464), .Y(n1451) );
  OAI21X1 U1065 ( .A(n1243), .B(n1323), .C(n1451), .Y(n2325) );
  NAND2X1 U1066 ( .A(\mem<26><3> ), .B(n1464), .Y(n1452) );
  OAI21X1 U1067 ( .A(n1243), .B(n1325), .C(n1452), .Y(n2324) );
  NAND2X1 U1068 ( .A(\mem<26><4> ), .B(n1464), .Y(n1453) );
  OAI21X1 U1069 ( .A(n1243), .B(n1327), .C(n1453), .Y(n2323) );
  NAND2X1 U1070 ( .A(\mem<26><5> ), .B(n1464), .Y(n1454) );
  OAI21X1 U1071 ( .A(n1243), .B(n1329), .C(n1454), .Y(n2322) );
  NAND2X1 U1072 ( .A(\mem<26><6> ), .B(n1464), .Y(n1455) );
  OAI21X1 U1073 ( .A(n1243), .B(n1331), .C(n1455), .Y(n2321) );
  NAND2X1 U1074 ( .A(\mem<26><7> ), .B(n1464), .Y(n1456) );
  OAI21X1 U1075 ( .A(n1243), .B(n1333), .C(n1456), .Y(n2320) );
  NAND2X1 U1076 ( .A(\mem<26><8> ), .B(n1464), .Y(n1457) );
  OAI21X1 U1077 ( .A(n1244), .B(n1335), .C(n1457), .Y(n2319) );
  NAND2X1 U1078 ( .A(\mem<26><9> ), .B(n1464), .Y(n1458) );
  OAI21X1 U1079 ( .A(n1244), .B(n1337), .C(n1458), .Y(n2318) );
  NAND2X1 U1080 ( .A(\mem<26><10> ), .B(n1464), .Y(n1459) );
  OAI21X1 U1081 ( .A(n1244), .B(n1339), .C(n1459), .Y(n2317) );
  NAND2X1 U1082 ( .A(\mem<26><11> ), .B(n1464), .Y(n1460) );
  OAI21X1 U1083 ( .A(n1244), .B(n1341), .C(n1460), .Y(n2316) );
  NAND2X1 U1084 ( .A(\mem<26><12> ), .B(n1464), .Y(n1461) );
  OAI21X1 U1085 ( .A(n1244), .B(n1343), .C(n1461), .Y(n2315) );
  NAND2X1 U1086 ( .A(\mem<26><13> ), .B(n1464), .Y(n1462) );
  OAI21X1 U1087 ( .A(n1244), .B(n1345), .C(n1462), .Y(n2314) );
  NAND2X1 U1088 ( .A(\mem<26><14> ), .B(n1464), .Y(n1463) );
  OAI21X1 U1089 ( .A(n1244), .B(n1347), .C(n1463), .Y(n2313) );
  NAND2X1 U1090 ( .A(\mem<26><15> ), .B(n1464), .Y(n1465) );
  OAI21X1 U1091 ( .A(n1244), .B(n1349), .C(n1465), .Y(n2312) );
  NAND3X1 U1092 ( .A(n1351), .B(n1355), .C(n1354), .Y(n1466) );
  NAND2X1 U1093 ( .A(\mem<25><0> ), .B(n1482), .Y(n1467) );
  OAI21X1 U1094 ( .A(n1245), .B(n1318), .C(n1467), .Y(n2311) );
  NAND2X1 U1095 ( .A(\mem<25><1> ), .B(n1482), .Y(n1468) );
  OAI21X1 U1096 ( .A(n1245), .B(n1321), .C(n1468), .Y(n2310) );
  NAND2X1 U1097 ( .A(\mem<25><2> ), .B(n1482), .Y(n1469) );
  OAI21X1 U1098 ( .A(n1245), .B(n1323), .C(n1469), .Y(n2309) );
  NAND2X1 U1099 ( .A(\mem<25><3> ), .B(n1482), .Y(n1470) );
  OAI21X1 U1100 ( .A(n1245), .B(n1325), .C(n1470), .Y(n2308) );
  NAND2X1 U1101 ( .A(\mem<25><4> ), .B(n1482), .Y(n1471) );
  OAI21X1 U1102 ( .A(n1245), .B(n1327), .C(n1471), .Y(n2307) );
  NAND2X1 U1103 ( .A(\mem<25><5> ), .B(n1482), .Y(n1472) );
  OAI21X1 U1104 ( .A(n1245), .B(n1329), .C(n1472), .Y(n2306) );
  NAND2X1 U1105 ( .A(\mem<25><6> ), .B(n1482), .Y(n1473) );
  OAI21X1 U1106 ( .A(n1245), .B(n1331), .C(n1473), .Y(n2305) );
  NAND2X1 U1107 ( .A(\mem<25><7> ), .B(n1482), .Y(n1474) );
  OAI21X1 U1108 ( .A(n1245), .B(n1333), .C(n1474), .Y(n2304) );
  NAND2X1 U1109 ( .A(\mem<25><8> ), .B(n1482), .Y(n1475) );
  OAI21X1 U1110 ( .A(n1246), .B(n1335), .C(n1475), .Y(n2303) );
  NAND2X1 U1111 ( .A(\mem<25><9> ), .B(n1482), .Y(n1476) );
  OAI21X1 U1112 ( .A(n1246), .B(n1337), .C(n1476), .Y(n2302) );
  NAND2X1 U1113 ( .A(\mem<25><10> ), .B(n1482), .Y(n1477) );
  OAI21X1 U1114 ( .A(n1246), .B(n1339), .C(n1477), .Y(n2301) );
  NAND2X1 U1115 ( .A(\mem<25><11> ), .B(n1482), .Y(n1478) );
  OAI21X1 U1116 ( .A(n1246), .B(n1341), .C(n1478), .Y(n2300) );
  NAND2X1 U1117 ( .A(\mem<25><12> ), .B(n1482), .Y(n1479) );
  OAI21X1 U1118 ( .A(n1246), .B(n1343), .C(n1479), .Y(n2299) );
  NAND2X1 U1119 ( .A(\mem<25><13> ), .B(n1482), .Y(n1480) );
  OAI21X1 U1120 ( .A(n1246), .B(n1345), .C(n1480), .Y(n2298) );
  NAND2X1 U1121 ( .A(\mem<25><14> ), .B(n1482), .Y(n1481) );
  OAI21X1 U1122 ( .A(n1246), .B(n1347), .C(n1481), .Y(n2297) );
  NAND2X1 U1123 ( .A(\mem<25><15> ), .B(n1482), .Y(n1483) );
  OAI21X1 U1124 ( .A(n1246), .B(n1349), .C(n1483), .Y(n2296) );
  NOR3X1 U1125 ( .A(n1351), .B(n1353), .C(n1192), .Y(n1879) );
  NAND2X1 U1126 ( .A(\mem<24><0> ), .B(n1499), .Y(n1484) );
  OAI21X1 U1127 ( .A(n100), .B(n1318), .C(n1484), .Y(n2295) );
  NAND2X1 U1128 ( .A(\mem<24><1> ), .B(n1499), .Y(n1485) );
  OAI21X1 U1129 ( .A(n100), .B(n1321), .C(n1485), .Y(n2294) );
  NAND2X1 U1130 ( .A(\mem<24><2> ), .B(n1499), .Y(n1486) );
  OAI21X1 U1131 ( .A(n100), .B(n1323), .C(n1486), .Y(n2293) );
  NAND2X1 U1132 ( .A(\mem<24><3> ), .B(n1499), .Y(n1487) );
  OAI21X1 U1133 ( .A(n100), .B(n1325), .C(n1487), .Y(n2292) );
  NAND2X1 U1134 ( .A(\mem<24><4> ), .B(n1499), .Y(n1488) );
  OAI21X1 U1135 ( .A(n100), .B(n1327), .C(n1488), .Y(n2291) );
  NAND2X1 U1136 ( .A(\mem<24><5> ), .B(n1499), .Y(n1489) );
  OAI21X1 U1137 ( .A(n100), .B(n1329), .C(n1489), .Y(n2290) );
  NAND2X1 U1138 ( .A(\mem<24><6> ), .B(n1499), .Y(n1490) );
  OAI21X1 U1139 ( .A(n100), .B(n1331), .C(n1490), .Y(n2289) );
  NAND2X1 U1140 ( .A(\mem<24><7> ), .B(n1499), .Y(n1491) );
  OAI21X1 U1141 ( .A(n100), .B(n1333), .C(n1491), .Y(n2288) );
  NAND2X1 U1142 ( .A(\mem<24><8> ), .B(n1499), .Y(n1492) );
  OAI21X1 U1143 ( .A(n100), .B(n1335), .C(n1492), .Y(n2287) );
  NAND2X1 U1144 ( .A(\mem<24><9> ), .B(n1499), .Y(n1493) );
  OAI21X1 U1145 ( .A(n100), .B(n1337), .C(n1493), .Y(n2286) );
  NAND2X1 U1146 ( .A(\mem<24><10> ), .B(n1499), .Y(n1494) );
  OAI21X1 U1147 ( .A(n100), .B(n1339), .C(n1494), .Y(n2285) );
  NAND2X1 U1148 ( .A(\mem<24><11> ), .B(n1499), .Y(n1495) );
  OAI21X1 U1149 ( .A(n100), .B(n1341), .C(n1495), .Y(n2284) );
  NAND2X1 U1150 ( .A(\mem<24><12> ), .B(n1499), .Y(n1496) );
  OAI21X1 U1151 ( .A(n100), .B(n1343), .C(n1496), .Y(n2283) );
  NAND2X1 U1152 ( .A(\mem<24><13> ), .B(n1499), .Y(n1497) );
  OAI21X1 U1153 ( .A(n100), .B(n1345), .C(n1497), .Y(n2282) );
  NAND2X1 U1154 ( .A(\mem<24><14> ), .B(n1499), .Y(n1498) );
  OAI21X1 U1155 ( .A(n100), .B(n1347), .C(n1498), .Y(n2281) );
  NAND2X1 U1156 ( .A(\mem<24><15> ), .B(n1499), .Y(n1500) );
  OAI21X1 U1157 ( .A(n100), .B(n1349), .C(n1500), .Y(n2280) );
  NAND2X1 U1158 ( .A(\mem<23><0> ), .B(n1516), .Y(n1501) );
  OAI21X1 U1159 ( .A(n1247), .B(n1318), .C(n1501), .Y(n2279) );
  NAND2X1 U1160 ( .A(\mem<23><1> ), .B(n1516), .Y(n1502) );
  OAI21X1 U1161 ( .A(n1247), .B(n1321), .C(n1502), .Y(n2278) );
  NAND2X1 U1162 ( .A(\mem<23><2> ), .B(n1516), .Y(n1503) );
  OAI21X1 U1163 ( .A(n1247), .B(n1323), .C(n1503), .Y(n2277) );
  NAND2X1 U1164 ( .A(\mem<23><3> ), .B(n1516), .Y(n1504) );
  OAI21X1 U1165 ( .A(n1247), .B(n1325), .C(n1504), .Y(n2276) );
  NAND2X1 U1166 ( .A(\mem<23><4> ), .B(n1516), .Y(n1505) );
  OAI21X1 U1167 ( .A(n1247), .B(n1327), .C(n1505), .Y(n2275) );
  NAND2X1 U1168 ( .A(\mem<23><5> ), .B(n1516), .Y(n1506) );
  OAI21X1 U1169 ( .A(n1247), .B(n1329), .C(n1506), .Y(n2274) );
  NAND2X1 U1170 ( .A(\mem<23><6> ), .B(n1516), .Y(n1507) );
  OAI21X1 U1171 ( .A(n1247), .B(n1331), .C(n1507), .Y(n2273) );
  NAND2X1 U1172 ( .A(\mem<23><7> ), .B(n1516), .Y(n1508) );
  OAI21X1 U1173 ( .A(n1247), .B(n1333), .C(n1508), .Y(n2272) );
  NAND2X1 U1174 ( .A(\mem<23><8> ), .B(n1516), .Y(n1509) );
  OAI21X1 U1175 ( .A(n1248), .B(n1335), .C(n1509), .Y(n2271) );
  NAND2X1 U1177 ( .A(\mem<23><9> ), .B(n1516), .Y(n1510) );
  OAI21X1 U1178 ( .A(n1248), .B(n1337), .C(n1510), .Y(n2270) );
  NAND2X1 U1179 ( .A(\mem<23><10> ), .B(n1516), .Y(n1511) );
  OAI21X1 U1180 ( .A(n1248), .B(n1339), .C(n1511), .Y(n2269) );
  NAND2X1 U1181 ( .A(\mem<23><11> ), .B(n1516), .Y(n1512) );
  OAI21X1 U1182 ( .A(n1248), .B(n1341), .C(n1512), .Y(n2268) );
  NAND2X1 U1183 ( .A(\mem<23><12> ), .B(n1516), .Y(n1513) );
  OAI21X1 U1184 ( .A(n1248), .B(n1343), .C(n1513), .Y(n2267) );
  NAND2X1 U1185 ( .A(\mem<23><13> ), .B(n1516), .Y(n1514) );
  OAI21X1 U1186 ( .A(n1248), .B(n1345), .C(n1514), .Y(n2266) );
  NAND2X1 U1187 ( .A(\mem<23><14> ), .B(n1516), .Y(n1515) );
  OAI21X1 U1188 ( .A(n1248), .B(n1347), .C(n1515), .Y(n2265) );
  NAND2X1 U1189 ( .A(\mem<23><15> ), .B(n1516), .Y(n1517) );
  OAI21X1 U1190 ( .A(n1248), .B(n1349), .C(n1517), .Y(n2264) );
  NAND2X1 U1191 ( .A(\mem<22><0> ), .B(n1251), .Y(n1518) );
  OAI21X1 U1192 ( .A(n1249), .B(n1318), .C(n1518), .Y(n2263) );
  NAND2X1 U1193 ( .A(\mem<22><1> ), .B(n1251), .Y(n1519) );
  OAI21X1 U1194 ( .A(n1249), .B(n1321), .C(n1519), .Y(n2262) );
  NAND2X1 U1195 ( .A(\mem<22><2> ), .B(n1251), .Y(n1520) );
  OAI21X1 U1196 ( .A(n1249), .B(n1323), .C(n1520), .Y(n2261) );
  NAND2X1 U1197 ( .A(\mem<22><3> ), .B(n1251), .Y(n1521) );
  OAI21X1 U1198 ( .A(n1249), .B(n1325), .C(n1521), .Y(n2260) );
  NAND2X1 U1199 ( .A(\mem<22><4> ), .B(n1251), .Y(n1522) );
  OAI21X1 U1200 ( .A(n1249), .B(n1327), .C(n1522), .Y(n2259) );
  NAND2X1 U1201 ( .A(\mem<22><5> ), .B(n1251), .Y(n1523) );
  OAI21X1 U1202 ( .A(n1249), .B(n1329), .C(n1523), .Y(n2258) );
  NAND2X1 U1203 ( .A(\mem<22><6> ), .B(n1251), .Y(n1524) );
  OAI21X1 U1204 ( .A(n1249), .B(n1331), .C(n1524), .Y(n2257) );
  NAND2X1 U1205 ( .A(\mem<22><7> ), .B(n1251), .Y(n1525) );
  OAI21X1 U1206 ( .A(n1249), .B(n1333), .C(n1525), .Y(n2256) );
  NAND2X1 U1207 ( .A(\mem<22><8> ), .B(n1252), .Y(n1526) );
  OAI21X1 U1208 ( .A(n1250), .B(n1335), .C(n1526), .Y(n2255) );
  NAND2X1 U1209 ( .A(\mem<22><9> ), .B(n1252), .Y(n1527) );
  OAI21X1 U1210 ( .A(n1250), .B(n1337), .C(n1527), .Y(n2254) );
  NAND2X1 U1211 ( .A(\mem<22><10> ), .B(n1252), .Y(n1528) );
  OAI21X1 U1212 ( .A(n1250), .B(n1339), .C(n1528), .Y(n2253) );
  NAND2X1 U1213 ( .A(\mem<22><11> ), .B(n1252), .Y(n1529) );
  OAI21X1 U1214 ( .A(n1250), .B(n1341), .C(n1529), .Y(n2252) );
  NAND2X1 U1215 ( .A(\mem<22><12> ), .B(n1252), .Y(n1530) );
  OAI21X1 U1216 ( .A(n1250), .B(n1343), .C(n1530), .Y(n2251) );
  NAND2X1 U1217 ( .A(\mem<22><13> ), .B(n1252), .Y(n1531) );
  OAI21X1 U1218 ( .A(n1250), .B(n1345), .C(n1531), .Y(n2250) );
  NAND2X1 U1219 ( .A(\mem<22><14> ), .B(n1252), .Y(n1532) );
  OAI21X1 U1220 ( .A(n1250), .B(n1347), .C(n1532), .Y(n2249) );
  NAND2X1 U1221 ( .A(\mem<22><15> ), .B(n1252), .Y(n1533) );
  OAI21X1 U1222 ( .A(n1250), .B(n1349), .C(n1533), .Y(n2248) );
  NAND2X1 U1223 ( .A(\mem<21><0> ), .B(n1255), .Y(n1534) );
  OAI21X1 U1224 ( .A(n1253), .B(n1318), .C(n1534), .Y(n2247) );
  NAND2X1 U1225 ( .A(\mem<21><1> ), .B(n1255), .Y(n1535) );
  OAI21X1 U1226 ( .A(n1253), .B(n1321), .C(n1535), .Y(n2246) );
  NAND2X1 U1227 ( .A(\mem<21><2> ), .B(n1255), .Y(n1536) );
  OAI21X1 U1228 ( .A(n1253), .B(n1323), .C(n1536), .Y(n2245) );
  NAND2X1 U1229 ( .A(\mem<21><3> ), .B(n1255), .Y(n1537) );
  OAI21X1 U1230 ( .A(n1253), .B(n1325), .C(n1537), .Y(n2244) );
  NAND2X1 U1231 ( .A(\mem<21><4> ), .B(n1255), .Y(n1538) );
  OAI21X1 U1232 ( .A(n1253), .B(n1327), .C(n1538), .Y(n2243) );
  NAND2X1 U1233 ( .A(\mem<21><5> ), .B(n1255), .Y(n1539) );
  OAI21X1 U1234 ( .A(n1253), .B(n1329), .C(n1539), .Y(n2242) );
  NAND2X1 U1235 ( .A(\mem<21><6> ), .B(n1255), .Y(n1540) );
  OAI21X1 U1236 ( .A(n1253), .B(n1331), .C(n1540), .Y(n2241) );
  NAND2X1 U1237 ( .A(\mem<21><7> ), .B(n1255), .Y(n1541) );
  OAI21X1 U1238 ( .A(n1253), .B(n1333), .C(n1541), .Y(n2240) );
  NAND2X1 U1239 ( .A(\mem<21><8> ), .B(n1256), .Y(n1542) );
  OAI21X1 U1240 ( .A(n1254), .B(n1335), .C(n1542), .Y(n2239) );
  NAND2X1 U1241 ( .A(\mem<21><9> ), .B(n1256), .Y(n1543) );
  OAI21X1 U1242 ( .A(n1254), .B(n1337), .C(n1543), .Y(n2238) );
  NAND2X1 U1243 ( .A(\mem<21><10> ), .B(n1256), .Y(n1544) );
  OAI21X1 U1244 ( .A(n1254), .B(n1339), .C(n1544), .Y(n2237) );
  NAND2X1 U1245 ( .A(\mem<21><11> ), .B(n1256), .Y(n1545) );
  OAI21X1 U1246 ( .A(n1254), .B(n1341), .C(n1545), .Y(n2236) );
  NAND2X1 U1247 ( .A(\mem<21><12> ), .B(n1256), .Y(n1546) );
  OAI21X1 U1248 ( .A(n1254), .B(n1343), .C(n1546), .Y(n2235) );
  NAND2X1 U1249 ( .A(\mem<21><13> ), .B(n1256), .Y(n1547) );
  OAI21X1 U1250 ( .A(n1254), .B(n1345), .C(n1547), .Y(n2234) );
  NAND2X1 U1251 ( .A(\mem<21><14> ), .B(n1256), .Y(n1548) );
  OAI21X1 U1252 ( .A(n1254), .B(n1347), .C(n1548), .Y(n2233) );
  NAND2X1 U1253 ( .A(\mem<21><15> ), .B(n1256), .Y(n1549) );
  OAI21X1 U1254 ( .A(n1254), .B(n1349), .C(n1549), .Y(n2232) );
  NAND2X1 U1255 ( .A(\mem<20><0> ), .B(n1259), .Y(n1550) );
  OAI21X1 U1256 ( .A(n1257), .B(n1318), .C(n1550), .Y(n2231) );
  NAND2X1 U1257 ( .A(\mem<20><1> ), .B(n1259), .Y(n1551) );
  OAI21X1 U1258 ( .A(n1257), .B(n1321), .C(n1551), .Y(n2230) );
  NAND2X1 U1259 ( .A(\mem<20><2> ), .B(n1259), .Y(n1552) );
  OAI21X1 U1260 ( .A(n1257), .B(n1323), .C(n1552), .Y(n2229) );
  NAND2X1 U1261 ( .A(\mem<20><3> ), .B(n1259), .Y(n1553) );
  OAI21X1 U1262 ( .A(n1257), .B(n1325), .C(n1553), .Y(n2228) );
  NAND2X1 U1263 ( .A(\mem<20><4> ), .B(n1259), .Y(n1554) );
  OAI21X1 U1264 ( .A(n1257), .B(n1327), .C(n1554), .Y(n2227) );
  NAND2X1 U1265 ( .A(\mem<20><5> ), .B(n1259), .Y(n1555) );
  OAI21X1 U1266 ( .A(n1257), .B(n1329), .C(n1555), .Y(n2226) );
  NAND2X1 U1267 ( .A(\mem<20><6> ), .B(n1259), .Y(n1556) );
  OAI21X1 U1268 ( .A(n1257), .B(n1331), .C(n1556), .Y(n2225) );
  NAND2X1 U1269 ( .A(\mem<20><7> ), .B(n1259), .Y(n1557) );
  OAI21X1 U1270 ( .A(n1257), .B(n1333), .C(n1557), .Y(n2224) );
  NAND2X1 U1271 ( .A(\mem<20><8> ), .B(n1260), .Y(n1558) );
  OAI21X1 U1272 ( .A(n1258), .B(n1335), .C(n1558), .Y(n2223) );
  NAND2X1 U1273 ( .A(\mem<20><9> ), .B(n1260), .Y(n1559) );
  OAI21X1 U1274 ( .A(n1258), .B(n1337), .C(n1559), .Y(n2222) );
  NAND2X1 U1275 ( .A(\mem<20><10> ), .B(n1260), .Y(n1560) );
  OAI21X1 U1276 ( .A(n1258), .B(n1339), .C(n1560), .Y(n2221) );
  NAND2X1 U1277 ( .A(\mem<20><11> ), .B(n1260), .Y(n1561) );
  OAI21X1 U1278 ( .A(n1258), .B(n1341), .C(n1561), .Y(n2220) );
  NAND2X1 U1279 ( .A(\mem<20><12> ), .B(n1260), .Y(n1562) );
  OAI21X1 U1280 ( .A(n1258), .B(n1343), .C(n1562), .Y(n2219) );
  NAND2X1 U1281 ( .A(\mem<20><13> ), .B(n1260), .Y(n1563) );
  OAI21X1 U1282 ( .A(n1258), .B(n1345), .C(n1563), .Y(n2218) );
  NAND2X1 U1283 ( .A(\mem<20><14> ), .B(n1260), .Y(n1564) );
  OAI21X1 U1284 ( .A(n1258), .B(n1347), .C(n1564), .Y(n2217) );
  NAND2X1 U1285 ( .A(\mem<20><15> ), .B(n1260), .Y(n1565) );
  OAI21X1 U1286 ( .A(n1258), .B(n1349), .C(n1565), .Y(n2216) );
  NAND2X1 U1287 ( .A(\mem<19><0> ), .B(n128), .Y(n1566) );
  OAI21X1 U1288 ( .A(n1261), .B(n1318), .C(n1566), .Y(n2215) );
  NAND2X1 U1289 ( .A(\mem<19><1> ), .B(n128), .Y(n1567) );
  OAI21X1 U1290 ( .A(n1261), .B(n1320), .C(n1567), .Y(n2214) );
  NAND2X1 U1291 ( .A(\mem<19><2> ), .B(n128), .Y(n1568) );
  OAI21X1 U1292 ( .A(n1261), .B(n1322), .C(n1568), .Y(n2213) );
  NAND2X1 U1293 ( .A(\mem<19><3> ), .B(n128), .Y(n1569) );
  OAI21X1 U1294 ( .A(n1261), .B(n1324), .C(n1569), .Y(n2212) );
  NAND2X1 U1295 ( .A(\mem<19><4> ), .B(n128), .Y(n1570) );
  OAI21X1 U1296 ( .A(n1261), .B(n1326), .C(n1570), .Y(n2211) );
  NAND2X1 U1297 ( .A(\mem<19><5> ), .B(n128), .Y(n1571) );
  OAI21X1 U1298 ( .A(n1261), .B(n1328), .C(n1571), .Y(n2210) );
  NAND2X1 U1299 ( .A(\mem<19><6> ), .B(n128), .Y(n1572) );
  OAI21X1 U1300 ( .A(n1261), .B(n1330), .C(n1572), .Y(n2209) );
  NAND2X1 U1301 ( .A(\mem<19><7> ), .B(n128), .Y(n1573) );
  OAI21X1 U1302 ( .A(n1261), .B(n1332), .C(n1573), .Y(n2208) );
  NAND2X1 U1303 ( .A(\mem<19><8> ), .B(n128), .Y(n1574) );
  OAI21X1 U1304 ( .A(n1262), .B(n1335), .C(n1574), .Y(n2207) );
  NAND2X1 U1305 ( .A(\mem<19><9> ), .B(n128), .Y(n1575) );
  OAI21X1 U1306 ( .A(n1262), .B(n1337), .C(n1575), .Y(n2206) );
  NAND2X1 U1307 ( .A(\mem<19><10> ), .B(n128), .Y(n1576) );
  OAI21X1 U1308 ( .A(n1262), .B(n1339), .C(n1576), .Y(n2205) );
  NAND2X1 U1309 ( .A(\mem<19><11> ), .B(n128), .Y(n1577) );
  OAI21X1 U1310 ( .A(n1262), .B(n1341), .C(n1577), .Y(n2204) );
  NAND2X1 U1311 ( .A(\mem<19><12> ), .B(n128), .Y(n1578) );
  OAI21X1 U1312 ( .A(n1262), .B(n1343), .C(n1578), .Y(n2203) );
  NAND2X1 U1313 ( .A(\mem<19><13> ), .B(n128), .Y(n1579) );
  OAI21X1 U1314 ( .A(n1262), .B(n1345), .C(n1579), .Y(n2202) );
  NAND2X1 U1315 ( .A(\mem<19><14> ), .B(n128), .Y(n1580) );
  OAI21X1 U1316 ( .A(n1262), .B(n1347), .C(n1580), .Y(n2201) );
  NAND2X1 U1317 ( .A(\mem<19><15> ), .B(n128), .Y(n1581) );
  OAI21X1 U1318 ( .A(n1262), .B(n1349), .C(n1581), .Y(n2200) );
  NAND2X1 U1319 ( .A(\mem<18><0> ), .B(n131), .Y(n1582) );
  OAI21X1 U1320 ( .A(n1263), .B(n1319), .C(n1582), .Y(n2199) );
  NAND2X1 U1321 ( .A(\mem<18><1> ), .B(n131), .Y(n1583) );
  OAI21X1 U1322 ( .A(n1263), .B(n1321), .C(n1583), .Y(n2198) );
  NAND2X1 U1323 ( .A(\mem<18><2> ), .B(n131), .Y(n1584) );
  OAI21X1 U1324 ( .A(n1263), .B(n1323), .C(n1584), .Y(n2197) );
  NAND2X1 U1325 ( .A(\mem<18><3> ), .B(n131), .Y(n1585) );
  OAI21X1 U1326 ( .A(n1263), .B(n1325), .C(n1585), .Y(n2196) );
  NAND2X1 U1327 ( .A(\mem<18><4> ), .B(n131), .Y(n1586) );
  OAI21X1 U1328 ( .A(n1263), .B(n1327), .C(n1586), .Y(n2195) );
  NAND2X1 U1329 ( .A(\mem<18><5> ), .B(n131), .Y(n1587) );
  OAI21X1 U1330 ( .A(n1263), .B(n1329), .C(n1587), .Y(n2194) );
  NAND2X1 U1331 ( .A(\mem<18><6> ), .B(n131), .Y(n1588) );
  OAI21X1 U1332 ( .A(n1263), .B(n1331), .C(n1588), .Y(n2193) );
  NAND2X1 U1333 ( .A(\mem<18><7> ), .B(n131), .Y(n1589) );
  OAI21X1 U1334 ( .A(n1263), .B(n1333), .C(n1589), .Y(n2192) );
  NAND2X1 U1335 ( .A(\mem<18><8> ), .B(n131), .Y(n1590) );
  OAI21X1 U1336 ( .A(n1264), .B(n1334), .C(n1590), .Y(n2191) );
  NAND2X1 U1337 ( .A(\mem<18><9> ), .B(n131), .Y(n1591) );
  OAI21X1 U1338 ( .A(n1264), .B(n1336), .C(n1591), .Y(n2190) );
  NAND2X1 U1339 ( .A(\mem<18><10> ), .B(n131), .Y(n1592) );
  OAI21X1 U1340 ( .A(n1264), .B(n1338), .C(n1592), .Y(n2189) );
  NAND2X1 U1341 ( .A(\mem<18><11> ), .B(n131), .Y(n1593) );
  OAI21X1 U1342 ( .A(n1264), .B(n1340), .C(n1593), .Y(n2188) );
  NAND2X1 U1343 ( .A(\mem<18><12> ), .B(n131), .Y(n1594) );
  OAI21X1 U1344 ( .A(n1264), .B(n1342), .C(n1594), .Y(n2187) );
  NAND2X1 U1345 ( .A(\mem<18><13> ), .B(n131), .Y(n1595) );
  OAI21X1 U1346 ( .A(n1264), .B(n1344), .C(n1595), .Y(n2186) );
  NAND2X1 U1347 ( .A(\mem<18><14> ), .B(n131), .Y(n1596) );
  OAI21X1 U1348 ( .A(n1264), .B(n1346), .C(n1596), .Y(n2185) );
  NAND2X1 U1349 ( .A(\mem<18><15> ), .B(n131), .Y(n1597) );
  OAI21X1 U1350 ( .A(n1264), .B(n1348), .C(n1597), .Y(n2184) );
  NAND2X1 U1351 ( .A(\mem<17><0> ), .B(n134), .Y(n1598) );
  OAI21X1 U1352 ( .A(n1265), .B(n1318), .C(n1598), .Y(n2183) );
  NAND2X1 U1353 ( .A(\mem<17><1> ), .B(n134), .Y(n1599) );
  OAI21X1 U1354 ( .A(n1265), .B(n1320), .C(n1599), .Y(n2182) );
  NAND2X1 U1355 ( .A(\mem<17><2> ), .B(n134), .Y(n1600) );
  OAI21X1 U1356 ( .A(n1265), .B(n1322), .C(n1600), .Y(n2181) );
  NAND2X1 U1357 ( .A(\mem<17><3> ), .B(n134), .Y(n1601) );
  OAI21X1 U1358 ( .A(n1265), .B(n1324), .C(n1601), .Y(n2180) );
  NAND2X1 U1359 ( .A(\mem<17><4> ), .B(n134), .Y(n1602) );
  OAI21X1 U1360 ( .A(n1265), .B(n1326), .C(n1602), .Y(n2179) );
  NAND2X1 U1361 ( .A(\mem<17><5> ), .B(n134), .Y(n1603) );
  OAI21X1 U1362 ( .A(n1265), .B(n1328), .C(n1603), .Y(n2178) );
  NAND2X1 U1363 ( .A(\mem<17><6> ), .B(n134), .Y(n1604) );
  OAI21X1 U1364 ( .A(n1265), .B(n1330), .C(n1604), .Y(n2177) );
  NAND2X1 U1365 ( .A(\mem<17><7> ), .B(n134), .Y(n1605) );
  OAI21X1 U1366 ( .A(n1265), .B(n1332), .C(n1605), .Y(n2176) );
  NAND2X1 U1367 ( .A(\mem<17><8> ), .B(n134), .Y(n1606) );
  OAI21X1 U1368 ( .A(n1266), .B(n1335), .C(n1606), .Y(n2175) );
  NAND2X1 U1369 ( .A(\mem<17><9> ), .B(n134), .Y(n1607) );
  OAI21X1 U1370 ( .A(n1266), .B(n1337), .C(n1607), .Y(n2174) );
  NAND2X1 U1371 ( .A(\mem<17><10> ), .B(n134), .Y(n1608) );
  OAI21X1 U1372 ( .A(n1266), .B(n1339), .C(n1608), .Y(n2173) );
  NAND2X1 U1373 ( .A(\mem<17><11> ), .B(n134), .Y(n1609) );
  OAI21X1 U1374 ( .A(n1266), .B(n1341), .C(n1609), .Y(n2172) );
  NAND2X1 U1375 ( .A(\mem<17><12> ), .B(n134), .Y(n1610) );
  OAI21X1 U1376 ( .A(n1266), .B(n1343), .C(n1610), .Y(n2171) );
  NAND2X1 U1377 ( .A(\mem<17><13> ), .B(n134), .Y(n1611) );
  OAI21X1 U1378 ( .A(n1266), .B(n1345), .C(n1611), .Y(n2170) );
  NAND2X1 U1379 ( .A(\mem<17><14> ), .B(n134), .Y(n1612) );
  OAI21X1 U1380 ( .A(n1266), .B(n1347), .C(n1612), .Y(n2169) );
  NAND2X1 U1381 ( .A(\mem<17><15> ), .B(n134), .Y(n1613) );
  OAI21X1 U1382 ( .A(n1266), .B(n1349), .C(n1613), .Y(n2168) );
  NAND2X1 U1383 ( .A(\mem<16><0> ), .B(n135), .Y(n1614) );
  OAI21X1 U1384 ( .A(n1267), .B(n1319), .C(n1614), .Y(n2167) );
  NAND2X1 U1385 ( .A(\mem<16><1> ), .B(n135), .Y(n1615) );
  OAI21X1 U1386 ( .A(n1267), .B(n1321), .C(n1615), .Y(n2166) );
  NAND2X1 U1387 ( .A(\mem<16><2> ), .B(n135), .Y(n1616) );
  OAI21X1 U1388 ( .A(n1267), .B(n1323), .C(n1616), .Y(n2165) );
  NAND2X1 U1389 ( .A(\mem<16><3> ), .B(n135), .Y(n1617) );
  OAI21X1 U1390 ( .A(n1267), .B(n1325), .C(n1617), .Y(n2164) );
  NAND2X1 U1391 ( .A(\mem<16><4> ), .B(n135), .Y(n1618) );
  OAI21X1 U1392 ( .A(n1267), .B(n1327), .C(n1618), .Y(n2163) );
  NAND2X1 U1393 ( .A(\mem<16><5> ), .B(n135), .Y(n1619) );
  OAI21X1 U1394 ( .A(n1267), .B(n1329), .C(n1619), .Y(n2162) );
  NAND2X1 U1395 ( .A(\mem<16><6> ), .B(n135), .Y(n1620) );
  OAI21X1 U1396 ( .A(n1267), .B(n1331), .C(n1620), .Y(n2161) );
  NAND2X1 U1397 ( .A(\mem<16><7> ), .B(n135), .Y(n1621) );
  OAI21X1 U1398 ( .A(n1267), .B(n1333), .C(n1621), .Y(n2160) );
  NAND2X1 U1399 ( .A(\mem<16><8> ), .B(n135), .Y(n1622) );
  OAI21X1 U1400 ( .A(n1267), .B(n1334), .C(n1622), .Y(n2159) );
  NAND2X1 U1401 ( .A(\mem<16><9> ), .B(n135), .Y(n1623) );
  OAI21X1 U1402 ( .A(n1267), .B(n1336), .C(n1623), .Y(n2158) );
  NAND2X1 U1403 ( .A(\mem<16><10> ), .B(n135), .Y(n1624) );
  OAI21X1 U1404 ( .A(n1267), .B(n1338), .C(n1624), .Y(n2157) );
  NAND2X1 U1405 ( .A(\mem<16><11> ), .B(n135), .Y(n1625) );
  OAI21X1 U1406 ( .A(n1267), .B(n1340), .C(n1625), .Y(n2156) );
  NAND2X1 U1407 ( .A(\mem<16><12> ), .B(n135), .Y(n1626) );
  OAI21X1 U1408 ( .A(n1267), .B(n1342), .C(n1626), .Y(n2155) );
  NAND2X1 U1409 ( .A(\mem<16><13> ), .B(n135), .Y(n1627) );
  OAI21X1 U1410 ( .A(n1267), .B(n1344), .C(n1627), .Y(n2154) );
  NAND2X1 U1411 ( .A(\mem<16><14> ), .B(n135), .Y(n1628) );
  OAI21X1 U1412 ( .A(n1267), .B(n1346), .C(n1628), .Y(n2153) );
  NAND2X1 U1413 ( .A(\mem<16><15> ), .B(n135), .Y(n1629) );
  OAI21X1 U1414 ( .A(n1267), .B(n1348), .C(n1629), .Y(n2152) );
  NAND3X1 U1415 ( .A(n1356), .B(n2408), .C(n1359), .Y(n1630) );
  NAND2X1 U1416 ( .A(\mem<15><0> ), .B(n138), .Y(n1631) );
  OAI21X1 U1417 ( .A(n1268), .B(n1319), .C(n1631), .Y(n2151) );
  NAND2X1 U1418 ( .A(\mem<15><1> ), .B(n138), .Y(n1632) );
  OAI21X1 U1419 ( .A(n1268), .B(n1321), .C(n1632), .Y(n2150) );
  NAND2X1 U1420 ( .A(\mem<15><2> ), .B(n138), .Y(n1633) );
  OAI21X1 U1421 ( .A(n1268), .B(n1323), .C(n1633), .Y(n2149) );
  NAND2X1 U1422 ( .A(\mem<15><3> ), .B(n138), .Y(n1634) );
  OAI21X1 U1423 ( .A(n1268), .B(n1325), .C(n1634), .Y(n2148) );
  NAND2X1 U1424 ( .A(\mem<15><4> ), .B(n138), .Y(n1635) );
  OAI21X1 U1425 ( .A(n1268), .B(n1327), .C(n1635), .Y(n2147) );
  NAND2X1 U1426 ( .A(\mem<15><5> ), .B(n138), .Y(n1636) );
  OAI21X1 U1427 ( .A(n1268), .B(n1329), .C(n1636), .Y(n2146) );
  NAND2X1 U1428 ( .A(\mem<15><6> ), .B(n138), .Y(n1637) );
  OAI21X1 U1429 ( .A(n1268), .B(n1331), .C(n1637), .Y(n2145) );
  NAND2X1 U1430 ( .A(\mem<15><7> ), .B(n138), .Y(n1638) );
  OAI21X1 U1431 ( .A(n1268), .B(n1333), .C(n1638), .Y(n2144) );
  NAND2X1 U1432 ( .A(\mem<15><8> ), .B(n138), .Y(n1639) );
  OAI21X1 U1433 ( .A(n1269), .B(n1334), .C(n1639), .Y(n2143) );
  NAND2X1 U1434 ( .A(\mem<15><9> ), .B(n138), .Y(n1640) );
  OAI21X1 U1435 ( .A(n1269), .B(n1336), .C(n1640), .Y(n2142) );
  NAND2X1 U1436 ( .A(\mem<15><10> ), .B(n138), .Y(n1641) );
  OAI21X1 U1437 ( .A(n1269), .B(n1338), .C(n1641), .Y(n2141) );
  NAND2X1 U1438 ( .A(\mem<15><11> ), .B(n138), .Y(n1642) );
  OAI21X1 U1439 ( .A(n1269), .B(n1340), .C(n1642), .Y(n2140) );
  NAND2X1 U1440 ( .A(\mem<15><12> ), .B(n138), .Y(n1643) );
  OAI21X1 U1441 ( .A(n1269), .B(n1342), .C(n1643), .Y(n2139) );
  NAND2X1 U1442 ( .A(\mem<15><13> ), .B(n138), .Y(n1644) );
  OAI21X1 U1443 ( .A(n1269), .B(n1344), .C(n1644), .Y(n2138) );
  NAND2X1 U1444 ( .A(\mem<15><14> ), .B(n138), .Y(n1645) );
  OAI21X1 U1445 ( .A(n1269), .B(n1346), .C(n1645), .Y(n2137) );
  NAND2X1 U1446 ( .A(\mem<15><15> ), .B(n138), .Y(n1646) );
  OAI21X1 U1447 ( .A(n1269), .B(n1348), .C(n1646), .Y(n2136) );
  NAND2X1 U1448 ( .A(\mem<14><0> ), .B(n1272), .Y(n1647) );
  OAI21X1 U1449 ( .A(n1270), .B(n1318), .C(n1647), .Y(n2135) );
  NAND2X1 U1450 ( .A(\mem<14><1> ), .B(n1272), .Y(n1648) );
  OAI21X1 U1451 ( .A(n1270), .B(n1320), .C(n1648), .Y(n2134) );
  NAND2X1 U1452 ( .A(\mem<14><2> ), .B(n1272), .Y(n1649) );
  OAI21X1 U1453 ( .A(n1270), .B(n1322), .C(n1649), .Y(n2133) );
  NAND2X1 U1454 ( .A(\mem<14><3> ), .B(n1272), .Y(n1650) );
  OAI21X1 U1455 ( .A(n1270), .B(n1324), .C(n1650), .Y(n2132) );
  NAND2X1 U1456 ( .A(\mem<14><4> ), .B(n1272), .Y(n1651) );
  OAI21X1 U1457 ( .A(n1270), .B(n1326), .C(n1651), .Y(n2131) );
  NAND2X1 U1458 ( .A(\mem<14><5> ), .B(n1272), .Y(n1652) );
  OAI21X1 U1459 ( .A(n1270), .B(n1328), .C(n1652), .Y(n2130) );
  NAND2X1 U1460 ( .A(\mem<14><6> ), .B(n1272), .Y(n1653) );
  OAI21X1 U1461 ( .A(n1270), .B(n1330), .C(n1653), .Y(n2129) );
  NAND2X1 U1462 ( .A(\mem<14><7> ), .B(n1272), .Y(n1654) );
  OAI21X1 U1463 ( .A(n1270), .B(n1332), .C(n1654), .Y(n2128) );
  NAND2X1 U1464 ( .A(\mem<14><8> ), .B(n1273), .Y(n1655) );
  OAI21X1 U1465 ( .A(n1271), .B(n1335), .C(n1655), .Y(n2127) );
  NAND2X1 U1466 ( .A(\mem<14><9> ), .B(n1273), .Y(n1656) );
  OAI21X1 U1467 ( .A(n1271), .B(n1337), .C(n1656), .Y(n2126) );
  NAND2X1 U1468 ( .A(\mem<14><10> ), .B(n1273), .Y(n1657) );
  OAI21X1 U1469 ( .A(n1271), .B(n1339), .C(n1657), .Y(n2125) );
  NAND2X1 U1470 ( .A(\mem<14><11> ), .B(n1273), .Y(n1658) );
  OAI21X1 U1471 ( .A(n1271), .B(n1341), .C(n1658), .Y(n2124) );
  NAND2X1 U1472 ( .A(\mem<14><12> ), .B(n1273), .Y(n1659) );
  OAI21X1 U1473 ( .A(n1271), .B(n1343), .C(n1659), .Y(n2123) );
  NAND2X1 U1474 ( .A(\mem<14><13> ), .B(n1273), .Y(n1660) );
  OAI21X1 U1475 ( .A(n1271), .B(n1345), .C(n1660), .Y(n2122) );
  NAND2X1 U1476 ( .A(\mem<14><14> ), .B(n1273), .Y(n1661) );
  OAI21X1 U1477 ( .A(n1271), .B(n1347), .C(n1661), .Y(n2121) );
  NAND2X1 U1478 ( .A(\mem<14><15> ), .B(n1273), .Y(n1662) );
  OAI21X1 U1479 ( .A(n1271), .B(n1349), .C(n1662), .Y(n2120) );
  NAND2X1 U1480 ( .A(\mem<13><0> ), .B(n1276), .Y(n1663) );
  OAI21X1 U1481 ( .A(n1274), .B(n1319), .C(n1663), .Y(n2119) );
  NAND2X1 U1482 ( .A(\mem<13><1> ), .B(n1276), .Y(n1664) );
  OAI21X1 U1483 ( .A(n1274), .B(n1321), .C(n1664), .Y(n2118) );
  NAND2X1 U1484 ( .A(\mem<13><2> ), .B(n1276), .Y(n1665) );
  OAI21X1 U1485 ( .A(n1274), .B(n1323), .C(n1665), .Y(n2117) );
  NAND2X1 U1486 ( .A(\mem<13><3> ), .B(n1276), .Y(n1666) );
  OAI21X1 U1487 ( .A(n1274), .B(n1325), .C(n1666), .Y(n2116) );
  NAND2X1 U1488 ( .A(\mem<13><4> ), .B(n1276), .Y(n1667) );
  OAI21X1 U1489 ( .A(n1274), .B(n1327), .C(n1667), .Y(n2115) );
  NAND2X1 U1490 ( .A(\mem<13><5> ), .B(n1276), .Y(n1668) );
  OAI21X1 U1491 ( .A(n1274), .B(n1329), .C(n1668), .Y(n2114) );
  NAND2X1 U1492 ( .A(\mem<13><6> ), .B(n1276), .Y(n1669) );
  OAI21X1 U1493 ( .A(n1274), .B(n1331), .C(n1669), .Y(n2113) );
  NAND2X1 U1494 ( .A(\mem<13><7> ), .B(n1276), .Y(n1670) );
  OAI21X1 U1495 ( .A(n1274), .B(n1333), .C(n1670), .Y(n2112) );
  NAND2X1 U1496 ( .A(\mem<13><8> ), .B(n1277), .Y(n1671) );
  OAI21X1 U1497 ( .A(n1275), .B(n1334), .C(n1671), .Y(n2111) );
  NAND2X1 U1498 ( .A(\mem<13><9> ), .B(n1277), .Y(n1672) );
  OAI21X1 U1499 ( .A(n1275), .B(n1336), .C(n1672), .Y(n2110) );
  NAND2X1 U1500 ( .A(\mem<13><10> ), .B(n1277), .Y(n1673) );
  OAI21X1 U1501 ( .A(n1275), .B(n1338), .C(n1673), .Y(n2109) );
  NAND2X1 U1502 ( .A(\mem<13><11> ), .B(n1277), .Y(n1674) );
  OAI21X1 U1503 ( .A(n1275), .B(n1340), .C(n1674), .Y(n2108) );
  NAND2X1 U1504 ( .A(\mem<13><12> ), .B(n1277), .Y(n1675) );
  OAI21X1 U1505 ( .A(n1275), .B(n1342), .C(n1675), .Y(n2107) );
  NAND2X1 U1506 ( .A(\mem<13><13> ), .B(n1277), .Y(n1676) );
  OAI21X1 U1507 ( .A(n1275), .B(n1344), .C(n1676), .Y(n2106) );
  NAND2X1 U1508 ( .A(\mem<13><14> ), .B(n1277), .Y(n1677) );
  OAI21X1 U1509 ( .A(n1275), .B(n1346), .C(n1677), .Y(n2105) );
  NAND2X1 U1510 ( .A(\mem<13><15> ), .B(n1277), .Y(n1678) );
  OAI21X1 U1511 ( .A(n1275), .B(n1348), .C(n1678), .Y(n2104) );
  NAND2X1 U1512 ( .A(\mem<12><0> ), .B(n1280), .Y(n1679) );
  OAI21X1 U1513 ( .A(n1278), .B(n1318), .C(n1679), .Y(n2103) );
  NAND2X1 U1514 ( .A(\mem<12><1> ), .B(n1280), .Y(n1680) );
  OAI21X1 U1515 ( .A(n1278), .B(n1320), .C(n1680), .Y(n2102) );
  NAND2X1 U1516 ( .A(\mem<12><2> ), .B(n1280), .Y(n1681) );
  OAI21X1 U1517 ( .A(n1278), .B(n1322), .C(n1681), .Y(n2101) );
  NAND2X1 U1518 ( .A(\mem<12><3> ), .B(n1280), .Y(n1682) );
  OAI21X1 U1519 ( .A(n1278), .B(n1324), .C(n1682), .Y(n2100) );
  NAND2X1 U1520 ( .A(\mem<12><4> ), .B(n1280), .Y(n1683) );
  OAI21X1 U1521 ( .A(n1278), .B(n1326), .C(n1683), .Y(n2099) );
  NAND2X1 U1522 ( .A(\mem<12><5> ), .B(n1280), .Y(n1684) );
  OAI21X1 U1523 ( .A(n1278), .B(n1328), .C(n1684), .Y(n2098) );
  NAND2X1 U1524 ( .A(\mem<12><6> ), .B(n1280), .Y(n1685) );
  OAI21X1 U1525 ( .A(n1278), .B(n1330), .C(n1685), .Y(n2097) );
  NAND2X1 U1526 ( .A(\mem<12><7> ), .B(n1280), .Y(n1686) );
  OAI21X1 U1527 ( .A(n1278), .B(n1332), .C(n1686), .Y(n2096) );
  NAND2X1 U1528 ( .A(\mem<12><8> ), .B(n1281), .Y(n1687) );
  OAI21X1 U1529 ( .A(n1279), .B(n1335), .C(n1687), .Y(n2095) );
  NAND2X1 U1530 ( .A(\mem<12><9> ), .B(n1281), .Y(n1688) );
  OAI21X1 U1531 ( .A(n1279), .B(n1337), .C(n1688), .Y(n2094) );
  NAND2X1 U1532 ( .A(\mem<12><10> ), .B(n1281), .Y(n1689) );
  OAI21X1 U1533 ( .A(n1279), .B(n1339), .C(n1689), .Y(n2093) );
  NAND2X1 U1534 ( .A(\mem<12><11> ), .B(n1281), .Y(n1690) );
  OAI21X1 U1535 ( .A(n1279), .B(n1341), .C(n1690), .Y(n2092) );
  NAND2X1 U1536 ( .A(\mem<12><12> ), .B(n1281), .Y(n1691) );
  OAI21X1 U1537 ( .A(n1279), .B(n1343), .C(n1691), .Y(n2091) );
  NAND2X1 U1538 ( .A(\mem<12><13> ), .B(n1281), .Y(n1692) );
  OAI21X1 U1539 ( .A(n1279), .B(n1345), .C(n1692), .Y(n2090) );
  NAND2X1 U1540 ( .A(\mem<12><14> ), .B(n1281), .Y(n1693) );
  OAI21X1 U1541 ( .A(n1279), .B(n1347), .C(n1693), .Y(n2089) );
  NAND2X1 U1542 ( .A(\mem<12><15> ), .B(n1281), .Y(n1694) );
  OAI21X1 U1543 ( .A(n1279), .B(n1349), .C(n1694), .Y(n2088) );
  NAND2X1 U1544 ( .A(\mem<11><0> ), .B(n1284), .Y(n1695) );
  OAI21X1 U1545 ( .A(n1282), .B(n1319), .C(n1695), .Y(n2087) );
  NAND2X1 U1546 ( .A(\mem<11><1> ), .B(n1284), .Y(n1696) );
  OAI21X1 U1547 ( .A(n1282), .B(n1320), .C(n1696), .Y(n2086) );
  NAND2X1 U1548 ( .A(\mem<11><2> ), .B(n1284), .Y(n1697) );
  OAI21X1 U1549 ( .A(n1282), .B(n1322), .C(n1697), .Y(n2085) );
  NAND2X1 U1550 ( .A(\mem<11><3> ), .B(n1284), .Y(n1698) );
  OAI21X1 U1551 ( .A(n1282), .B(n1324), .C(n1698), .Y(n2084) );
  NAND2X1 U1552 ( .A(\mem<11><4> ), .B(n1284), .Y(n1699) );
  OAI21X1 U1553 ( .A(n1282), .B(n1326), .C(n1699), .Y(n2083) );
  NAND2X1 U1554 ( .A(\mem<11><5> ), .B(n1284), .Y(n1700) );
  OAI21X1 U1555 ( .A(n1282), .B(n1328), .C(n1700), .Y(n2082) );
  NAND2X1 U1556 ( .A(\mem<11><6> ), .B(n1284), .Y(n1701) );
  OAI21X1 U1557 ( .A(n1282), .B(n1330), .C(n1701), .Y(n2081) );
  NAND2X1 U1558 ( .A(\mem<11><7> ), .B(n1284), .Y(n1702) );
  OAI21X1 U1559 ( .A(n1282), .B(n1332), .C(n1702), .Y(n2080) );
  NAND2X1 U1560 ( .A(\mem<11><8> ), .B(n1285), .Y(n1703) );
  OAI21X1 U1561 ( .A(n1283), .B(n1334), .C(n1703), .Y(n2079) );
  NAND2X1 U1562 ( .A(\mem<11><9> ), .B(n1285), .Y(n1704) );
  OAI21X1 U1563 ( .A(n1283), .B(n1336), .C(n1704), .Y(n2078) );
  NAND2X1 U1564 ( .A(\mem<11><10> ), .B(n1285), .Y(n1705) );
  OAI21X1 U1565 ( .A(n1283), .B(n1338), .C(n1705), .Y(n2077) );
  NAND2X1 U1566 ( .A(\mem<11><11> ), .B(n1285), .Y(n1706) );
  OAI21X1 U1567 ( .A(n1283), .B(n1340), .C(n1706), .Y(n2076) );
  NAND2X1 U1568 ( .A(\mem<11><12> ), .B(n1285), .Y(n1707) );
  OAI21X1 U1569 ( .A(n1283), .B(n1342), .C(n1707), .Y(n2075) );
  NAND2X1 U1570 ( .A(\mem<11><13> ), .B(n1285), .Y(n1708) );
  OAI21X1 U1571 ( .A(n1283), .B(n1344), .C(n1708), .Y(n2074) );
  NAND2X1 U1572 ( .A(\mem<11><14> ), .B(n1285), .Y(n1709) );
  OAI21X1 U1573 ( .A(n1283), .B(n1346), .C(n1709), .Y(n2073) );
  NAND2X1 U1574 ( .A(\mem<11><15> ), .B(n1285), .Y(n1710) );
  OAI21X1 U1575 ( .A(n1283), .B(n1348), .C(n1710), .Y(n2072) );
  NAND2X1 U1576 ( .A(\mem<10><0> ), .B(n1288), .Y(n1711) );
  OAI21X1 U1577 ( .A(n1286), .B(n1319), .C(n1711), .Y(n2071) );
  NAND2X1 U1578 ( .A(\mem<10><1> ), .B(n1288), .Y(n1712) );
  OAI21X1 U1579 ( .A(n1286), .B(n1320), .C(n1712), .Y(n2070) );
  NAND2X1 U1580 ( .A(\mem<10><2> ), .B(n1288), .Y(n1713) );
  OAI21X1 U1581 ( .A(n1286), .B(n1322), .C(n1713), .Y(n2069) );
  NAND2X1 U1582 ( .A(\mem<10><3> ), .B(n1288), .Y(n1714) );
  OAI21X1 U1583 ( .A(n1286), .B(n1324), .C(n1714), .Y(n2068) );
  NAND2X1 U1584 ( .A(\mem<10><4> ), .B(n1288), .Y(n1715) );
  OAI21X1 U1585 ( .A(n1286), .B(n1326), .C(n1715), .Y(n2067) );
  NAND2X1 U1586 ( .A(\mem<10><5> ), .B(n1288), .Y(n1716) );
  OAI21X1 U1587 ( .A(n1286), .B(n1328), .C(n1716), .Y(n2066) );
  NAND2X1 U1588 ( .A(\mem<10><6> ), .B(n1288), .Y(n1717) );
  OAI21X1 U1589 ( .A(n1286), .B(n1330), .C(n1717), .Y(n2065) );
  NAND2X1 U1590 ( .A(\mem<10><7> ), .B(n1288), .Y(n1718) );
  OAI21X1 U1591 ( .A(n1286), .B(n1332), .C(n1718), .Y(n2064) );
  NAND2X1 U1592 ( .A(\mem<10><8> ), .B(n1289), .Y(n1719) );
  OAI21X1 U1593 ( .A(n1287), .B(n1334), .C(n1719), .Y(n2063) );
  NAND2X1 U1594 ( .A(\mem<10><9> ), .B(n1289), .Y(n1720) );
  OAI21X1 U1595 ( .A(n1287), .B(n1336), .C(n1720), .Y(n2062) );
  NAND2X1 U1596 ( .A(\mem<10><10> ), .B(n1289), .Y(n1721) );
  OAI21X1 U1597 ( .A(n1287), .B(n1338), .C(n1721), .Y(n2061) );
  NAND2X1 U1598 ( .A(\mem<10><11> ), .B(n1289), .Y(n1722) );
  OAI21X1 U1599 ( .A(n1287), .B(n1340), .C(n1722), .Y(n2060) );
  NAND2X1 U1600 ( .A(\mem<10><12> ), .B(n1289), .Y(n1723) );
  OAI21X1 U1601 ( .A(n1287), .B(n1342), .C(n1723), .Y(n2059) );
  NAND2X1 U1602 ( .A(\mem<10><13> ), .B(n1289), .Y(n1724) );
  OAI21X1 U1603 ( .A(n1287), .B(n1344), .C(n1724), .Y(n2058) );
  NAND2X1 U1604 ( .A(\mem<10><14> ), .B(n1289), .Y(n1725) );
  OAI21X1 U1605 ( .A(n1287), .B(n1346), .C(n1725), .Y(n2057) );
  NAND2X1 U1606 ( .A(\mem<10><15> ), .B(n1289), .Y(n1726) );
  OAI21X1 U1607 ( .A(n1287), .B(n1348), .C(n1726), .Y(n2056) );
  NAND2X1 U1608 ( .A(\mem<9><0> ), .B(n1292), .Y(n1727) );
  OAI21X1 U1609 ( .A(n1290), .B(n1319), .C(n1727), .Y(n2055) );
  NAND2X1 U1610 ( .A(\mem<9><1> ), .B(n1292), .Y(n1728) );
  OAI21X1 U1611 ( .A(n1290), .B(n1320), .C(n1728), .Y(n2054) );
  NAND2X1 U1612 ( .A(\mem<9><2> ), .B(n1292), .Y(n1729) );
  OAI21X1 U1613 ( .A(n1290), .B(n1322), .C(n1729), .Y(n2053) );
  NAND2X1 U1614 ( .A(\mem<9><3> ), .B(n1292), .Y(n1730) );
  OAI21X1 U1615 ( .A(n1290), .B(n1324), .C(n1730), .Y(n2052) );
  NAND2X1 U1616 ( .A(\mem<9><4> ), .B(n1292), .Y(n1731) );
  OAI21X1 U1617 ( .A(n1290), .B(n1326), .C(n1731), .Y(n2051) );
  NAND2X1 U1618 ( .A(\mem<9><5> ), .B(n1292), .Y(n1732) );
  OAI21X1 U1619 ( .A(n1290), .B(n1328), .C(n1732), .Y(n2050) );
  NAND2X1 U1620 ( .A(\mem<9><6> ), .B(n1292), .Y(n1733) );
  OAI21X1 U1621 ( .A(n1290), .B(n1330), .C(n1733), .Y(n2049) );
  NAND2X1 U1622 ( .A(\mem<9><7> ), .B(n1292), .Y(n1734) );
  OAI21X1 U1623 ( .A(n1290), .B(n1332), .C(n1734), .Y(n2048) );
  NAND2X1 U1624 ( .A(\mem<9><8> ), .B(n1293), .Y(n1735) );
  OAI21X1 U1625 ( .A(n1291), .B(n1334), .C(n1735), .Y(n2047) );
  NAND2X1 U1626 ( .A(\mem<9><9> ), .B(n1293), .Y(n1736) );
  OAI21X1 U1627 ( .A(n1291), .B(n1336), .C(n1736), .Y(n2046) );
  NAND2X1 U1628 ( .A(\mem<9><10> ), .B(n1293), .Y(n1737) );
  OAI21X1 U1629 ( .A(n1291), .B(n1338), .C(n1737), .Y(n2045) );
  NAND2X1 U1630 ( .A(\mem<9><11> ), .B(n1293), .Y(n1738) );
  OAI21X1 U1631 ( .A(n1291), .B(n1340), .C(n1738), .Y(n2044) );
  NAND2X1 U1632 ( .A(\mem<9><12> ), .B(n1293), .Y(n1739) );
  OAI21X1 U1633 ( .A(n1291), .B(n1342), .C(n1739), .Y(n2043) );
  NAND2X1 U1634 ( .A(\mem<9><13> ), .B(n1293), .Y(n1740) );
  OAI21X1 U1635 ( .A(n1291), .B(n1344), .C(n1740), .Y(n2042) );
  NAND2X1 U1636 ( .A(\mem<9><14> ), .B(n1293), .Y(n1741) );
  OAI21X1 U1637 ( .A(n1291), .B(n1346), .C(n1741), .Y(n2041) );
  NAND2X1 U1638 ( .A(\mem<9><15> ), .B(n1293), .Y(n1742) );
  OAI21X1 U1639 ( .A(n1291), .B(n1348), .C(n1742), .Y(n2040) );
  NAND2X1 U1640 ( .A(\mem<8><0> ), .B(n1295), .Y(n1744) );
  OAI21X1 U1641 ( .A(n1294), .B(n1319), .C(n1744), .Y(n2039) );
  NAND2X1 U1642 ( .A(\mem<8><1> ), .B(n1295), .Y(n1745) );
  OAI21X1 U1643 ( .A(n1294), .B(n1320), .C(n1745), .Y(n2038) );
  NAND2X1 U1644 ( .A(\mem<8><2> ), .B(n1295), .Y(n1746) );
  OAI21X1 U1645 ( .A(n1294), .B(n1322), .C(n1746), .Y(n2037) );
  NAND2X1 U1646 ( .A(\mem<8><3> ), .B(n1295), .Y(n1747) );
  OAI21X1 U1647 ( .A(n1294), .B(n1324), .C(n1747), .Y(n2036) );
  NAND2X1 U1648 ( .A(\mem<8><4> ), .B(n1295), .Y(n1748) );
  OAI21X1 U1649 ( .A(n1294), .B(n1326), .C(n1748), .Y(n2035) );
  NAND2X1 U1650 ( .A(\mem<8><5> ), .B(n1295), .Y(n1749) );
  OAI21X1 U1651 ( .A(n1294), .B(n1328), .C(n1749), .Y(n2034) );
  NAND2X1 U1652 ( .A(\mem<8><6> ), .B(n1295), .Y(n1750) );
  OAI21X1 U1653 ( .A(n1294), .B(n1330), .C(n1750), .Y(n2033) );
  NAND2X1 U1654 ( .A(\mem<8><7> ), .B(n1295), .Y(n1751) );
  OAI21X1 U1655 ( .A(n1294), .B(n1332), .C(n1751), .Y(n2032) );
  NAND2X1 U1656 ( .A(\mem<8><8> ), .B(n1296), .Y(n1752) );
  OAI21X1 U1657 ( .A(n1294), .B(n1334), .C(n1752), .Y(n2031) );
  NAND2X1 U1658 ( .A(\mem<8><9> ), .B(n1296), .Y(n1753) );
  OAI21X1 U1659 ( .A(n1294), .B(n1336), .C(n1753), .Y(n2030) );
  NAND2X1 U1660 ( .A(\mem<8><10> ), .B(n1296), .Y(n1754) );
  OAI21X1 U1661 ( .A(n1294), .B(n1338), .C(n1754), .Y(n2029) );
  NAND2X1 U1662 ( .A(\mem<8><11> ), .B(n1296), .Y(n1755) );
  OAI21X1 U1663 ( .A(n1294), .B(n1340), .C(n1755), .Y(n2028) );
  NAND2X1 U1664 ( .A(\mem<8><12> ), .B(n1296), .Y(n1756) );
  OAI21X1 U1665 ( .A(n1294), .B(n1342), .C(n1756), .Y(n2027) );
  NAND2X1 U1666 ( .A(\mem<8><13> ), .B(n1296), .Y(n1757) );
  OAI21X1 U1667 ( .A(n1294), .B(n1344), .C(n1757), .Y(n2026) );
  NAND2X1 U1668 ( .A(\mem<8><14> ), .B(n1296), .Y(n1758) );
  OAI21X1 U1669 ( .A(n1294), .B(n1346), .C(n1758), .Y(n2025) );
  NAND2X1 U1670 ( .A(\mem<8><15> ), .B(n1296), .Y(n1759) );
  OAI21X1 U1671 ( .A(n1294), .B(n1348), .C(n1759), .Y(n2024) );
  NAND3X1 U1672 ( .A(n1357), .B(n2408), .C(n1359), .Y(n1760) );
  NAND2X1 U1673 ( .A(\mem<7><0> ), .B(n1299), .Y(n1761) );
  OAI21X1 U1674 ( .A(n1297), .B(n1319), .C(n1761), .Y(n2023) );
  NAND2X1 U1675 ( .A(\mem<7><1> ), .B(n1299), .Y(n1762) );
  OAI21X1 U1676 ( .A(n1297), .B(n1320), .C(n1762), .Y(n2022) );
  NAND2X1 U1677 ( .A(\mem<7><2> ), .B(n1299), .Y(n1763) );
  OAI21X1 U1678 ( .A(n1297), .B(n1322), .C(n1763), .Y(n2021) );
  NAND2X1 U1679 ( .A(\mem<7><3> ), .B(n1299), .Y(n1764) );
  OAI21X1 U1680 ( .A(n1297), .B(n1324), .C(n1764), .Y(n2020) );
  NAND2X1 U1681 ( .A(\mem<7><4> ), .B(n1299), .Y(n1765) );
  OAI21X1 U1682 ( .A(n1297), .B(n1326), .C(n1765), .Y(n2019) );
  NAND2X1 U1683 ( .A(\mem<7><5> ), .B(n1299), .Y(n1766) );
  OAI21X1 U1684 ( .A(n1297), .B(n1328), .C(n1766), .Y(n2018) );
  NAND2X1 U1685 ( .A(\mem<7><6> ), .B(n1299), .Y(n1767) );
  OAI21X1 U1686 ( .A(n1297), .B(n1330), .C(n1767), .Y(n2017) );
  NAND2X1 U1687 ( .A(\mem<7><7> ), .B(n1299), .Y(n1768) );
  OAI21X1 U1688 ( .A(n1297), .B(n1332), .C(n1768), .Y(n2016) );
  NAND2X1 U1689 ( .A(\mem<7><8> ), .B(n1300), .Y(n1769) );
  OAI21X1 U1690 ( .A(n1298), .B(n1334), .C(n1769), .Y(n2015) );
  NAND2X1 U1691 ( .A(\mem<7><9> ), .B(n1300), .Y(n1770) );
  OAI21X1 U1692 ( .A(n1298), .B(n1336), .C(n1770), .Y(n2014) );
  NAND2X1 U1693 ( .A(\mem<7><10> ), .B(n1300), .Y(n1771) );
  OAI21X1 U1694 ( .A(n1298), .B(n1338), .C(n1771), .Y(n2013) );
  NAND2X1 U1695 ( .A(\mem<7><11> ), .B(n1300), .Y(n1772) );
  OAI21X1 U1696 ( .A(n1298), .B(n1340), .C(n1772), .Y(n2012) );
  NAND2X1 U1697 ( .A(\mem<7><12> ), .B(n1300), .Y(n1773) );
  OAI21X1 U1698 ( .A(n1298), .B(n1342), .C(n1773), .Y(n2011) );
  NAND2X1 U1699 ( .A(\mem<7><13> ), .B(n1300), .Y(n1774) );
  OAI21X1 U1700 ( .A(n1298), .B(n1344), .C(n1774), .Y(n2010) );
  NAND2X1 U1701 ( .A(\mem<7><14> ), .B(n1300), .Y(n1775) );
  OAI21X1 U1702 ( .A(n1298), .B(n1346), .C(n1775), .Y(n2009) );
  NAND2X1 U1703 ( .A(\mem<7><15> ), .B(n1300), .Y(n1776) );
  OAI21X1 U1704 ( .A(n1298), .B(n1348), .C(n1776), .Y(n2008) );
  NAND2X1 U1705 ( .A(\mem<6><0> ), .B(n1303), .Y(n1777) );
  OAI21X1 U1706 ( .A(n1301), .B(n1319), .C(n1777), .Y(n2007) );
  NAND2X1 U1707 ( .A(\mem<6><1> ), .B(n1303), .Y(n1778) );
  OAI21X1 U1708 ( .A(n1301), .B(n1320), .C(n1778), .Y(n2006) );
  NAND2X1 U1709 ( .A(\mem<6><2> ), .B(n1303), .Y(n1779) );
  OAI21X1 U1710 ( .A(n1301), .B(n1322), .C(n1779), .Y(n2005) );
  NAND2X1 U1711 ( .A(\mem<6><3> ), .B(n1303), .Y(n1780) );
  OAI21X1 U1712 ( .A(n1301), .B(n1324), .C(n1780), .Y(n2004) );
  NAND2X1 U1713 ( .A(\mem<6><4> ), .B(n1303), .Y(n1781) );
  OAI21X1 U1714 ( .A(n1301), .B(n1326), .C(n1781), .Y(n2003) );
  NAND2X1 U1715 ( .A(\mem<6><5> ), .B(n1303), .Y(n1782) );
  OAI21X1 U1716 ( .A(n1301), .B(n1328), .C(n1782), .Y(n2002) );
  NAND2X1 U1717 ( .A(\mem<6><6> ), .B(n1303), .Y(n1783) );
  OAI21X1 U1718 ( .A(n1301), .B(n1330), .C(n1783), .Y(n2001) );
  NAND2X1 U1719 ( .A(\mem<6><7> ), .B(n1303), .Y(n1784) );
  OAI21X1 U1720 ( .A(n1301), .B(n1332), .C(n1784), .Y(n2000) );
  NAND2X1 U1721 ( .A(\mem<6><8> ), .B(n1304), .Y(n1785) );
  OAI21X1 U1722 ( .A(n1302), .B(n1334), .C(n1785), .Y(n1999) );
  NAND2X1 U1723 ( .A(\mem<6><9> ), .B(n1304), .Y(n1786) );
  OAI21X1 U1724 ( .A(n1302), .B(n1336), .C(n1786), .Y(n1998) );
  NAND2X1 U1725 ( .A(\mem<6><10> ), .B(n1304), .Y(n1787) );
  OAI21X1 U1726 ( .A(n1302), .B(n1338), .C(n1787), .Y(n1997) );
  NAND2X1 U1727 ( .A(\mem<6><11> ), .B(n1304), .Y(n1788) );
  OAI21X1 U1728 ( .A(n1302), .B(n1340), .C(n1788), .Y(n1996) );
  NAND2X1 U1729 ( .A(\mem<6><12> ), .B(n1304), .Y(n1789) );
  OAI21X1 U1730 ( .A(n1302), .B(n1342), .C(n1789), .Y(n1995) );
  NAND2X1 U1731 ( .A(\mem<6><13> ), .B(n1304), .Y(n1790) );
  OAI21X1 U1732 ( .A(n1302), .B(n1344), .C(n1790), .Y(n1994) );
  NAND2X1 U1733 ( .A(\mem<6><14> ), .B(n1304), .Y(n1791) );
  OAI21X1 U1734 ( .A(n1302), .B(n1346), .C(n1791), .Y(n1993) );
  NAND2X1 U1735 ( .A(\mem<6><15> ), .B(n1304), .Y(n1792) );
  OAI21X1 U1736 ( .A(n1302), .B(n1348), .C(n1792), .Y(n1992) );
  NAND2X1 U1737 ( .A(\mem<5><0> ), .B(n1307), .Y(n1794) );
  OAI21X1 U1738 ( .A(n1305), .B(n1319), .C(n1794), .Y(n1991) );
  NAND2X1 U1739 ( .A(\mem<5><1> ), .B(n1307), .Y(n1795) );
  OAI21X1 U1740 ( .A(n1305), .B(n1320), .C(n1795), .Y(n1990) );
  NAND2X1 U1741 ( .A(\mem<5><2> ), .B(n1307), .Y(n1796) );
  OAI21X1 U1742 ( .A(n1305), .B(n1322), .C(n1796), .Y(n1989) );
  NAND2X1 U1743 ( .A(\mem<5><3> ), .B(n1307), .Y(n1797) );
  OAI21X1 U1744 ( .A(n1305), .B(n1324), .C(n1797), .Y(n1988) );
  NAND2X1 U1745 ( .A(\mem<5><4> ), .B(n1307), .Y(n1798) );
  OAI21X1 U1746 ( .A(n1305), .B(n1326), .C(n1798), .Y(n1987) );
  NAND2X1 U1747 ( .A(\mem<5><5> ), .B(n1307), .Y(n1799) );
  OAI21X1 U1748 ( .A(n1305), .B(n1328), .C(n1799), .Y(n1986) );
  NAND2X1 U1749 ( .A(\mem<5><6> ), .B(n1307), .Y(n1800) );
  OAI21X1 U1750 ( .A(n1305), .B(n1330), .C(n1800), .Y(n1985) );
  NAND2X1 U1751 ( .A(\mem<5><7> ), .B(n1307), .Y(n1801) );
  OAI21X1 U1752 ( .A(n1305), .B(n1332), .C(n1801), .Y(n1984) );
  NAND2X1 U1753 ( .A(\mem<5><8> ), .B(n1308), .Y(n1802) );
  OAI21X1 U1754 ( .A(n1306), .B(n1334), .C(n1802), .Y(n1983) );
  NAND2X1 U1755 ( .A(\mem<5><9> ), .B(n1308), .Y(n1803) );
  OAI21X1 U1756 ( .A(n1306), .B(n1336), .C(n1803), .Y(n1982) );
  NAND2X1 U1757 ( .A(\mem<5><10> ), .B(n1308), .Y(n1804) );
  OAI21X1 U1758 ( .A(n1306), .B(n1338), .C(n1804), .Y(n1981) );
  NAND2X1 U1759 ( .A(\mem<5><11> ), .B(n1308), .Y(n1805) );
  OAI21X1 U1760 ( .A(n1306), .B(n1340), .C(n1805), .Y(n1980) );
  NAND2X1 U1761 ( .A(\mem<5><12> ), .B(n1308), .Y(n1806) );
  OAI21X1 U1762 ( .A(n1306), .B(n1342), .C(n1806), .Y(n1979) );
  NAND2X1 U1763 ( .A(\mem<5><13> ), .B(n1308), .Y(n1807) );
  OAI21X1 U1764 ( .A(n1306), .B(n1344), .C(n1807), .Y(n1978) );
  NAND2X1 U1765 ( .A(\mem<5><14> ), .B(n1308), .Y(n1808) );
  OAI21X1 U1766 ( .A(n1306), .B(n1346), .C(n1808), .Y(n1977) );
  NAND2X1 U1767 ( .A(\mem<5><15> ), .B(n1308), .Y(n1809) );
  OAI21X1 U1768 ( .A(n1306), .B(n1348), .C(n1809), .Y(n1976) );
  NAND2X1 U1769 ( .A(\mem<4><0> ), .B(n63), .Y(n1811) );
  OAI21X1 U1770 ( .A(n1309), .B(n1319), .C(n1811), .Y(n1975) );
  NAND2X1 U1771 ( .A(\mem<4><1> ), .B(n63), .Y(n1812) );
  OAI21X1 U1772 ( .A(n1309), .B(n1320), .C(n1812), .Y(n1974) );
  NAND2X1 U1773 ( .A(\mem<4><2> ), .B(n63), .Y(n1813) );
  OAI21X1 U1774 ( .A(n1309), .B(n1322), .C(n1813), .Y(n1973) );
  NAND2X1 U1775 ( .A(\mem<4><3> ), .B(n63), .Y(n1814) );
  OAI21X1 U1776 ( .A(n1309), .B(n1324), .C(n1814), .Y(n1972) );
  NAND2X1 U1777 ( .A(\mem<4><4> ), .B(n63), .Y(n1815) );
  OAI21X1 U1778 ( .A(n1309), .B(n1326), .C(n1815), .Y(n1971) );
  NAND2X1 U1779 ( .A(\mem<4><5> ), .B(n63), .Y(n1816) );
  OAI21X1 U1780 ( .A(n1309), .B(n1328), .C(n1816), .Y(n1970) );
  NAND2X1 U1781 ( .A(\mem<4><6> ), .B(n63), .Y(n1817) );
  OAI21X1 U1782 ( .A(n1309), .B(n1330), .C(n1817), .Y(n1969) );
  NAND2X1 U1783 ( .A(\mem<4><7> ), .B(n63), .Y(n1818) );
  OAI21X1 U1784 ( .A(n1309), .B(n1332), .C(n1818), .Y(n1968) );
  NAND2X1 U1785 ( .A(\mem<4><8> ), .B(n63), .Y(n1819) );
  OAI21X1 U1786 ( .A(n1310), .B(n1334), .C(n1819), .Y(n1967) );
  NAND2X1 U1787 ( .A(\mem<4><9> ), .B(n63), .Y(n1820) );
  OAI21X1 U1788 ( .A(n1310), .B(n1336), .C(n1820), .Y(n1966) );
  NAND2X1 U1789 ( .A(\mem<4><10> ), .B(n63), .Y(n1821) );
  OAI21X1 U1790 ( .A(n1310), .B(n1338), .C(n1821), .Y(n1965) );
  NAND2X1 U1791 ( .A(\mem<4><11> ), .B(n63), .Y(n1822) );
  OAI21X1 U1792 ( .A(n1310), .B(n1340), .C(n1822), .Y(n1964) );
  NAND2X1 U1793 ( .A(\mem<4><12> ), .B(n63), .Y(n1823) );
  OAI21X1 U1794 ( .A(n1310), .B(n1342), .C(n1823), .Y(n1963) );
  NAND2X1 U1795 ( .A(\mem<4><13> ), .B(n63), .Y(n1824) );
  OAI21X1 U1796 ( .A(n1310), .B(n1344), .C(n1824), .Y(n1962) );
  NAND2X1 U1797 ( .A(\mem<4><14> ), .B(n63), .Y(n1825) );
  OAI21X1 U1798 ( .A(n1310), .B(n1346), .C(n1825), .Y(n1961) );
  NAND2X1 U1799 ( .A(\mem<4><15> ), .B(n63), .Y(n1826) );
  OAI21X1 U1800 ( .A(n1310), .B(n1348), .C(n1826), .Y(n1960) );
  NAND2X1 U1801 ( .A(\mem<3><0> ), .B(n65), .Y(n1828) );
  OAI21X1 U1802 ( .A(n1311), .B(n1319), .C(n1828), .Y(n1959) );
  NAND2X1 U1803 ( .A(\mem<3><1> ), .B(n65), .Y(n1829) );
  OAI21X1 U1804 ( .A(n1311), .B(n1320), .C(n1829), .Y(n1958) );
  NAND2X1 U1805 ( .A(\mem<3><2> ), .B(n65), .Y(n1830) );
  OAI21X1 U1806 ( .A(n1311), .B(n1322), .C(n1830), .Y(n1957) );
  NAND2X1 U1807 ( .A(\mem<3><3> ), .B(n65), .Y(n1831) );
  OAI21X1 U1808 ( .A(n1311), .B(n1324), .C(n1831), .Y(n1956) );
  NAND2X1 U1809 ( .A(\mem<3><4> ), .B(n65), .Y(n1832) );
  OAI21X1 U1810 ( .A(n1311), .B(n1326), .C(n1832), .Y(n1955) );
  NAND2X1 U1811 ( .A(\mem<3><5> ), .B(n65), .Y(n1833) );
  OAI21X1 U1812 ( .A(n1311), .B(n1328), .C(n1833), .Y(n1954) );
  NAND2X1 U1813 ( .A(\mem<3><6> ), .B(n65), .Y(n1834) );
  OAI21X1 U1814 ( .A(n1311), .B(n1330), .C(n1834), .Y(n1953) );
  NAND2X1 U1815 ( .A(\mem<3><7> ), .B(n65), .Y(n1835) );
  OAI21X1 U1816 ( .A(n1311), .B(n1332), .C(n1835), .Y(n1952) );
  NAND2X1 U1817 ( .A(\mem<3><8> ), .B(n65), .Y(n1836) );
  OAI21X1 U1818 ( .A(n1312), .B(n1334), .C(n1836), .Y(n1951) );
  NAND2X1 U1819 ( .A(\mem<3><9> ), .B(n65), .Y(n1837) );
  OAI21X1 U1820 ( .A(n1312), .B(n1336), .C(n1837), .Y(n1950) );
  NAND2X1 U1821 ( .A(\mem<3><10> ), .B(n65), .Y(n1838) );
  OAI21X1 U1822 ( .A(n1312), .B(n1338), .C(n1838), .Y(n1949) );
  NAND2X1 U1823 ( .A(\mem<3><11> ), .B(n65), .Y(n1839) );
  OAI21X1 U1824 ( .A(n1312), .B(n1340), .C(n1839), .Y(n1948) );
  NAND2X1 U1825 ( .A(\mem<3><12> ), .B(n65), .Y(n1840) );
  OAI21X1 U1826 ( .A(n1312), .B(n1342), .C(n1840), .Y(n1947) );
  NAND2X1 U1827 ( .A(\mem<3><13> ), .B(n65), .Y(n1841) );
  OAI21X1 U1828 ( .A(n1312), .B(n1344), .C(n1841), .Y(n1946) );
  NAND2X1 U1829 ( .A(\mem<3><14> ), .B(n65), .Y(n1842) );
  OAI21X1 U1830 ( .A(n1312), .B(n1346), .C(n1842), .Y(n1945) );
  NAND2X1 U1831 ( .A(\mem<3><15> ), .B(n65), .Y(n1843) );
  OAI21X1 U1832 ( .A(n1312), .B(n1348), .C(n1843), .Y(n1944) );
  NAND2X1 U1833 ( .A(\mem<2><0> ), .B(n163), .Y(n1845) );
  OAI21X1 U1834 ( .A(n1313), .B(n1319), .C(n1845), .Y(n1943) );
  NAND2X1 U1835 ( .A(\mem<2><1> ), .B(n163), .Y(n1846) );
  OAI21X1 U1836 ( .A(n1313), .B(n1320), .C(n1846), .Y(n1942) );
  NAND2X1 U1837 ( .A(\mem<2><2> ), .B(n163), .Y(n1847) );
  OAI21X1 U1838 ( .A(n1313), .B(n1322), .C(n1847), .Y(n1941) );
  NAND2X1 U1839 ( .A(\mem<2><3> ), .B(n163), .Y(n1848) );
  OAI21X1 U1840 ( .A(n1313), .B(n1324), .C(n1848), .Y(n1940) );
  NAND2X1 U1841 ( .A(\mem<2><4> ), .B(n163), .Y(n1849) );
  OAI21X1 U1842 ( .A(n1313), .B(n1326), .C(n1849), .Y(n1939) );
  NAND2X1 U1843 ( .A(\mem<2><5> ), .B(n163), .Y(n1850) );
  OAI21X1 U1844 ( .A(n1313), .B(n1328), .C(n1850), .Y(n1938) );
  NAND2X1 U1845 ( .A(\mem<2><6> ), .B(n163), .Y(n1851) );
  OAI21X1 U1846 ( .A(n1313), .B(n1330), .C(n1851), .Y(n1937) );
  NAND2X1 U1847 ( .A(\mem<2><7> ), .B(n163), .Y(n1852) );
  OAI21X1 U1848 ( .A(n1313), .B(n1332), .C(n1852), .Y(n1936) );
  NAND2X1 U1849 ( .A(\mem<2><8> ), .B(n163), .Y(n1853) );
  OAI21X1 U1850 ( .A(n1314), .B(n1334), .C(n1853), .Y(n1935) );
  NAND2X1 U1851 ( .A(\mem<2><9> ), .B(n163), .Y(n1854) );
  OAI21X1 U1852 ( .A(n1314), .B(n1336), .C(n1854), .Y(n1934) );
  NAND2X1 U1853 ( .A(\mem<2><10> ), .B(n163), .Y(n1855) );
  OAI21X1 U1854 ( .A(n1314), .B(n1338), .C(n1855), .Y(n1933) );
  NAND2X1 U1855 ( .A(\mem<2><11> ), .B(n163), .Y(n1856) );
  OAI21X1 U1856 ( .A(n1314), .B(n1340), .C(n1856), .Y(n1932) );
  NAND2X1 U1857 ( .A(\mem<2><12> ), .B(n163), .Y(n1857) );
  OAI21X1 U1858 ( .A(n1314), .B(n1342), .C(n1857), .Y(n1931) );
  NAND2X1 U1859 ( .A(\mem<2><13> ), .B(n163), .Y(n1858) );
  OAI21X1 U1860 ( .A(n1314), .B(n1344), .C(n1858), .Y(n1930) );
  NAND2X1 U1861 ( .A(\mem<2><14> ), .B(n163), .Y(n1859) );
  OAI21X1 U1862 ( .A(n1314), .B(n1346), .C(n1859), .Y(n1929) );
  NAND2X1 U1863 ( .A(\mem<2><15> ), .B(n163), .Y(n1860) );
  OAI21X1 U1864 ( .A(n1314), .B(n1348), .C(n1860), .Y(n1928) );
  NAND2X1 U1865 ( .A(\mem<1><0> ), .B(n166), .Y(n1862) );
  OAI21X1 U1866 ( .A(n1315), .B(n1319), .C(n1862), .Y(n1927) );
  NAND2X1 U1867 ( .A(\mem<1><1> ), .B(n166), .Y(n1863) );
  OAI21X1 U1868 ( .A(n1315), .B(n1320), .C(n1863), .Y(n1926) );
  NAND2X1 U1869 ( .A(\mem<1><2> ), .B(n166), .Y(n1864) );
  OAI21X1 U1870 ( .A(n1315), .B(n1322), .C(n1864), .Y(n1925) );
  NAND2X1 U1871 ( .A(\mem<1><3> ), .B(n166), .Y(n1865) );
  OAI21X1 U1872 ( .A(n1315), .B(n1324), .C(n1865), .Y(n1924) );
  NAND2X1 U1873 ( .A(\mem<1><4> ), .B(n166), .Y(n1866) );
  OAI21X1 U1874 ( .A(n1315), .B(n1326), .C(n1866), .Y(n1923) );
  NAND2X1 U1875 ( .A(\mem<1><5> ), .B(n166), .Y(n1867) );
  OAI21X1 U1876 ( .A(n1315), .B(n1328), .C(n1867), .Y(n1922) );
  NAND2X1 U1877 ( .A(\mem<1><6> ), .B(n166), .Y(n1868) );
  OAI21X1 U1878 ( .A(n1315), .B(n1330), .C(n1868), .Y(n1921) );
  NAND2X1 U1879 ( .A(\mem<1><7> ), .B(n166), .Y(n1869) );
  OAI21X1 U1880 ( .A(n1315), .B(n1332), .C(n1869), .Y(n1920) );
  NAND2X1 U1881 ( .A(\mem<1><8> ), .B(n166), .Y(n1870) );
  OAI21X1 U1882 ( .A(n1316), .B(n1334), .C(n1870), .Y(n1919) );
  NAND2X1 U1883 ( .A(\mem<1><9> ), .B(n166), .Y(n1871) );
  OAI21X1 U1884 ( .A(n1316), .B(n1336), .C(n1871), .Y(n1918) );
  NAND2X1 U1885 ( .A(\mem<1><10> ), .B(n166), .Y(n1872) );
  OAI21X1 U1886 ( .A(n1316), .B(n1338), .C(n1872), .Y(n1917) );
  NAND2X1 U1887 ( .A(\mem<1><11> ), .B(n166), .Y(n1873) );
  OAI21X1 U1888 ( .A(n1316), .B(n1340), .C(n1873), .Y(n1916) );
  NAND2X1 U1889 ( .A(\mem<1><12> ), .B(n166), .Y(n1874) );
  OAI21X1 U1890 ( .A(n1316), .B(n1342), .C(n1874), .Y(n1915) );
  NAND2X1 U1891 ( .A(\mem<1><13> ), .B(n166), .Y(n1875) );
  OAI21X1 U1892 ( .A(n1316), .B(n1344), .C(n1875), .Y(n1914) );
  NAND2X1 U1893 ( .A(\mem<1><14> ), .B(n166), .Y(n1876) );
  OAI21X1 U1894 ( .A(n1316), .B(n1346), .C(n1876), .Y(n1913) );
  NAND2X1 U1895 ( .A(\mem<1><15> ), .B(n166), .Y(n1877) );
  OAI21X1 U1896 ( .A(n1316), .B(n1348), .C(n1877), .Y(n1912) );
  NAND2X1 U1897 ( .A(\mem<0><0> ), .B(n167), .Y(n1880) );
  OAI21X1 U1898 ( .A(n1317), .B(n1319), .C(n1880), .Y(n1911) );
  NAND2X1 U1899 ( .A(\mem<0><1> ), .B(n167), .Y(n1881) );
  OAI21X1 U1900 ( .A(n1317), .B(n1320), .C(n1881), .Y(n1910) );
  NAND2X1 U1901 ( .A(\mem<0><2> ), .B(n167), .Y(n1882) );
  OAI21X1 U1902 ( .A(n1317), .B(n1322), .C(n1882), .Y(n1909) );
  NAND2X1 U1903 ( .A(\mem<0><3> ), .B(n167), .Y(n1883) );
  OAI21X1 U1904 ( .A(n1317), .B(n1324), .C(n1883), .Y(n1908) );
  NAND2X1 U1905 ( .A(\mem<0><4> ), .B(n167), .Y(n1884) );
  OAI21X1 U1906 ( .A(n1317), .B(n1326), .C(n1884), .Y(n1907) );
  NAND2X1 U1907 ( .A(\mem<0><5> ), .B(n167), .Y(n1885) );
  OAI21X1 U1908 ( .A(n1317), .B(n1328), .C(n1885), .Y(n1906) );
  NAND2X1 U1909 ( .A(\mem<0><6> ), .B(n167), .Y(n1886) );
  OAI21X1 U1910 ( .A(n1317), .B(n1330), .C(n1886), .Y(n1905) );
  NAND2X1 U1911 ( .A(\mem<0><7> ), .B(n167), .Y(n1887) );
  OAI21X1 U1912 ( .A(n1317), .B(n1332), .C(n1887), .Y(n1904) );
  NAND2X1 U1913 ( .A(\mem<0><8> ), .B(n167), .Y(n1888) );
  OAI21X1 U1914 ( .A(n1317), .B(n1334), .C(n1888), .Y(n1903) );
  NAND2X1 U1915 ( .A(\mem<0><9> ), .B(n167), .Y(n1889) );
  OAI21X1 U1916 ( .A(n1317), .B(n1336), .C(n1889), .Y(n1902) );
  NAND2X1 U1917 ( .A(\mem<0><10> ), .B(n167), .Y(n1890) );
  OAI21X1 U1918 ( .A(n1317), .B(n1338), .C(n1890), .Y(n1901) );
  NAND2X1 U1919 ( .A(\mem<0><11> ), .B(n167), .Y(n1891) );
  OAI21X1 U1920 ( .A(n1317), .B(n1340), .C(n1891), .Y(n1900) );
  NAND2X1 U1921 ( .A(\mem<0><12> ), .B(n167), .Y(n1892) );
  OAI21X1 U1922 ( .A(n1317), .B(n1342), .C(n1892), .Y(n1899) );
  NAND2X1 U1923 ( .A(\mem<0><13> ), .B(n167), .Y(n1893) );
  OAI21X1 U1924 ( .A(n1317), .B(n1344), .C(n1893), .Y(n1898) );
  NAND2X1 U1925 ( .A(\mem<0><14> ), .B(n167), .Y(n1894) );
  OAI21X1 U1926 ( .A(n1317), .B(n1346), .C(n1894), .Y(n1897) );
  NAND2X1 U1927 ( .A(\mem<0><15> ), .B(n167), .Y(n1895) );
  OAI21X1 U1928 ( .A(n1317), .B(n1348), .C(n1895), .Y(n1896) );
endmodule


module memc_Size16_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1881), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1882), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1883), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1884), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1885), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1886), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1887), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1888), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1889), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1890), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1891), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1892), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1893), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1894), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1895), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1896), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1897), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1898), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1899), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1900), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1901), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1902), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1903), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1904), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1905), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1906), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1907), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1908), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1909), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1910), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1911), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1912), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1913), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1914), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1915), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1916), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1917), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1918), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1919), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1920), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1921), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1922), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1923), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1924), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1925), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1926), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1927), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1928), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1929), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1930), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1931), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1932), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1933), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1934), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1935), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1936), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1937), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1938), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1939), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1940), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1941), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1942), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1943), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1944), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1945), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1946), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1947), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1948), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1949), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1950), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1951), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1952), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1953), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1954), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1955), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1956), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1957), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1958), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1959), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1960), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1961), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1962), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1963), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1964), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1965), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1966), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1967), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1968), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1969), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1970), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1971), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1972), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1973), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1974), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1975), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1976), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1977), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1978), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1979), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1980), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1981), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1982), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1983), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1984), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1985), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1986), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1987), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1988), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1989), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1990), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1991), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1992), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1993), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1994), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1995), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1996), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1997), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1998), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1999), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2000), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2001), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2002), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2003), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2004), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2005), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2006), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2007), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2008), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2009), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2010), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2011), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2012), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2013), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2014), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2015), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2016), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2017), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2018), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2019), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2020), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2021), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2022), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2023), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2024), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2025), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2026), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2027), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2028), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2029), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2030), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2031), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2032), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2033), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2034), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2035), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2036), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2037), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2038), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2039), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2040), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2041), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2042), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2043), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2044), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2045), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2046), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2047), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2048), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2049), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2050), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2051), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2052), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2053), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2054), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2055), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2056), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2057), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2058), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2059), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2060), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2061), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2062), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2063), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2064), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2065), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2066), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2067), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2068), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2069), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2070), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2071), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2072), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2073), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2074), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2075), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2076), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2077), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2078), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2079), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2080), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2081), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2082), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2083), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2084), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2085), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2086), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2087), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2088), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2089), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2090), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2091), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2092), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2093), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2094), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2095), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2096), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2097), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2098), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2099), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2100), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2101), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2102), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2103), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2104), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2105), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2106), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2107), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2108), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2109), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2110), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2111), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2112), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2113), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2114), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2115), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2116), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2117), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2118), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2119), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2120), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2121), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2122), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2123), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2124), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2125), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2126), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2127), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2128), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2129), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2130), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2131), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2132), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2133), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2134), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2135), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2136), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2137), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2138), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2139), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2140), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2141), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2142), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2143), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2144), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2145), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2146), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2147), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2148), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2149), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2150), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2151), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2152), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2153), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2154), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2155), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2156), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2157), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2158), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2159), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2160), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2161), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2162), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2163), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2164), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2165), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2166), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2167), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2168), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2169), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2170), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2171), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2172), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2173), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2174), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2175), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2176), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2177), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2178), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2179), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2180), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2181), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2182), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2183), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2184), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2185), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2186), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2187), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2188), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2189), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2190), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2191), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2192), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2193), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2194), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2195), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2196), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2197), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2198), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2199), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2200), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2201), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2202), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2203), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2204), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2205), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2206), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2207), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2208), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2209), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2210), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2211), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2212), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2213), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2214), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2215), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2216), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2217), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2218), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2219), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2220), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2221), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2222), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2223), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2224), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2225), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2226), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2227), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2228), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2229), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2230), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2231), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2232), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2233), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2234), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2235), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2236), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2237), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2238), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2239), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2240), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2241), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2242), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2243), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2244), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2245), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2246), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2247), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2248), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2249), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2250), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2251), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2252), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2253), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2254), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2255), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2256), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2257), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2258), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2259), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2260), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2261), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2262), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2263), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2264), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2265), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2266), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2267), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2268), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2269), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2270), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2271), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2272), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2273), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2274), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2275), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2276), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2277), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2278), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2279), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2280), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2281), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2282), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2283), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2284), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2285), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2286), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2287), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2288), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2289), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2290), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2291), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2292), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2293), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2294), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2295), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2296), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2297), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2298), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2299), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2300), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2301), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2302), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2303), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2304), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2305), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2306), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2307), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2308), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2309), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2310), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2311), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2312), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2313), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2314), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2315), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2316), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2317), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2318), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2319), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2320), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2321), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2322), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2323), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2324), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2325), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2326), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2327), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2328), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2329), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2330), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2331), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2332), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2333), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2334), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2335), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2336), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2337), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2338), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2339), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2340), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2341), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2342), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2343), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2344), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2345), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2346), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2347), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2348), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2349), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2350), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2351), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2352), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2353), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2354), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2355), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2356), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2357), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2358), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2359), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2360), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2361), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2362), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2363), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2364), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2365), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2366), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2367), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2368), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2369), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2370), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2371), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2372), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2373), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2374), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2375), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2376), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2377), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2378), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2379), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2380), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2381), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2382), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2383), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2384), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2385), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2386), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2387), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2388), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2389), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2390), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2391), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2392), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2393) );
  INVX4 U2 ( .A(n66), .Y(n67) );
  INVX4 U3 ( .A(n64), .Y(n65) );
  INVX4 U4 ( .A(n62), .Y(n63) );
  INVX4 U5 ( .A(n60), .Y(n61) );
  INVX4 U6 ( .A(n58), .Y(n59) );
  INVX4 U7 ( .A(n56), .Y(n57) );
  INVX4 U8 ( .A(n91), .Y(n92) );
  INVX4 U9 ( .A(n89), .Y(n90) );
  INVX4 U10 ( .A(n87), .Y(n88) );
  INVX4 U11 ( .A(n85), .Y(n86) );
  INVX4 U12 ( .A(n83), .Y(n84) );
  INVX4 U13 ( .A(n78), .Y(n79) );
  INVX4 U14 ( .A(n76), .Y(n77) );
  INVX4 U15 ( .A(n74), .Y(n75) );
  INVX4 U16 ( .A(n42), .Y(n43) );
  INVX4 U17 ( .A(n40), .Y(n41) );
  INVX4 U18 ( .A(n39), .Y(n1) );
  INVX1 U19 ( .A(n1192), .Y(n1194) );
  INVX1 U20 ( .A(n1175), .Y(N31) );
  INVX1 U21 ( .A(n1178), .Y(N28) );
  INVX1 U22 ( .A(n1180), .Y(N26) );
  INVX1 U23 ( .A(n1181), .Y(N25) );
  INVX1 U24 ( .A(rst), .Y(n1344) );
  INVX1 U25 ( .A(n1187), .Y(N19) );
  INVX1 U26 ( .A(n1188), .Y(N18) );
  INVX1 U27 ( .A(n1236), .Y(n1211) );
  INVX1 U28 ( .A(n1347), .Y(n1197) );
  INVX1 U29 ( .A(n1213), .Y(n1215) );
  INVX1 U30 ( .A(n1213), .Y(n1214) );
  INVX1 U31 ( .A(n1198), .Y(n1199) );
  INVX1 U32 ( .A(n1213), .Y(n1216) );
  INVX1 U33 ( .A(n1212), .Y(n1217) );
  INVX1 U34 ( .A(n1198), .Y(n1200) );
  INVX1 U35 ( .A(n1212), .Y(n1219) );
  INVX1 U36 ( .A(n1212), .Y(n1218) );
  INVX1 U37 ( .A(n1198), .Y(n1201) );
  INVX1 U38 ( .A(n1212), .Y(n1220) );
  INVX1 U39 ( .A(n1213), .Y(n1221) );
  INVX1 U40 ( .A(n1197), .Y(n1202) );
  INVX2 U41 ( .A(n1213), .Y(n1222) );
  INVX1 U42 ( .A(n1211), .Y(n1223) );
  INVX1 U43 ( .A(n1197), .Y(n1203) );
  INVX1 U44 ( .A(n1211), .Y(n1224) );
  INVX1 U45 ( .A(n1211), .Y(n1225) );
  INVX1 U46 ( .A(n1197), .Y(n1204) );
  INVX1 U47 ( .A(n1211), .Y(n1226) );
  INVX1 U48 ( .A(n1211), .Y(n1227) );
  INVX2 U49 ( .A(n1197), .Y(n1205) );
  INVX1 U50 ( .A(n1212), .Y(n1228) );
  INVX1 U51 ( .A(n1211), .Y(n1229) );
  INVX1 U52 ( .A(n1197), .Y(n1206) );
  INVX1 U53 ( .A(n1211), .Y(n1231) );
  INVX1 U54 ( .A(n1211), .Y(n1230) );
  INVX1 U55 ( .A(n1197), .Y(n1207) );
  INVX1 U56 ( .A(n1210), .Y(n1232) );
  INVX1 U57 ( .A(n1210), .Y(n1233) );
  INVX2 U58 ( .A(n1198), .Y(n1208) );
  INVX1 U59 ( .A(n1210), .Y(n1235) );
  INVX2 U60 ( .A(n1210), .Y(n1234) );
  INVX2 U61 ( .A(n1198), .Y(n1209) );
  INVX1 U62 ( .A(n1183), .Y(N23) );
  INVX1 U63 ( .A(n1174), .Y(N32) );
  INVX1 U64 ( .A(n1176), .Y(N30) );
  INVX1 U65 ( .A(n1177), .Y(N29) );
  INVX1 U66 ( .A(n1179), .Y(N27) );
  INVX1 U67 ( .A(n1182), .Y(N24) );
  INVX1 U68 ( .A(n1184), .Y(N22) );
  INVX1 U69 ( .A(n1185), .Y(N21) );
  INVX1 U70 ( .A(n1186), .Y(N20) );
  INVX1 U71 ( .A(n1189), .Y(N17) );
  BUFX2 U72 ( .A(n125), .Y(n1240) );
  BUFX2 U73 ( .A(n127), .Y(n1244) );
  BUFX2 U74 ( .A(n129), .Y(n1246) );
  BUFX2 U75 ( .A(n131), .Y(n1248) );
  BUFX2 U76 ( .A(n133), .Y(n1250) );
  BUFX2 U77 ( .A(n135), .Y(n1252) );
  BUFX2 U78 ( .A(n137), .Y(n1254) );
  BUFX2 U79 ( .A(n139), .Y(n1257) );
  BUFX2 U80 ( .A(n141), .Y(n1260) );
  BUFX2 U81 ( .A(n143), .Y(n1263) );
  BUFX2 U82 ( .A(n145), .Y(n1266) );
  BUFX2 U83 ( .A(n147), .Y(n1269) );
  BUFX2 U84 ( .A(n149), .Y(n1271) );
  BUFX2 U85 ( .A(n151), .Y(n1273) );
  BUFX2 U86 ( .A(n153), .Y(n1277) );
  BUFX2 U87 ( .A(n155), .Y(n1279) );
  BUFX2 U88 ( .A(n157), .Y(n1281) );
  BUFX2 U89 ( .A(n159), .Y(n1283) );
  BUFX2 U90 ( .A(n161), .Y(n1285) );
  BUFX2 U91 ( .A(n163), .Y(n1287) );
  BUFX2 U92 ( .A(n165), .Y(n1289) );
  BUFX2 U93 ( .A(n167), .Y(n1292) );
  BUFX2 U94 ( .A(n169), .Y(n1294) );
  BUFX2 U95 ( .A(n171), .Y(n1296) );
  BUFX2 U96 ( .A(n173), .Y(n1298) );
  BUFX2 U97 ( .A(n175), .Y(n1300) );
  BUFX2 U98 ( .A(n177), .Y(n1302) );
  BUFX2 U99 ( .A(n179), .Y(n1304) );
  INVX1 U100 ( .A(N12), .Y(n1350) );
  INVX2 U101 ( .A(n1350), .Y(n1196) );
  INVX1 U102 ( .A(n1349), .Y(n1192) );
  INVX1 U103 ( .A(n1192), .Y(n1193) );
  INVX1 U104 ( .A(n1350), .Y(n1195) );
  INVX1 U105 ( .A(n1346), .Y(n1237) );
  INVX1 U106 ( .A(n1237), .Y(n1212) );
  INVX1 U107 ( .A(n1237), .Y(n1213) );
  INVX1 U108 ( .A(n1346), .Y(n1236) );
  INVX1 U109 ( .A(n1352), .Y(n1191) );
  INVX1 U110 ( .A(n1345), .Y(n1210) );
  INVX1 U111 ( .A(N14), .Y(n1353) );
  BUFX2 U112 ( .A(n127), .Y(n1245) );
  INVX1 U113 ( .A(n1352), .Y(n1351) );
  INVX1 U114 ( .A(N13), .Y(n1352) );
  INVX1 U115 ( .A(n1353), .Y(n1190) );
  INVX1 U116 ( .A(n122), .Y(n1291) );
  INVX1 U117 ( .A(n123), .Y(n1306) );
  BUFX2 U118 ( .A(n143), .Y(n1264) );
  BUFX2 U119 ( .A(n145), .Y(n1267) );
  BUFX2 U120 ( .A(n147), .Y(n1270) );
  BUFX2 U121 ( .A(n149), .Y(n1272) );
  BUFX2 U122 ( .A(n151), .Y(n1274) );
  BUFX2 U123 ( .A(n163), .Y(n1288) );
  BUFX2 U124 ( .A(n165), .Y(n1290) );
  BUFX2 U125 ( .A(n153), .Y(n1278) );
  BUFX2 U126 ( .A(n155), .Y(n1280) );
  BUFX2 U127 ( .A(n157), .Y(n1282) );
  BUFX2 U128 ( .A(n159), .Y(n1284) );
  BUFX2 U129 ( .A(n161), .Y(n1286) );
  INVX1 U130 ( .A(n1347), .Y(n1198) );
  BUFX2 U131 ( .A(n125), .Y(n1241) );
  BUFX2 U132 ( .A(n167), .Y(n1293) );
  BUFX2 U133 ( .A(n169), .Y(n1295) );
  BUFX2 U134 ( .A(n171), .Y(n1297) );
  BUFX2 U135 ( .A(n173), .Y(n1299) );
  BUFX2 U136 ( .A(n175), .Y(n1301) );
  BUFX2 U137 ( .A(n177), .Y(n1303) );
  BUFX2 U138 ( .A(n179), .Y(n1305) );
  BUFX2 U139 ( .A(n129), .Y(n1247) );
  BUFX2 U140 ( .A(n131), .Y(n1249) );
  BUFX2 U141 ( .A(n133), .Y(n1251) );
  BUFX2 U142 ( .A(n135), .Y(n1253) );
  BUFX2 U143 ( .A(n137), .Y(n1255) );
  BUFX2 U144 ( .A(n139), .Y(n1258) );
  BUFX2 U145 ( .A(n141), .Y(n1261) );
  INVX1 U146 ( .A(n120), .Y(n1256) );
  INVX1 U147 ( .A(n121), .Y(n1275) );
  INVX1 U148 ( .A(n80), .Y(n2) );
  BUFX2 U149 ( .A(n81), .Y(n3) );
  INVX4 U150 ( .A(n37), .Y(n106) );
  INVX4 U151 ( .A(n36), .Y(n105) );
  INVX4 U152 ( .A(n35), .Y(n104) );
  INVX4 U153 ( .A(n34), .Y(n103) );
  INVX4 U154 ( .A(n33), .Y(n102) );
  INVX4 U155 ( .A(n32), .Y(n101) );
  INVX4 U156 ( .A(n31), .Y(n100) );
  INVX4 U157 ( .A(n30), .Y(n99) );
  INVX4 U158 ( .A(n93), .Y(n1310) );
  BUFX2 U159 ( .A(n55), .Y(n4) );
  INVX1 U160 ( .A(n47), .Y(n5) );
  BUFX2 U161 ( .A(n48), .Y(n6) );
  INVX1 U162 ( .A(n44), .Y(n7) );
  BUFX2 U163 ( .A(n45), .Y(n8) );
  INVX1 U164 ( .A(n71), .Y(n9) );
  BUFX2 U165 ( .A(n73), .Y(n10) );
  INVX1 U166 ( .A(n68), .Y(n11) );
  BUFX2 U167 ( .A(n70), .Y(n12) );
  BUFX2 U168 ( .A(n54), .Y(n13) );
  INVX1 U169 ( .A(n50), .Y(n14) );
  BUFX2 U170 ( .A(n51), .Y(n15) );
  INVX1 U171 ( .A(write), .Y(n16) );
  INVX1 U172 ( .A(write), .Y(n1238) );
  AND2X2 U173 ( .A(n1344), .B(n16), .Y(n17) );
  AND2X2 U174 ( .A(n1344), .B(n1238), .Y(n18) );
  AND2X2 U175 ( .A(\data_in<0> ), .B(n1309), .Y(n19) );
  AND2X2 U176 ( .A(\data_in<1> ), .B(n1309), .Y(n20) );
  AND2X2 U177 ( .A(\data_in<2> ), .B(n1309), .Y(n21) );
  AND2X2 U178 ( .A(\data_in<3> ), .B(n1309), .Y(n22) );
  AND2X2 U179 ( .A(\data_in<4> ), .B(n1309), .Y(n23) );
  AND2X2 U180 ( .A(\data_in<5> ), .B(n1309), .Y(n24) );
  AND2X2 U181 ( .A(\data_in<6> ), .B(n1309), .Y(n25) );
  AND2X2 U182 ( .A(\data_in<7> ), .B(n1309), .Y(n26) );
  AND2X2 U183 ( .A(\data_in<8> ), .B(n1309), .Y(n27) );
  AND2X2 U184 ( .A(\data_in<9> ), .B(n1309), .Y(n28) );
  AND2X2 U185 ( .A(\data_in<10> ), .B(n1309), .Y(n29) );
  AND2X2 U186 ( .A(n1309), .B(n122), .Y(n30) );
  AND2X2 U187 ( .A(n1309), .B(n166), .Y(n31) );
  AND2X2 U188 ( .A(n1309), .B(n168), .Y(n32) );
  AND2X2 U189 ( .A(n1309), .B(n170), .Y(n33) );
  AND2X2 U190 ( .A(n1309), .B(n172), .Y(n34) );
  AND2X2 U191 ( .A(n1309), .B(n174), .Y(n35) );
  AND2X2 U192 ( .A(n1309), .B(n176), .Y(n36) );
  AND2X2 U193 ( .A(n1309), .B(n178), .Y(n37) );
  AND2X2 U194 ( .A(n1344), .B(n16), .Y(n38) );
  AND2X2 U195 ( .A(n1308), .B(n162), .Y(n39) );
  AND2X2 U196 ( .A(n1308), .B(n164), .Y(n40) );
  AND2X2 U197 ( .A(n1308), .B(n123), .Y(n42) );
  AND2X2 U198 ( .A(n1307), .B(n142), .Y(n44) );
  INVX1 U199 ( .A(n44), .Y(n45) );
  INVX1 U200 ( .A(n44), .Y(n46) );
  AND2X2 U201 ( .A(n1307), .B(n144), .Y(n47) );
  INVX1 U202 ( .A(n47), .Y(n48) );
  INVX1 U203 ( .A(n47), .Y(n49) );
  AND2X2 U204 ( .A(n1307), .B(n120), .Y(n50) );
  INVX1 U205 ( .A(n50), .Y(n51) );
  INVX1 U206 ( .A(n50), .Y(n52) );
  AND2X2 U207 ( .A(n1307), .B(n124), .Y(n53) );
  INVX1 U208 ( .A(n53), .Y(n54) );
  INVX1 U209 ( .A(n53), .Y(n55) );
  AND2X2 U210 ( .A(n1307), .B(n126), .Y(n56) );
  AND2X2 U211 ( .A(n1307), .B(n128), .Y(n58) );
  AND2X2 U212 ( .A(n1307), .B(n130), .Y(n60) );
  AND2X2 U213 ( .A(n1307), .B(n132), .Y(n62) );
  AND2X2 U214 ( .A(n1307), .B(n134), .Y(n64) );
  AND2X2 U215 ( .A(n1307), .B(n136), .Y(n66) );
  AND2X2 U216 ( .A(n1307), .B(n138), .Y(n68) );
  INVX1 U217 ( .A(n68), .Y(n69) );
  INVX1 U218 ( .A(n68), .Y(n70) );
  AND2X2 U219 ( .A(n1307), .B(n140), .Y(n71) );
  INVX1 U220 ( .A(n71), .Y(n72) );
  INVX1 U221 ( .A(n71), .Y(n73) );
  AND2X2 U222 ( .A(n1308), .B(n146), .Y(n74) );
  AND2X2 U223 ( .A(n1308), .B(n148), .Y(n76) );
  AND2X2 U224 ( .A(n1308), .B(n150), .Y(n78) );
  AND2X2 U225 ( .A(n1308), .B(n121), .Y(n80) );
  INVX1 U226 ( .A(n80), .Y(n81) );
  INVX1 U227 ( .A(n80), .Y(n82) );
  AND2X2 U228 ( .A(n1308), .B(n152), .Y(n83) );
  AND2X2 U229 ( .A(n1308), .B(n154), .Y(n85) );
  AND2X2 U230 ( .A(n1308), .B(n156), .Y(n87) );
  AND2X2 U231 ( .A(n1308), .B(n158), .Y(n89) );
  AND2X2 U232 ( .A(n1308), .B(n160), .Y(n91) );
  AND2X2 U233 ( .A(n1344), .B(write), .Y(n93) );
  AND2X2 U234 ( .A(\data_in<11> ), .B(n1309), .Y(n94) );
  AND2X2 U235 ( .A(\data_in<12> ), .B(n1309), .Y(n95) );
  AND2X2 U236 ( .A(\data_in<13> ), .B(n1309), .Y(n96) );
  AND2X2 U237 ( .A(\data_in<14> ), .B(n1309), .Y(n97) );
  AND2X2 U238 ( .A(\data_in<15> ), .B(n1309), .Y(n98) );
  INVX1 U239 ( .A(n1350), .Y(n1349) );
  INVX1 U240 ( .A(n1346), .Y(n1345) );
  AND2X1 U241 ( .A(n1349), .B(n1347), .Y(n107) );
  INVX1 U242 ( .A(n1348), .Y(n1347) );
  AND2X1 U243 ( .A(n2393), .B(N14), .Y(n108) );
  BUFX2 U244 ( .A(n1386), .Y(n109) );
  INVX1 U245 ( .A(n109), .Y(n1778) );
  BUFX2 U246 ( .A(n1403), .Y(n110) );
  INVX1 U247 ( .A(n110), .Y(n1795) );
  BUFX2 U248 ( .A(n1420), .Y(n111) );
  INVX1 U249 ( .A(n111), .Y(n1812) );
  BUFX2 U250 ( .A(n1437), .Y(n112) );
  INVX1 U251 ( .A(n112), .Y(n1829) );
  BUFX2 U252 ( .A(n1454), .Y(n113) );
  INVX1 U253 ( .A(n113), .Y(n1846) );
  BUFX2 U254 ( .A(n1615), .Y(n114) );
  INVX1 U255 ( .A(n114), .Y(n1728) );
  BUFX2 U256 ( .A(n1745), .Y(n115) );
  INVX1 U257 ( .A(n115), .Y(n1863) );
  AND2X1 U258 ( .A(n1345), .B(n107), .Y(n116) );
  AND2X1 U259 ( .A(n1351), .B(n108), .Y(n117) );
  AND2X1 U260 ( .A(n1346), .B(n107), .Y(n118) );
  AND2X1 U261 ( .A(n1352), .B(n108), .Y(n119) );
  AND2X1 U262 ( .A(n117), .B(n1864), .Y(n120) );
  AND2X1 U263 ( .A(n1864), .B(n119), .Y(n121) );
  AND2X1 U264 ( .A(n1864), .B(n1728), .Y(n122) );
  AND2X1 U265 ( .A(n1864), .B(n1863), .Y(n123) );
  AND2X1 U266 ( .A(n116), .B(n117), .Y(n124) );
  INVX1 U267 ( .A(n124), .Y(n125) );
  AND2X1 U268 ( .A(n117), .B(n118), .Y(n126) );
  INVX1 U269 ( .A(n126), .Y(n127) );
  AND2X1 U270 ( .A(n117), .B(n1778), .Y(n128) );
  INVX1 U271 ( .A(n128), .Y(n129) );
  AND2X1 U272 ( .A(n117), .B(n1795), .Y(n130) );
  INVX1 U273 ( .A(n130), .Y(n131) );
  AND2X1 U274 ( .A(n117), .B(n1812), .Y(n132) );
  INVX1 U275 ( .A(n132), .Y(n133) );
  AND2X1 U276 ( .A(n117), .B(n1829), .Y(n134) );
  INVX1 U277 ( .A(n134), .Y(n135) );
  AND2X1 U278 ( .A(n117), .B(n1846), .Y(n136) );
  INVX1 U279 ( .A(n136), .Y(n137) );
  AND2X1 U280 ( .A(n116), .B(n119), .Y(n138) );
  INVX1 U281 ( .A(n138), .Y(n139) );
  AND2X1 U282 ( .A(n118), .B(n119), .Y(n140) );
  INVX1 U283 ( .A(n140), .Y(n141) );
  AND2X1 U284 ( .A(n1778), .B(n119), .Y(n142) );
  INVX1 U285 ( .A(n142), .Y(n143) );
  AND2X1 U286 ( .A(n1795), .B(n119), .Y(n144) );
  INVX1 U287 ( .A(n144), .Y(n145) );
  AND2X1 U288 ( .A(n1812), .B(n119), .Y(n146) );
  INVX1 U289 ( .A(n146), .Y(n147) );
  AND2X1 U290 ( .A(n1829), .B(n119), .Y(n148) );
  INVX1 U291 ( .A(n148), .Y(n149) );
  AND2X1 U292 ( .A(n1846), .B(n119), .Y(n150) );
  INVX1 U293 ( .A(n150), .Y(n151) );
  AND2X1 U294 ( .A(n116), .B(n1728), .Y(n152) );
  INVX1 U295 ( .A(n152), .Y(n153) );
  AND2X1 U296 ( .A(n118), .B(n1728), .Y(n154) );
  INVX1 U297 ( .A(n154), .Y(n155) );
  AND2X1 U298 ( .A(n1778), .B(n1728), .Y(n156) );
  INVX1 U299 ( .A(n156), .Y(n157) );
  AND2X1 U300 ( .A(n1795), .B(n1728), .Y(n158) );
  INVX1 U301 ( .A(n158), .Y(n159) );
  AND2X1 U302 ( .A(n1812), .B(n1728), .Y(n160) );
  INVX1 U303 ( .A(n160), .Y(n161) );
  AND2X1 U304 ( .A(n1829), .B(n1728), .Y(n162) );
  INVX1 U305 ( .A(n162), .Y(n163) );
  AND2X1 U306 ( .A(n1846), .B(n1728), .Y(n164) );
  INVX1 U307 ( .A(n164), .Y(n165) );
  AND2X1 U308 ( .A(n116), .B(n1863), .Y(n166) );
  INVX1 U309 ( .A(n166), .Y(n167) );
  AND2X1 U310 ( .A(n118), .B(n1863), .Y(n168) );
  INVX1 U311 ( .A(n168), .Y(n169) );
  AND2X1 U312 ( .A(n1778), .B(n1863), .Y(n170) );
  INVX1 U313 ( .A(n170), .Y(n171) );
  AND2X1 U314 ( .A(n1795), .B(n1863), .Y(n172) );
  INVX1 U315 ( .A(n172), .Y(n173) );
  AND2X1 U316 ( .A(n1812), .B(n1863), .Y(n174) );
  INVX1 U317 ( .A(n174), .Y(n175) );
  AND2X1 U318 ( .A(n1829), .B(n1863), .Y(n176) );
  INVX1 U319 ( .A(n176), .Y(n177) );
  AND2X1 U320 ( .A(n1846), .B(n1863), .Y(n178) );
  INVX1 U321 ( .A(n178), .Y(n179) );
  BUFX2 U322 ( .A(n51), .Y(n180) );
  BUFX2 U323 ( .A(n81), .Y(n1276) );
  BUFX2 U324 ( .A(n48), .Y(n1268) );
  BUFX2 U325 ( .A(n45), .Y(n1265) );
  BUFX2 U326 ( .A(n73), .Y(n1262) );
  BUFX2 U327 ( .A(n70), .Y(n1259) );
  INVX4 U328 ( .A(n1311), .Y(n1307) );
  BUFX2 U329 ( .A(n55), .Y(n1243) );
  BUFX2 U330 ( .A(n54), .Y(n1242) );
  INVX1 U331 ( .A(N11), .Y(n1348) );
  MUX2X1 U332 ( .B(n182), .A(n183), .S(n1199), .Y(n181) );
  MUX2X1 U333 ( .B(n185), .A(n186), .S(n1199), .Y(n184) );
  MUX2X1 U334 ( .B(n188), .A(n189), .S(n1199), .Y(n187) );
  MUX2X1 U335 ( .B(n191), .A(n192), .S(n1199), .Y(n190) );
  MUX2X1 U336 ( .B(n194), .A(n195), .S(n1191), .Y(n193) );
  MUX2X1 U337 ( .B(n197), .A(n198), .S(n1199), .Y(n196) );
  MUX2X1 U338 ( .B(n200), .A(n201), .S(n1199), .Y(n199) );
  MUX2X1 U339 ( .B(n203), .A(n204), .S(n1199), .Y(n202) );
  MUX2X1 U340 ( .B(n206), .A(n207), .S(n1199), .Y(n205) );
  MUX2X1 U341 ( .B(n209), .A(n210), .S(n1191), .Y(n208) );
  MUX2X1 U342 ( .B(n212), .A(n213), .S(n1200), .Y(n211) );
  MUX2X1 U343 ( .B(n216), .A(n217), .S(n1200), .Y(n215) );
  MUX2X1 U344 ( .B(n219), .A(n220), .S(n1200), .Y(n218) );
  MUX2X1 U345 ( .B(n222), .A(n223), .S(n1200), .Y(n221) );
  MUX2X1 U346 ( .B(n225), .A(n226), .S(n1191), .Y(n224) );
  MUX2X1 U347 ( .B(n228), .A(n229), .S(n1200), .Y(n227) );
  MUX2X1 U348 ( .B(n231), .A(n232), .S(n1200), .Y(n230) );
  MUX2X1 U349 ( .B(n234), .A(n235), .S(n1200), .Y(n233) );
  MUX2X1 U350 ( .B(n237), .A(n238), .S(n1200), .Y(n236) );
  MUX2X1 U351 ( .B(n240), .A(n241), .S(n1191), .Y(n239) );
  MUX2X1 U352 ( .B(n243), .A(n244), .S(n1200), .Y(n242) );
  MUX2X1 U353 ( .B(n246), .A(n247), .S(n1200), .Y(n245) );
  MUX2X1 U354 ( .B(n249), .A(n250), .S(n1200), .Y(n248) );
  MUX2X1 U355 ( .B(n252), .A(n253), .S(n1200), .Y(n251) );
  MUX2X1 U356 ( .B(n255), .A(n256), .S(n1191), .Y(n254) );
  MUX2X1 U357 ( .B(n258), .A(n259), .S(n1201), .Y(n257) );
  MUX2X1 U358 ( .B(n261), .A(n262), .S(n1201), .Y(n260) );
  MUX2X1 U359 ( .B(n264), .A(n265), .S(n1201), .Y(n263) );
  MUX2X1 U360 ( .B(n267), .A(n268), .S(n1201), .Y(n266) );
  MUX2X1 U361 ( .B(n270), .A(n271), .S(n1191), .Y(n269) );
  MUX2X1 U362 ( .B(n273), .A(n274), .S(n1201), .Y(n272) );
  MUX2X1 U363 ( .B(n276), .A(n277), .S(n1201), .Y(n275) );
  MUX2X1 U364 ( .B(n279), .A(n280), .S(n1201), .Y(n278) );
  MUX2X1 U365 ( .B(n282), .A(n283), .S(n1201), .Y(n281) );
  MUX2X1 U366 ( .B(n285), .A(n286), .S(n1191), .Y(n284) );
  MUX2X1 U367 ( .B(n288), .A(n289), .S(n1201), .Y(n287) );
  MUX2X1 U368 ( .B(n291), .A(n292), .S(n1201), .Y(n290) );
  MUX2X1 U369 ( .B(n294), .A(n295), .S(n1201), .Y(n293) );
  MUX2X1 U370 ( .B(n297), .A(n298), .S(n1201), .Y(n296) );
  MUX2X1 U371 ( .B(n300), .A(n301), .S(n1191), .Y(n299) );
  MUX2X1 U372 ( .B(n303), .A(n304), .S(n1202), .Y(n302) );
  MUX2X1 U373 ( .B(n306), .A(n307), .S(n1202), .Y(n305) );
  MUX2X1 U374 ( .B(n309), .A(n310), .S(n1202), .Y(n308) );
  MUX2X1 U375 ( .B(n312), .A(n313), .S(n1202), .Y(n311) );
  MUX2X1 U376 ( .B(n315), .A(n316), .S(n1191), .Y(n314) );
  MUX2X1 U377 ( .B(n318), .A(n319), .S(n1202), .Y(n317) );
  MUX2X1 U378 ( .B(n321), .A(n322), .S(n1202), .Y(n320) );
  MUX2X1 U379 ( .B(n324), .A(n325), .S(n1202), .Y(n323) );
  MUX2X1 U380 ( .B(n327), .A(n328), .S(n1202), .Y(n326) );
  MUX2X1 U381 ( .B(n330), .A(n331), .S(n1191), .Y(n329) );
  MUX2X1 U382 ( .B(n333), .A(n334), .S(n1202), .Y(n332) );
  MUX2X1 U383 ( .B(n336), .A(n337), .S(n1202), .Y(n335) );
  MUX2X1 U384 ( .B(n339), .A(n340), .S(n1202), .Y(n338) );
  MUX2X1 U385 ( .B(n342), .A(n343), .S(n1202), .Y(n341) );
  MUX2X1 U386 ( .B(n345), .A(n346), .S(n1191), .Y(n344) );
  MUX2X1 U387 ( .B(n348), .A(n349), .S(n1203), .Y(n347) );
  MUX2X1 U388 ( .B(n351), .A(n352), .S(n1203), .Y(n350) );
  MUX2X1 U389 ( .B(n354), .A(n355), .S(n1203), .Y(n353) );
  MUX2X1 U390 ( .B(n357), .A(n358), .S(n1203), .Y(n356) );
  MUX2X1 U391 ( .B(n360), .A(n361), .S(n1191), .Y(n359) );
  MUX2X1 U392 ( .B(n363), .A(n364), .S(n1203), .Y(n362) );
  MUX2X1 U393 ( .B(n366), .A(n367), .S(n1203), .Y(n365) );
  MUX2X1 U394 ( .B(n369), .A(n370), .S(n1203), .Y(n368) );
  MUX2X1 U395 ( .B(n372), .A(n373), .S(n1203), .Y(n371) );
  MUX2X1 U396 ( .B(n375), .A(n376), .S(n1351), .Y(n374) );
  MUX2X1 U397 ( .B(n378), .A(n379), .S(n1203), .Y(n377) );
  MUX2X1 U398 ( .B(n381), .A(n382), .S(n1203), .Y(n380) );
  MUX2X1 U399 ( .B(n384), .A(n385), .S(n1203), .Y(n383) );
  MUX2X1 U400 ( .B(n387), .A(n388), .S(n1203), .Y(n386) );
  MUX2X1 U401 ( .B(n390), .A(n391), .S(n1351), .Y(n389) );
  MUX2X1 U402 ( .B(n393), .A(n394), .S(n1204), .Y(n392) );
  MUX2X1 U403 ( .B(n396), .A(n397), .S(n1204), .Y(n395) );
  MUX2X1 U404 ( .B(n399), .A(n400), .S(n1204), .Y(n398) );
  MUX2X1 U405 ( .B(n402), .A(n403), .S(n1204), .Y(n401) );
  MUX2X1 U406 ( .B(n405), .A(n406), .S(n1351), .Y(n404) );
  MUX2X1 U407 ( .B(n408), .A(n409), .S(n1204), .Y(n407) );
  MUX2X1 U408 ( .B(n411), .A(n412), .S(n1204), .Y(n410) );
  MUX2X1 U409 ( .B(n414), .A(n415), .S(n1204), .Y(n413) );
  MUX2X1 U410 ( .B(n417), .A(n418), .S(n1204), .Y(n416) );
  MUX2X1 U411 ( .B(n420), .A(n421), .S(n1351), .Y(n419) );
  MUX2X1 U412 ( .B(n423), .A(n424), .S(n1204), .Y(n422) );
  MUX2X1 U413 ( .B(n426), .A(n427), .S(n1204), .Y(n425) );
  MUX2X1 U414 ( .B(n429), .A(n430), .S(n1204), .Y(n428) );
  MUX2X1 U415 ( .B(n432), .A(n433), .S(n1204), .Y(n431) );
  MUX2X1 U416 ( .B(n435), .A(n436), .S(n1351), .Y(n434) );
  MUX2X1 U417 ( .B(n438), .A(n439), .S(n1205), .Y(n437) );
  MUX2X1 U418 ( .B(n441), .A(n442), .S(n1205), .Y(n440) );
  MUX2X1 U419 ( .B(n444), .A(n445), .S(n1205), .Y(n443) );
  MUX2X1 U420 ( .B(n447), .A(n448), .S(n1205), .Y(n446) );
  MUX2X1 U421 ( .B(n450), .A(n451), .S(n1351), .Y(n449) );
  MUX2X1 U422 ( .B(n453), .A(n454), .S(n1205), .Y(n452) );
  MUX2X1 U423 ( .B(n456), .A(n457), .S(n1205), .Y(n455) );
  MUX2X1 U424 ( .B(n459), .A(n460), .S(n1205), .Y(n458) );
  MUX2X1 U425 ( .B(n462), .A(n463), .S(n1205), .Y(n461) );
  MUX2X1 U426 ( .B(n465), .A(n466), .S(n1351), .Y(n464) );
  MUX2X1 U427 ( .B(n468), .A(n469), .S(n1205), .Y(n467) );
  MUX2X1 U428 ( .B(n471), .A(n472), .S(n1205), .Y(n470) );
  MUX2X1 U429 ( .B(n474), .A(n475), .S(n1205), .Y(n473) );
  MUX2X1 U430 ( .B(n477), .A(n478), .S(n1205), .Y(n476) );
  MUX2X1 U431 ( .B(n480), .A(n481), .S(n1351), .Y(n479) );
  MUX2X1 U432 ( .B(n483), .A(n484), .S(n1206), .Y(n482) );
  MUX2X1 U433 ( .B(n486), .A(n487), .S(n1206), .Y(n485) );
  MUX2X1 U434 ( .B(n489), .A(n490), .S(n1206), .Y(n488) );
  MUX2X1 U435 ( .B(n492), .A(n493), .S(n1206), .Y(n491) );
  MUX2X1 U436 ( .B(n495), .A(n496), .S(n1351), .Y(n494) );
  MUX2X1 U437 ( .B(n498), .A(n499), .S(n1206), .Y(n497) );
  MUX2X1 U438 ( .B(n501), .A(n502), .S(n1206), .Y(n500) );
  MUX2X1 U439 ( .B(n504), .A(n505), .S(n1206), .Y(n503) );
  MUX2X1 U440 ( .B(n507), .A(n508), .S(n1206), .Y(n506) );
  MUX2X1 U441 ( .B(n510), .A(n511), .S(n1351), .Y(n509) );
  MUX2X1 U442 ( .B(n513), .A(n514), .S(n1206), .Y(n512) );
  MUX2X1 U443 ( .B(n516), .A(n517), .S(n1206), .Y(n515) );
  MUX2X1 U444 ( .B(n519), .A(n520), .S(n1206), .Y(n518) );
  MUX2X1 U445 ( .B(n522), .A(n523), .S(n1206), .Y(n521) );
  MUX2X1 U446 ( .B(n525), .A(n526), .S(n1351), .Y(n524) );
  MUX2X1 U447 ( .B(n528), .A(n529), .S(n1207), .Y(n527) );
  MUX2X1 U448 ( .B(n531), .A(n532), .S(n1207), .Y(n530) );
  MUX2X1 U449 ( .B(n534), .A(n535), .S(n1207), .Y(n533) );
  MUX2X1 U450 ( .B(n537), .A(n538), .S(n1207), .Y(n536) );
  MUX2X1 U451 ( .B(n540), .A(n541), .S(n1351), .Y(n539) );
  MUX2X1 U452 ( .B(n543), .A(n544), .S(n1207), .Y(n542) );
  MUX2X1 U453 ( .B(n546), .A(n547), .S(n1207), .Y(n545) );
  MUX2X1 U454 ( .B(n549), .A(n550), .S(n1207), .Y(n548) );
  MUX2X1 U455 ( .B(n552), .A(n553), .S(n1207), .Y(n551) );
  MUX2X1 U456 ( .B(n555), .A(n556), .S(n1191), .Y(n554) );
  MUX2X1 U457 ( .B(n558), .A(n559), .S(n1207), .Y(n557) );
  MUX2X1 U458 ( .B(n561), .A(n562), .S(n1207), .Y(n560) );
  MUX2X1 U459 ( .B(n564), .A(n565), .S(n1207), .Y(n563) );
  MUX2X1 U460 ( .B(n567), .A(n568), .S(n1207), .Y(n566) );
  MUX2X1 U461 ( .B(n570), .A(n571), .S(n1191), .Y(n569) );
  MUX2X1 U462 ( .B(n573), .A(n574), .S(n1208), .Y(n572) );
  MUX2X1 U463 ( .B(n576), .A(n577), .S(n1208), .Y(n575) );
  MUX2X1 U464 ( .B(n579), .A(n580), .S(n1208), .Y(n578) );
  MUX2X1 U465 ( .B(n582), .A(n583), .S(n1208), .Y(n581) );
  MUX2X1 U466 ( .B(n585), .A(n586), .S(n1191), .Y(n584) );
  MUX2X1 U467 ( .B(n588), .A(n589), .S(n1208), .Y(n587) );
  MUX2X1 U468 ( .B(n591), .A(n592), .S(n1208), .Y(n590) );
  MUX2X1 U469 ( .B(n594), .A(n595), .S(n1208), .Y(n593) );
  MUX2X1 U470 ( .B(n597), .A(n598), .S(n1208), .Y(n596) );
  MUX2X1 U471 ( .B(n600), .A(n601), .S(n1191), .Y(n599) );
  MUX2X1 U472 ( .B(n603), .A(n604), .S(n1208), .Y(n602) );
  MUX2X1 U473 ( .B(n606), .A(n607), .S(n1208), .Y(n605) );
  MUX2X1 U474 ( .B(n609), .A(n610), .S(n1208), .Y(n608) );
  MUX2X1 U475 ( .B(n612), .A(n613), .S(n1208), .Y(n611) );
  MUX2X1 U476 ( .B(n615), .A(n616), .S(n1191), .Y(n614) );
  MUX2X1 U477 ( .B(n618), .A(n619), .S(n1209), .Y(n617) );
  MUX2X1 U478 ( .B(n621), .A(n622), .S(n1209), .Y(n620) );
  MUX2X1 U479 ( .B(n624), .A(n625), .S(n1209), .Y(n623) );
  MUX2X1 U480 ( .B(n627), .A(n628), .S(n1209), .Y(n626) );
  MUX2X1 U481 ( .B(n630), .A(n631), .S(n1191), .Y(n629) );
  MUX2X1 U482 ( .B(n633), .A(n634), .S(n1209), .Y(n632) );
  MUX2X1 U483 ( .B(n636), .A(n637), .S(n1209), .Y(n635) );
  MUX2X1 U484 ( .B(n639), .A(n640), .S(n1209), .Y(n638) );
  MUX2X1 U485 ( .B(n642), .A(n643), .S(n1209), .Y(n641) );
  MUX2X1 U486 ( .B(n645), .A(n646), .S(n1191), .Y(n644) );
  MUX2X1 U487 ( .B(n648), .A(n649), .S(n1209), .Y(n647) );
  MUX2X1 U488 ( .B(n1163), .A(n1164), .S(n1209), .Y(n650) );
  MUX2X1 U489 ( .B(n1166), .A(n1167), .S(n1209), .Y(n1165) );
  MUX2X1 U490 ( .B(n1169), .A(n1170), .S(n1209), .Y(n1168) );
  MUX2X1 U491 ( .B(n1172), .A(n1173), .S(n1191), .Y(n1171) );
  MUX2X1 U492 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1214), .Y(n183) );
  MUX2X1 U493 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1214), .Y(n182) );
  MUX2X1 U494 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1214), .Y(n186) );
  MUX2X1 U495 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1214), .Y(n185) );
  MUX2X1 U496 ( .B(n184), .A(n181), .S(n1196), .Y(n195) );
  MUX2X1 U497 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1215), .Y(n189) );
  MUX2X1 U498 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1215), .Y(n188) );
  MUX2X1 U499 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1215), .Y(n192) );
  MUX2X1 U500 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1215), .Y(n191) );
  MUX2X1 U501 ( .B(n190), .A(n187), .S(n1196), .Y(n194) );
  MUX2X1 U502 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1215), .Y(n198) );
  MUX2X1 U503 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1215), .Y(n197) );
  MUX2X1 U504 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1215), .Y(n201) );
  MUX2X1 U505 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1215), .Y(n200) );
  MUX2X1 U506 ( .B(n199), .A(n196), .S(n1196), .Y(n210) );
  MUX2X1 U507 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1215), .Y(n204) );
  MUX2X1 U508 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1215), .Y(n203) );
  MUX2X1 U509 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1215), .Y(n207) );
  MUX2X1 U510 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1215), .Y(n206) );
  MUX2X1 U511 ( .B(n205), .A(n202), .S(n1196), .Y(n209) );
  MUX2X1 U512 ( .B(n208), .A(n193), .S(n1190), .Y(n1174) );
  MUX2X1 U513 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1216), .Y(n213) );
  MUX2X1 U514 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1216), .Y(n212) );
  MUX2X1 U515 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1216), .Y(n217) );
  MUX2X1 U516 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1216), .Y(n216) );
  MUX2X1 U517 ( .B(n215), .A(n211), .S(n1196), .Y(n226) );
  MUX2X1 U518 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1216), .Y(n220) );
  MUX2X1 U519 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1216), .Y(n219) );
  MUX2X1 U520 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1216), .Y(n223) );
  MUX2X1 U521 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1216), .Y(n222) );
  MUX2X1 U522 ( .B(n221), .A(n218), .S(n1196), .Y(n225) );
  MUX2X1 U523 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1216), .Y(n229) );
  MUX2X1 U524 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1216), .Y(n228) );
  MUX2X1 U525 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1216), .Y(n232) );
  MUX2X1 U526 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1216), .Y(n231) );
  MUX2X1 U527 ( .B(n230), .A(n227), .S(n1196), .Y(n241) );
  MUX2X1 U528 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1217), .Y(n235) );
  MUX2X1 U529 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1217), .Y(n234) );
  MUX2X1 U530 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1217), .Y(n238) );
  MUX2X1 U531 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1217), .Y(n237) );
  MUX2X1 U532 ( .B(n236), .A(n233), .S(n1196), .Y(n240) );
  MUX2X1 U533 ( .B(n239), .A(n224), .S(n1190), .Y(n1175) );
  MUX2X1 U534 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1217), .Y(n244) );
  MUX2X1 U535 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1217), .Y(n243) );
  MUX2X1 U536 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1217), .Y(n247) );
  MUX2X1 U537 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1217), .Y(n246) );
  MUX2X1 U538 ( .B(n245), .A(n242), .S(n1196), .Y(n256) );
  MUX2X1 U539 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1217), .Y(n250) );
  MUX2X1 U540 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1217), .Y(n249) );
  MUX2X1 U541 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1217), .Y(n253) );
  MUX2X1 U542 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1217), .Y(n252) );
  MUX2X1 U543 ( .B(n251), .A(n248), .S(n1196), .Y(n255) );
  MUX2X1 U544 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1218), .Y(n259) );
  MUX2X1 U545 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1218), .Y(n258) );
  MUX2X1 U546 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1218), .Y(n262) );
  MUX2X1 U547 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1218), .Y(n261) );
  MUX2X1 U548 ( .B(n260), .A(n257), .S(n1196), .Y(n271) );
  MUX2X1 U549 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1218), .Y(n265) );
  MUX2X1 U550 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1218), .Y(n264) );
  MUX2X1 U551 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1218), .Y(n268) );
  MUX2X1 U552 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1218), .Y(n267) );
  MUX2X1 U553 ( .B(n266), .A(n263), .S(n1196), .Y(n270) );
  MUX2X1 U554 ( .B(n269), .A(n254), .S(n1190), .Y(n1176) );
  MUX2X1 U555 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1218), .Y(n274) );
  MUX2X1 U556 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1218), .Y(n273) );
  MUX2X1 U557 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1218), .Y(n277) );
  MUX2X1 U558 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1218), .Y(n276) );
  MUX2X1 U559 ( .B(n275), .A(n272), .S(n1196), .Y(n286) );
  MUX2X1 U560 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1219), .Y(n280) );
  MUX2X1 U561 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1219), .Y(n279) );
  MUX2X1 U562 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1219), .Y(n283) );
  MUX2X1 U563 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1219), .Y(n282) );
  MUX2X1 U564 ( .B(n281), .A(n278), .S(n1196), .Y(n285) );
  MUX2X1 U565 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1219), .Y(n289) );
  MUX2X1 U566 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1219), .Y(n288) );
  MUX2X1 U567 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1219), .Y(n292) );
  MUX2X1 U568 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1219), .Y(n291) );
  MUX2X1 U569 ( .B(n290), .A(n287), .S(n1196), .Y(n301) );
  MUX2X1 U570 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1219), .Y(n295) );
  MUX2X1 U571 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1219), .Y(n294) );
  MUX2X1 U572 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1219), .Y(n298) );
  MUX2X1 U573 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1219), .Y(n297) );
  MUX2X1 U574 ( .B(n296), .A(n293), .S(n1196), .Y(n300) );
  MUX2X1 U575 ( .B(n299), .A(n284), .S(n1190), .Y(n1177) );
  MUX2X1 U576 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1220), .Y(n304) );
  MUX2X1 U577 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1220), .Y(n303) );
  MUX2X1 U578 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1220), .Y(n307) );
  MUX2X1 U579 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1220), .Y(n306) );
  MUX2X1 U580 ( .B(n305), .A(n302), .S(n1196), .Y(n316) );
  MUX2X1 U581 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1220), .Y(n310) );
  MUX2X1 U582 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1220), .Y(n309) );
  MUX2X1 U583 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1220), .Y(n313) );
  MUX2X1 U584 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1220), .Y(n312) );
  MUX2X1 U585 ( .B(n311), .A(n308), .S(n1196), .Y(n315) );
  MUX2X1 U586 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1220), .Y(n319) );
  MUX2X1 U587 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1220), .Y(n318) );
  MUX2X1 U588 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1220), .Y(n322) );
  MUX2X1 U589 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1220), .Y(n321) );
  MUX2X1 U590 ( .B(n320), .A(n317), .S(n1196), .Y(n331) );
  MUX2X1 U591 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1221), .Y(n325) );
  MUX2X1 U592 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1221), .Y(n324) );
  MUX2X1 U593 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1221), .Y(n328) );
  MUX2X1 U594 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1221), .Y(n327) );
  MUX2X1 U595 ( .B(n326), .A(n323), .S(n1196), .Y(n330) );
  MUX2X1 U596 ( .B(n329), .A(n314), .S(n1190), .Y(n1178) );
  MUX2X1 U597 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1221), .Y(n334) );
  MUX2X1 U598 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1221), .Y(n333) );
  MUX2X1 U599 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1221), .Y(n337) );
  MUX2X1 U600 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1221), .Y(n336) );
  MUX2X1 U601 ( .B(n335), .A(n332), .S(n1196), .Y(n346) );
  MUX2X1 U602 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1221), .Y(n340) );
  MUX2X1 U603 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1221), .Y(n339) );
  MUX2X1 U604 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1221), .Y(n343) );
  MUX2X1 U605 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1221), .Y(n342) );
  MUX2X1 U606 ( .B(n341), .A(n338), .S(n1196), .Y(n345) );
  MUX2X1 U607 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1222), .Y(n349) );
  MUX2X1 U608 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1222), .Y(n348) );
  MUX2X1 U609 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1222), .Y(n352) );
  MUX2X1 U610 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1222), .Y(n351) );
  MUX2X1 U611 ( .B(n350), .A(n347), .S(n1196), .Y(n361) );
  MUX2X1 U612 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1222), .Y(n355) );
  MUX2X1 U613 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1222), .Y(n354) );
  MUX2X1 U614 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1222), .Y(n358) );
  MUX2X1 U615 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1222), .Y(n357) );
  MUX2X1 U616 ( .B(n356), .A(n353), .S(n1196), .Y(n360) );
  MUX2X1 U617 ( .B(n359), .A(n344), .S(n1190), .Y(n1179) );
  MUX2X1 U618 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1222), .Y(n364) );
  MUX2X1 U619 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1222), .Y(n363) );
  MUX2X1 U620 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1222), .Y(n367) );
  MUX2X1 U621 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1222), .Y(n366) );
  MUX2X1 U622 ( .B(n365), .A(n362), .S(n1195), .Y(n376) );
  MUX2X1 U623 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1223), .Y(n370) );
  MUX2X1 U624 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1223), .Y(n369) );
  MUX2X1 U625 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1223), .Y(n373) );
  MUX2X1 U626 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1223), .Y(n372) );
  MUX2X1 U627 ( .B(n371), .A(n368), .S(n1195), .Y(n375) );
  MUX2X1 U628 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1223), .Y(n379) );
  MUX2X1 U629 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1223), .Y(n378) );
  MUX2X1 U630 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1223), .Y(n382) );
  MUX2X1 U631 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1223), .Y(n381) );
  MUX2X1 U632 ( .B(n380), .A(n377), .S(n1195), .Y(n391) );
  MUX2X1 U633 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1223), .Y(n385) );
  MUX2X1 U634 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1223), .Y(n384) );
  MUX2X1 U635 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1223), .Y(n388) );
  MUX2X1 U636 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1223), .Y(n387) );
  MUX2X1 U637 ( .B(n386), .A(n383), .S(n1195), .Y(n390) );
  MUX2X1 U638 ( .B(n389), .A(n374), .S(n1190), .Y(n1180) );
  MUX2X1 U639 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1224), .Y(n394) );
  MUX2X1 U640 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1224), .Y(n393) );
  MUX2X1 U641 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1224), .Y(n397) );
  MUX2X1 U642 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1224), .Y(n396) );
  MUX2X1 U643 ( .B(n395), .A(n392), .S(n1195), .Y(n406) );
  MUX2X1 U644 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1224), .Y(n400) );
  MUX2X1 U645 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1224), .Y(n399) );
  MUX2X1 U646 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1224), .Y(n403) );
  MUX2X1 U647 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1224), .Y(n402) );
  MUX2X1 U648 ( .B(n401), .A(n398), .S(n1195), .Y(n405) );
  MUX2X1 U649 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1224), .Y(n409) );
  MUX2X1 U650 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1224), .Y(n408) );
  MUX2X1 U651 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1224), .Y(n412) );
  MUX2X1 U652 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1224), .Y(n411) );
  MUX2X1 U653 ( .B(n410), .A(n407), .S(n1195), .Y(n421) );
  MUX2X1 U654 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1225), .Y(n415) );
  MUX2X1 U655 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1225), .Y(n414) );
  MUX2X1 U656 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1225), .Y(n418) );
  MUX2X1 U657 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1225), .Y(n417) );
  MUX2X1 U658 ( .B(n416), .A(n413), .S(n1195), .Y(n420) );
  MUX2X1 U659 ( .B(n419), .A(n404), .S(n1190), .Y(n1181) );
  MUX2X1 U660 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1225), .Y(n424) );
  MUX2X1 U661 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1225), .Y(n423) );
  MUX2X1 U662 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1225), .Y(n427) );
  MUX2X1 U663 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1225), .Y(n426) );
  MUX2X1 U664 ( .B(n425), .A(n422), .S(n1195), .Y(n436) );
  MUX2X1 U665 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1225), .Y(n430) );
  MUX2X1 U666 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1225), .Y(n429) );
  MUX2X1 U667 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1225), .Y(n433) );
  MUX2X1 U668 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1225), .Y(n432) );
  MUX2X1 U669 ( .B(n431), .A(n428), .S(n1195), .Y(n435) );
  MUX2X1 U670 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1226), .Y(n439) );
  MUX2X1 U671 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1226), .Y(n438) );
  MUX2X1 U672 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1226), .Y(n442) );
  MUX2X1 U673 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1226), .Y(n441) );
  MUX2X1 U674 ( .B(n440), .A(n437), .S(n1195), .Y(n451) );
  MUX2X1 U675 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1226), .Y(n445) );
  MUX2X1 U676 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1226), .Y(n444) );
  MUX2X1 U677 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1226), .Y(n448) );
  MUX2X1 U678 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1226), .Y(n447) );
  MUX2X1 U679 ( .B(n446), .A(n443), .S(n1195), .Y(n450) );
  MUX2X1 U680 ( .B(n449), .A(n434), .S(n1190), .Y(n1182) );
  MUX2X1 U681 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1226), .Y(n454) );
  MUX2X1 U682 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1226), .Y(n453) );
  MUX2X1 U683 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1226), .Y(n457) );
  MUX2X1 U684 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1226), .Y(n456) );
  MUX2X1 U685 ( .B(n455), .A(n452), .S(n1194), .Y(n466) );
  MUX2X1 U686 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1227), .Y(n460) );
  MUX2X1 U687 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1227), .Y(n459) );
  MUX2X1 U688 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1227), .Y(n463) );
  MUX2X1 U689 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1227), .Y(n462) );
  MUX2X1 U690 ( .B(n461), .A(n458), .S(n1194), .Y(n465) );
  MUX2X1 U691 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1227), .Y(n469) );
  MUX2X1 U692 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1227), .Y(n468) );
  MUX2X1 U693 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1227), .Y(n472) );
  MUX2X1 U694 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1227), .Y(n471) );
  MUX2X1 U695 ( .B(n470), .A(n467), .S(n1194), .Y(n481) );
  MUX2X1 U696 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1227), .Y(n475) );
  MUX2X1 U697 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1227), .Y(n474) );
  MUX2X1 U698 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1227), .Y(n478) );
  MUX2X1 U699 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1227), .Y(n477) );
  MUX2X1 U700 ( .B(n476), .A(n473), .S(n1194), .Y(n480) );
  MUX2X1 U701 ( .B(n479), .A(n464), .S(n1190), .Y(n1183) );
  MUX2X1 U702 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1228), .Y(n484) );
  MUX2X1 U703 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1228), .Y(n483) );
  MUX2X1 U704 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1228), .Y(n487) );
  MUX2X1 U705 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1228), .Y(n486) );
  MUX2X1 U706 ( .B(n485), .A(n482), .S(n1194), .Y(n496) );
  MUX2X1 U707 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1228), .Y(n490) );
  MUX2X1 U708 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1228), .Y(n489) );
  MUX2X1 U709 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1228), .Y(n493) );
  MUX2X1 U710 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1228), .Y(n492) );
  MUX2X1 U711 ( .B(n491), .A(n488), .S(n1194), .Y(n495) );
  MUX2X1 U712 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1228), .Y(n499) );
  MUX2X1 U713 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1228), .Y(n498) );
  MUX2X1 U714 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1228), .Y(n502) );
  MUX2X1 U715 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1228), .Y(n501) );
  MUX2X1 U716 ( .B(n500), .A(n497), .S(n1194), .Y(n511) );
  MUX2X1 U717 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1229), .Y(n505) );
  MUX2X1 U718 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1229), .Y(n504) );
  MUX2X1 U719 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1229), .Y(n508) );
  MUX2X1 U720 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1229), .Y(n507) );
  MUX2X1 U721 ( .B(n506), .A(n503), .S(n1194), .Y(n510) );
  MUX2X1 U722 ( .B(n509), .A(n494), .S(n1190), .Y(n1184) );
  MUX2X1 U723 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1229), .Y(n514) );
  MUX2X1 U724 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1229), .Y(n513) );
  MUX2X1 U725 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1229), .Y(n517) );
  MUX2X1 U726 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1229), .Y(n516) );
  MUX2X1 U727 ( .B(n515), .A(n512), .S(n1194), .Y(n526) );
  MUX2X1 U728 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1229), .Y(n520) );
  MUX2X1 U729 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1229), .Y(n519) );
  MUX2X1 U730 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1229), .Y(n523) );
  MUX2X1 U731 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1229), .Y(n522) );
  MUX2X1 U732 ( .B(n521), .A(n518), .S(n1194), .Y(n525) );
  MUX2X1 U733 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1230), .Y(n529) );
  MUX2X1 U734 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1230), .Y(n528) );
  MUX2X1 U735 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1230), .Y(n532) );
  MUX2X1 U736 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1230), .Y(n531) );
  MUX2X1 U737 ( .B(n530), .A(n527), .S(n1194), .Y(n541) );
  MUX2X1 U738 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1230), .Y(n535) );
  MUX2X1 U739 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1230), .Y(n534) );
  MUX2X1 U740 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1230), .Y(n538) );
  MUX2X1 U741 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1230), .Y(n537) );
  MUX2X1 U742 ( .B(n536), .A(n533), .S(n1194), .Y(n540) );
  MUX2X1 U743 ( .B(n539), .A(n524), .S(n1190), .Y(n1185) );
  MUX2X1 U744 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1230), .Y(n544) );
  MUX2X1 U745 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1230), .Y(n543) );
  MUX2X1 U746 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1230), .Y(n547) );
  MUX2X1 U747 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1230), .Y(n546) );
  MUX2X1 U748 ( .B(n545), .A(n542), .S(n1193), .Y(n556) );
  MUX2X1 U749 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1231), .Y(n550) );
  MUX2X1 U750 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1231), .Y(n549) );
  MUX2X1 U751 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1231), .Y(n553) );
  MUX2X1 U752 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1231), .Y(n552) );
  MUX2X1 U753 ( .B(n551), .A(n548), .S(n1193), .Y(n555) );
  MUX2X1 U754 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1231), .Y(n559) );
  MUX2X1 U755 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1231), .Y(n558) );
  MUX2X1 U756 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1231), .Y(n562) );
  MUX2X1 U757 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1231), .Y(n561) );
  MUX2X1 U758 ( .B(n560), .A(n557), .S(n1193), .Y(n571) );
  MUX2X1 U759 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1231), .Y(n565) );
  MUX2X1 U760 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1231), .Y(n564) );
  MUX2X1 U761 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1231), .Y(n568) );
  MUX2X1 U762 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1231), .Y(n567) );
  MUX2X1 U763 ( .B(n566), .A(n563), .S(n1193), .Y(n570) );
  MUX2X1 U764 ( .B(n569), .A(n554), .S(n1190), .Y(n1186) );
  MUX2X1 U765 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1232), .Y(n574) );
  MUX2X1 U766 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1232), .Y(n573) );
  MUX2X1 U767 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1232), .Y(n577) );
  MUX2X1 U768 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1232), .Y(n576) );
  MUX2X1 U769 ( .B(n575), .A(n572), .S(n1193), .Y(n586) );
  MUX2X1 U770 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1232), .Y(n580) );
  MUX2X1 U771 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1232), .Y(n579) );
  MUX2X1 U772 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1232), .Y(n583) );
  MUX2X1 U773 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1232), .Y(n582) );
  MUX2X1 U774 ( .B(n581), .A(n578), .S(n1195), .Y(n585) );
  MUX2X1 U775 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1232), .Y(n589) );
  MUX2X1 U776 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1232), .Y(n588) );
  MUX2X1 U777 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1232), .Y(n592) );
  MUX2X1 U778 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1232), .Y(n591) );
  MUX2X1 U779 ( .B(n590), .A(n587), .S(n1193), .Y(n601) );
  MUX2X1 U780 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1233), .Y(n595) );
  MUX2X1 U781 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1233), .Y(n594) );
  MUX2X1 U782 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1233), .Y(n598) );
  MUX2X1 U783 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1233), .Y(n597) );
  MUX2X1 U784 ( .B(n596), .A(n593), .S(n1193), .Y(n600) );
  MUX2X1 U785 ( .B(n599), .A(n584), .S(n1190), .Y(n1187) );
  MUX2X1 U786 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1233), .Y(n604) );
  MUX2X1 U787 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1233), .Y(n603) );
  MUX2X1 U788 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1233), .Y(n607) );
  MUX2X1 U789 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1233), .Y(n606) );
  MUX2X1 U790 ( .B(n605), .A(n602), .S(n1195), .Y(n616) );
  MUX2X1 U791 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1233), .Y(n610) );
  MUX2X1 U792 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1233), .Y(n609) );
  MUX2X1 U793 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1233), .Y(n613) );
  MUX2X1 U794 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1233), .Y(n612) );
  MUX2X1 U795 ( .B(n611), .A(n608), .S(n1193), .Y(n615) );
  MUX2X1 U796 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1234), .Y(n619) );
  MUX2X1 U797 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1234), .Y(n618) );
  MUX2X1 U798 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1234), .Y(n622) );
  MUX2X1 U799 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1234), .Y(n621) );
  MUX2X1 U800 ( .B(n620), .A(n617), .S(n1193), .Y(n631) );
  MUX2X1 U801 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1234), .Y(n625) );
  MUX2X1 U802 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1234), .Y(n624) );
  MUX2X1 U803 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1234), .Y(n628) );
  MUX2X1 U804 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1234), .Y(n627) );
  MUX2X1 U805 ( .B(n626), .A(n623), .S(n1193), .Y(n630) );
  MUX2X1 U806 ( .B(n629), .A(n614), .S(n1190), .Y(n1188) );
  MUX2X1 U807 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1234), .Y(n634) );
  MUX2X1 U808 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1234), .Y(n633) );
  MUX2X1 U809 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1234), .Y(n637) );
  MUX2X1 U810 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1234), .Y(n636) );
  MUX2X1 U811 ( .B(n635), .A(n632), .S(n1193), .Y(n646) );
  MUX2X1 U812 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1235), .Y(n640) );
  MUX2X1 U813 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1235), .Y(n639) );
  MUX2X1 U814 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1235), .Y(n643) );
  MUX2X1 U815 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1235), .Y(n642) );
  MUX2X1 U816 ( .B(n641), .A(n638), .S(n1193), .Y(n645) );
  MUX2X1 U817 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1235), .Y(n649) );
  MUX2X1 U818 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1235), .Y(n648) );
  MUX2X1 U819 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1235), .Y(n1164) );
  MUX2X1 U820 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1235), .Y(n1163) );
  MUX2X1 U821 ( .B(n650), .A(n647), .S(n1193), .Y(n1173) );
  MUX2X1 U822 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1235), .Y(n1167) );
  MUX2X1 U823 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1235), .Y(n1166) );
  MUX2X1 U824 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1235), .Y(n1170) );
  MUX2X1 U825 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1235), .Y(n1169) );
  MUX2X1 U826 ( .B(n1168), .A(n1165), .S(n1193), .Y(n1172) );
  MUX2X1 U827 ( .B(n1171), .A(n644), .S(n1190), .Y(n1189) );
  INVX4 U828 ( .A(n1310), .Y(n1308) );
  INVX1 U829 ( .A(n93), .Y(n1311) );
  AND2X1 U830 ( .A(n1344), .B(N23), .Y(n1239) );
  INVX1 U831 ( .A(N10), .Y(n1346) );
  INVX8 U832 ( .A(n1310), .Y(n1309) );
  INVX8 U833 ( .A(n19), .Y(n1312) );
  INVX8 U834 ( .A(n19), .Y(n1313) );
  INVX8 U835 ( .A(n20), .Y(n1314) );
  INVX8 U836 ( .A(n20), .Y(n1315) );
  INVX8 U837 ( .A(n21), .Y(n1316) );
  INVX8 U838 ( .A(n21), .Y(n1317) );
  INVX8 U839 ( .A(n22), .Y(n1318) );
  INVX8 U840 ( .A(n22), .Y(n1319) );
  INVX8 U841 ( .A(n23), .Y(n1320) );
  INVX8 U842 ( .A(n23), .Y(n1321) );
  INVX8 U843 ( .A(n24), .Y(n1322) );
  INVX8 U844 ( .A(n24), .Y(n1323) );
  INVX8 U845 ( .A(n25), .Y(n1324) );
  INVX8 U846 ( .A(n25), .Y(n1325) );
  INVX8 U847 ( .A(n26), .Y(n1326) );
  INVX8 U848 ( .A(n26), .Y(n1327) );
  INVX8 U849 ( .A(n27), .Y(n1328) );
  INVX8 U850 ( .A(n27), .Y(n1329) );
  INVX8 U851 ( .A(n28), .Y(n1330) );
  INVX8 U852 ( .A(n28), .Y(n1331) );
  INVX8 U853 ( .A(n29), .Y(n1332) );
  INVX8 U854 ( .A(n29), .Y(n1333) );
  INVX8 U855 ( .A(n94), .Y(n1334) );
  INVX8 U856 ( .A(n94), .Y(n1335) );
  INVX8 U857 ( .A(n95), .Y(n1336) );
  INVX8 U858 ( .A(n95), .Y(n1337) );
  INVX8 U859 ( .A(n96), .Y(n1338) );
  INVX8 U860 ( .A(n96), .Y(n1339) );
  INVX8 U861 ( .A(n97), .Y(n1340) );
  INVX8 U862 ( .A(n97), .Y(n1341) );
  INVX8 U863 ( .A(n98), .Y(n1342) );
  INVX8 U864 ( .A(n98), .Y(n1343) );
  AND2X2 U865 ( .A(n18), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U866 ( .A(N31), .B(n38), .Y(\data_out<1> ) );
  AND2X2 U867 ( .A(n17), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U868 ( .A(n18), .B(N29), .Y(\data_out<3> ) );
  AND2X2 U869 ( .A(n18), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U870 ( .A(n17), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U871 ( .A(N26), .B(n18), .Y(\data_out<6> ) );
  AND2X2 U872 ( .A(N25), .B(n38), .Y(\data_out<7> ) );
  AND2X2 U873 ( .A(N24), .B(n17), .Y(\data_out<8> ) );
  AND2X2 U874 ( .A(n1238), .B(n1239), .Y(\data_out<9> ) );
  AND2X2 U875 ( .A(n17), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U876 ( .A(n38), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U877 ( .A(n18), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U878 ( .A(N19), .B(n38), .Y(\data_out<13> ) );
  AND2X2 U879 ( .A(N18), .B(n38), .Y(\data_out<14> ) );
  AND2X2 U880 ( .A(n17), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U881 ( .A(\mem<31><0> ), .B(n1242), .Y(n1354) );
  OAI21X1 U882 ( .A(n1241), .B(n1312), .C(n1354), .Y(n2392) );
  NAND2X1 U883 ( .A(\mem<31><1> ), .B(n4), .Y(n1355) );
  OAI21X1 U884 ( .A(n1315), .B(n1240), .C(n1355), .Y(n2391) );
  NAND2X1 U885 ( .A(\mem<31><2> ), .B(n13), .Y(n1356) );
  OAI21X1 U886 ( .A(n1317), .B(n1240), .C(n1356), .Y(n2390) );
  NAND2X1 U887 ( .A(\mem<31><3> ), .B(n1243), .Y(n1357) );
  OAI21X1 U888 ( .A(n1318), .B(n1240), .C(n1357), .Y(n2389) );
  NAND2X1 U889 ( .A(\mem<31><4> ), .B(n4), .Y(n1358) );
  OAI21X1 U890 ( .A(n1321), .B(n1240), .C(n1358), .Y(n2388) );
  NAND2X1 U891 ( .A(\mem<31><5> ), .B(n1242), .Y(n1359) );
  OAI21X1 U892 ( .A(n1323), .B(n1240), .C(n1359), .Y(n2387) );
  NAND2X1 U893 ( .A(\mem<31><6> ), .B(n1242), .Y(n1360) );
  OAI21X1 U894 ( .A(n1324), .B(n1240), .C(n1360), .Y(n2386) );
  NAND2X1 U895 ( .A(\mem<31><7> ), .B(n1243), .Y(n1361) );
  OAI21X1 U896 ( .A(n1327), .B(n1240), .C(n1361), .Y(n2385) );
  NAND2X1 U897 ( .A(\mem<31><8> ), .B(n1243), .Y(n1362) );
  OAI21X1 U898 ( .A(n1329), .B(n1240), .C(n1362), .Y(n2384) );
  NAND2X1 U899 ( .A(\mem<31><9> ), .B(n13), .Y(n1363) );
  OAI21X1 U900 ( .A(n1331), .B(n1241), .C(n1363), .Y(n2383) );
  NAND2X1 U901 ( .A(\mem<31><10> ), .B(n13), .Y(n1364) );
  OAI21X1 U902 ( .A(n1333), .B(n1241), .C(n1364), .Y(n2382) );
  NAND2X1 U903 ( .A(\mem<31><11> ), .B(n13), .Y(n1365) );
  OAI21X1 U904 ( .A(n1335), .B(n1241), .C(n1365), .Y(n2381) );
  NAND2X1 U905 ( .A(\mem<31><12> ), .B(n1243), .Y(n1366) );
  OAI21X1 U906 ( .A(n1337), .B(n1241), .C(n1366), .Y(n2380) );
  NAND2X1 U907 ( .A(\mem<31><13> ), .B(n4), .Y(n1367) );
  OAI21X1 U908 ( .A(n1339), .B(n1241), .C(n1367), .Y(n2379) );
  NAND2X1 U909 ( .A(\mem<31><14> ), .B(n1242), .Y(n1368) );
  OAI21X1 U910 ( .A(n1341), .B(n1241), .C(n1368), .Y(n2378) );
  NAND2X1 U911 ( .A(\mem<31><15> ), .B(n4), .Y(n1369) );
  OAI21X1 U912 ( .A(n1343), .B(n1241), .C(n1369), .Y(n2377) );
  NAND2X1 U913 ( .A(\mem<30><0> ), .B(n57), .Y(n1370) );
  OAI21X1 U914 ( .A(n1244), .B(n1312), .C(n1370), .Y(n2376) );
  NAND2X1 U915 ( .A(\mem<30><1> ), .B(n57), .Y(n1371) );
  OAI21X1 U916 ( .A(n1244), .B(n1315), .C(n1371), .Y(n2375) );
  NAND2X1 U917 ( .A(\mem<30><2> ), .B(n57), .Y(n1372) );
  OAI21X1 U918 ( .A(n1244), .B(n1317), .C(n1372), .Y(n2374) );
  NAND2X1 U919 ( .A(\mem<30><3> ), .B(n57), .Y(n1373) );
  OAI21X1 U920 ( .A(n1244), .B(n1318), .C(n1373), .Y(n2373) );
  NAND2X1 U921 ( .A(\mem<30><4> ), .B(n57), .Y(n1374) );
  OAI21X1 U922 ( .A(n1244), .B(n1321), .C(n1374), .Y(n2372) );
  NAND2X1 U923 ( .A(\mem<30><5> ), .B(n57), .Y(n1375) );
  OAI21X1 U924 ( .A(n1244), .B(n1323), .C(n1375), .Y(n2371) );
  NAND2X1 U925 ( .A(\mem<30><6> ), .B(n57), .Y(n1376) );
  OAI21X1 U926 ( .A(n1244), .B(n1324), .C(n1376), .Y(n2370) );
  NAND2X1 U927 ( .A(\mem<30><7> ), .B(n57), .Y(n1377) );
  OAI21X1 U928 ( .A(n1244), .B(n1327), .C(n1377), .Y(n2369) );
  NAND2X1 U929 ( .A(\mem<30><8> ), .B(n57), .Y(n1378) );
  OAI21X1 U930 ( .A(n1245), .B(n1328), .C(n1378), .Y(n2368) );
  NAND2X1 U931 ( .A(\mem<30><9> ), .B(n57), .Y(n1379) );
  OAI21X1 U932 ( .A(n1245), .B(n1330), .C(n1379), .Y(n2367) );
  NAND2X1 U933 ( .A(\mem<30><10> ), .B(n57), .Y(n1380) );
  OAI21X1 U934 ( .A(n1245), .B(n1332), .C(n1380), .Y(n2366) );
  NAND2X1 U935 ( .A(\mem<30><11> ), .B(n57), .Y(n1381) );
  OAI21X1 U936 ( .A(n1245), .B(n1334), .C(n1381), .Y(n2365) );
  NAND2X1 U937 ( .A(\mem<30><12> ), .B(n57), .Y(n1382) );
  OAI21X1 U938 ( .A(n1245), .B(n1336), .C(n1382), .Y(n2364) );
  NAND2X1 U939 ( .A(\mem<30><13> ), .B(n57), .Y(n1383) );
  OAI21X1 U940 ( .A(n1245), .B(n1338), .C(n1383), .Y(n2363) );
  NAND2X1 U941 ( .A(\mem<30><14> ), .B(n57), .Y(n1384) );
  OAI21X1 U942 ( .A(n1245), .B(n1340), .C(n1384), .Y(n2362) );
  NAND2X1 U943 ( .A(\mem<30><15> ), .B(n57), .Y(n1385) );
  OAI21X1 U944 ( .A(n1245), .B(n1342), .C(n1385), .Y(n2361) );
  NAND3X1 U945 ( .A(n1345), .B(n1349), .C(n1348), .Y(n1386) );
  NAND2X1 U946 ( .A(\mem<29><0> ), .B(n59), .Y(n1387) );
  OAI21X1 U947 ( .A(n1246), .B(n1312), .C(n1387), .Y(n2360) );
  NAND2X1 U948 ( .A(\mem<29><1> ), .B(n59), .Y(n1388) );
  OAI21X1 U949 ( .A(n1246), .B(n1314), .C(n1388), .Y(n2359) );
  NAND2X1 U950 ( .A(\mem<29><2> ), .B(n59), .Y(n1389) );
  OAI21X1 U951 ( .A(n1246), .B(n1316), .C(n1389), .Y(n2358) );
  NAND2X1 U952 ( .A(\mem<29><3> ), .B(n59), .Y(n1390) );
  OAI21X1 U953 ( .A(n1246), .B(n1319), .C(n1390), .Y(n2357) );
  NAND2X1 U954 ( .A(\mem<29><4> ), .B(n59), .Y(n1391) );
  OAI21X1 U955 ( .A(n1246), .B(n1320), .C(n1391), .Y(n2356) );
  NAND2X1 U956 ( .A(\mem<29><5> ), .B(n59), .Y(n1392) );
  OAI21X1 U957 ( .A(n1246), .B(n1322), .C(n1392), .Y(n2355) );
  NAND2X1 U958 ( .A(\mem<29><6> ), .B(n59), .Y(n1393) );
  OAI21X1 U959 ( .A(n1246), .B(n1325), .C(n1393), .Y(n2354) );
  NAND2X1 U960 ( .A(\mem<29><7> ), .B(n59), .Y(n1394) );
  OAI21X1 U961 ( .A(n1246), .B(n1327), .C(n1394), .Y(n2353) );
  NAND2X1 U962 ( .A(\mem<29><8> ), .B(n59), .Y(n1395) );
  OAI21X1 U963 ( .A(n1247), .B(n1329), .C(n1395), .Y(n2352) );
  NAND2X1 U964 ( .A(\mem<29><9> ), .B(n59), .Y(n1396) );
  OAI21X1 U965 ( .A(n1247), .B(n1331), .C(n1396), .Y(n2351) );
  NAND2X1 U966 ( .A(\mem<29><10> ), .B(n59), .Y(n1397) );
  OAI21X1 U967 ( .A(n1247), .B(n1333), .C(n1397), .Y(n2350) );
  NAND2X1 U968 ( .A(\mem<29><11> ), .B(n59), .Y(n1398) );
  OAI21X1 U969 ( .A(n1247), .B(n1335), .C(n1398), .Y(n2349) );
  NAND2X1 U970 ( .A(\mem<29><12> ), .B(n59), .Y(n1399) );
  OAI21X1 U971 ( .A(n1247), .B(n1337), .C(n1399), .Y(n2348) );
  NAND2X1 U972 ( .A(\mem<29><13> ), .B(n59), .Y(n1400) );
  OAI21X1 U973 ( .A(n1247), .B(n1339), .C(n1400), .Y(n2347) );
  NAND2X1 U974 ( .A(\mem<29><14> ), .B(n59), .Y(n1401) );
  OAI21X1 U975 ( .A(n1247), .B(n1341), .C(n1401), .Y(n2346) );
  NAND2X1 U976 ( .A(\mem<29><15> ), .B(n59), .Y(n1402) );
  OAI21X1 U977 ( .A(n1247), .B(n1343), .C(n1402), .Y(n2345) );
  NAND3X1 U978 ( .A(n1349), .B(n1348), .C(n1346), .Y(n1403) );
  NAND2X1 U979 ( .A(\mem<28><0> ), .B(n61), .Y(n1404) );
  OAI21X1 U980 ( .A(n1248), .B(n1312), .C(n1404), .Y(n2344) );
  NAND2X1 U981 ( .A(\mem<28><1> ), .B(n61), .Y(n1405) );
  OAI21X1 U982 ( .A(n1248), .B(n1315), .C(n1405), .Y(n2343) );
  NAND2X1 U983 ( .A(\mem<28><2> ), .B(n61), .Y(n1406) );
  OAI21X1 U984 ( .A(n1248), .B(n1317), .C(n1406), .Y(n2342) );
  NAND2X1 U985 ( .A(\mem<28><3> ), .B(n61), .Y(n1407) );
  OAI21X1 U986 ( .A(n1248), .B(n1318), .C(n1407), .Y(n2341) );
  NAND2X1 U987 ( .A(\mem<28><4> ), .B(n61), .Y(n1408) );
  OAI21X1 U988 ( .A(n1248), .B(n1321), .C(n1408), .Y(n2340) );
  NAND2X1 U989 ( .A(\mem<28><5> ), .B(n61), .Y(n1409) );
  OAI21X1 U990 ( .A(n1248), .B(n1323), .C(n1409), .Y(n2339) );
  NAND2X1 U991 ( .A(\mem<28><6> ), .B(n61), .Y(n1410) );
  OAI21X1 U992 ( .A(n1248), .B(n1324), .C(n1410), .Y(n2338) );
  NAND2X1 U993 ( .A(\mem<28><7> ), .B(n61), .Y(n1411) );
  OAI21X1 U994 ( .A(n1248), .B(n1327), .C(n1411), .Y(n2337) );
  NAND2X1 U995 ( .A(\mem<28><8> ), .B(n61), .Y(n1412) );
  OAI21X1 U996 ( .A(n1249), .B(n1328), .C(n1412), .Y(n2336) );
  NAND2X1 U997 ( .A(\mem<28><9> ), .B(n61), .Y(n1413) );
  OAI21X1 U998 ( .A(n1249), .B(n1330), .C(n1413), .Y(n2335) );
  NAND2X1 U999 ( .A(\mem<28><10> ), .B(n61), .Y(n1414) );
  OAI21X1 U1000 ( .A(n1249), .B(n1332), .C(n1414), .Y(n2334) );
  NAND2X1 U1001 ( .A(\mem<28><11> ), .B(n61), .Y(n1415) );
  OAI21X1 U1002 ( .A(n1249), .B(n1334), .C(n1415), .Y(n2333) );
  NAND2X1 U1003 ( .A(\mem<28><12> ), .B(n61), .Y(n1416) );
  OAI21X1 U1004 ( .A(n1249), .B(n1336), .C(n1416), .Y(n2332) );
  NAND2X1 U1005 ( .A(\mem<28><13> ), .B(n61), .Y(n1417) );
  OAI21X1 U1006 ( .A(n1249), .B(n1338), .C(n1417), .Y(n2331) );
  NAND2X1 U1007 ( .A(\mem<28><14> ), .B(n61), .Y(n1418) );
  OAI21X1 U1008 ( .A(n1249), .B(n1340), .C(n1418), .Y(n2330) );
  NAND2X1 U1009 ( .A(\mem<28><15> ), .B(n61), .Y(n1419) );
  OAI21X1 U1010 ( .A(n1249), .B(n1342), .C(n1419), .Y(n2329) );
  NAND3X1 U1011 ( .A(n1345), .B(n1347), .C(n1350), .Y(n1420) );
  NAND2X1 U1012 ( .A(\mem<27><0> ), .B(n63), .Y(n1421) );
  OAI21X1 U1013 ( .A(n1250), .B(n1312), .C(n1421), .Y(n2328) );
  NAND2X1 U1014 ( .A(\mem<27><1> ), .B(n63), .Y(n1422) );
  OAI21X1 U1015 ( .A(n1250), .B(n1314), .C(n1422), .Y(n2327) );
  NAND2X1 U1016 ( .A(\mem<27><2> ), .B(n63), .Y(n1423) );
  OAI21X1 U1017 ( .A(n1250), .B(n1316), .C(n1423), .Y(n2326) );
  NAND2X1 U1018 ( .A(\mem<27><3> ), .B(n63), .Y(n1424) );
  OAI21X1 U1019 ( .A(n1250), .B(n1319), .C(n1424), .Y(n2325) );
  NAND2X1 U1020 ( .A(\mem<27><4> ), .B(n63), .Y(n1425) );
  OAI21X1 U1021 ( .A(n1250), .B(n1320), .C(n1425), .Y(n2324) );
  NAND2X1 U1022 ( .A(\mem<27><5> ), .B(n63), .Y(n1426) );
  OAI21X1 U1023 ( .A(n1250), .B(n1322), .C(n1426), .Y(n2323) );
  NAND2X1 U1024 ( .A(\mem<27><6> ), .B(n63), .Y(n1427) );
  OAI21X1 U1025 ( .A(n1250), .B(n1325), .C(n1427), .Y(n2322) );
  NAND2X1 U1026 ( .A(\mem<27><7> ), .B(n63), .Y(n1428) );
  OAI21X1 U1027 ( .A(n1250), .B(n1327), .C(n1428), .Y(n2321) );
  NAND2X1 U1028 ( .A(\mem<27><8> ), .B(n63), .Y(n1429) );
  OAI21X1 U1029 ( .A(n1251), .B(n1329), .C(n1429), .Y(n2320) );
  NAND2X1 U1030 ( .A(\mem<27><9> ), .B(n63), .Y(n1430) );
  OAI21X1 U1031 ( .A(n1251), .B(n1331), .C(n1430), .Y(n2319) );
  NAND2X1 U1032 ( .A(\mem<27><10> ), .B(n63), .Y(n1431) );
  OAI21X1 U1033 ( .A(n1251), .B(n1333), .C(n1431), .Y(n2318) );
  NAND2X1 U1034 ( .A(\mem<27><11> ), .B(n63), .Y(n1432) );
  OAI21X1 U1035 ( .A(n1251), .B(n1335), .C(n1432), .Y(n2317) );
  NAND2X1 U1036 ( .A(\mem<27><12> ), .B(n63), .Y(n1433) );
  OAI21X1 U1037 ( .A(n1251), .B(n1337), .C(n1433), .Y(n2316) );
  NAND2X1 U1038 ( .A(\mem<27><13> ), .B(n63), .Y(n1434) );
  OAI21X1 U1039 ( .A(n1251), .B(n1339), .C(n1434), .Y(n2315) );
  NAND2X1 U1040 ( .A(\mem<27><14> ), .B(n63), .Y(n1435) );
  OAI21X1 U1041 ( .A(n1251), .B(n1341), .C(n1435), .Y(n2314) );
  NAND2X1 U1042 ( .A(\mem<27><15> ), .B(n63), .Y(n1436) );
  OAI21X1 U1043 ( .A(n1251), .B(n1343), .C(n1436), .Y(n2313) );
  NAND3X1 U1044 ( .A(n1350), .B(n1347), .C(n1346), .Y(n1437) );
  NAND2X1 U1045 ( .A(\mem<26><0> ), .B(n65), .Y(n1438) );
  OAI21X1 U1046 ( .A(n1252), .B(n1312), .C(n1438), .Y(n2312) );
  NAND2X1 U1047 ( .A(\mem<26><1> ), .B(n65), .Y(n1439) );
  OAI21X1 U1048 ( .A(n1252), .B(n1315), .C(n1439), .Y(n2311) );
  NAND2X1 U1049 ( .A(\mem<26><2> ), .B(n65), .Y(n1440) );
  OAI21X1 U1050 ( .A(n1252), .B(n1317), .C(n1440), .Y(n2310) );
  NAND2X1 U1051 ( .A(\mem<26><3> ), .B(n65), .Y(n1441) );
  OAI21X1 U1052 ( .A(n1252), .B(n1318), .C(n1441), .Y(n2309) );
  NAND2X1 U1053 ( .A(\mem<26><4> ), .B(n65), .Y(n1442) );
  OAI21X1 U1054 ( .A(n1252), .B(n1321), .C(n1442), .Y(n2308) );
  NAND2X1 U1055 ( .A(\mem<26><5> ), .B(n65), .Y(n1443) );
  OAI21X1 U1056 ( .A(n1252), .B(n1323), .C(n1443), .Y(n2307) );
  NAND2X1 U1057 ( .A(\mem<26><6> ), .B(n65), .Y(n1444) );
  OAI21X1 U1058 ( .A(n1252), .B(n1324), .C(n1444), .Y(n2306) );
  NAND2X1 U1059 ( .A(\mem<26><7> ), .B(n65), .Y(n1445) );
  OAI21X1 U1060 ( .A(n1252), .B(n1327), .C(n1445), .Y(n2305) );
  NAND2X1 U1061 ( .A(\mem<26><8> ), .B(n65), .Y(n1446) );
  OAI21X1 U1062 ( .A(n1253), .B(n1328), .C(n1446), .Y(n2304) );
  NAND2X1 U1063 ( .A(\mem<26><9> ), .B(n65), .Y(n1447) );
  OAI21X1 U1064 ( .A(n1253), .B(n1330), .C(n1447), .Y(n2303) );
  NAND2X1 U1065 ( .A(\mem<26><10> ), .B(n65), .Y(n1448) );
  OAI21X1 U1066 ( .A(n1253), .B(n1332), .C(n1448), .Y(n2302) );
  NAND2X1 U1067 ( .A(\mem<26><11> ), .B(n65), .Y(n1449) );
  OAI21X1 U1068 ( .A(n1253), .B(n1334), .C(n1449), .Y(n2301) );
  NAND2X1 U1069 ( .A(\mem<26><12> ), .B(n65), .Y(n1450) );
  OAI21X1 U1070 ( .A(n1253), .B(n1336), .C(n1450), .Y(n2300) );
  NAND2X1 U1071 ( .A(\mem<26><13> ), .B(n65), .Y(n1451) );
  OAI21X1 U1072 ( .A(n1253), .B(n1338), .C(n1451), .Y(n2299) );
  NAND2X1 U1073 ( .A(\mem<26><14> ), .B(n65), .Y(n1452) );
  OAI21X1 U1074 ( .A(n1253), .B(n1340), .C(n1452), .Y(n2298) );
  NAND2X1 U1075 ( .A(\mem<26><15> ), .B(n65), .Y(n1453) );
  OAI21X1 U1076 ( .A(n1253), .B(n1342), .C(n1453), .Y(n2297) );
  NAND3X1 U1077 ( .A(n1345), .B(n1350), .C(n1348), .Y(n1454) );
  NAND2X1 U1078 ( .A(\mem<25><0> ), .B(n67), .Y(n1455) );
  OAI21X1 U1079 ( .A(n1254), .B(n1312), .C(n1455), .Y(n2296) );
  NAND2X1 U1080 ( .A(\mem<25><1> ), .B(n67), .Y(n1456) );
  OAI21X1 U1081 ( .A(n1254), .B(n1314), .C(n1456), .Y(n2295) );
  NAND2X1 U1082 ( .A(\mem<25><2> ), .B(n67), .Y(n1457) );
  OAI21X1 U1083 ( .A(n1254), .B(n1316), .C(n1457), .Y(n2294) );
  NAND2X1 U1084 ( .A(\mem<25><3> ), .B(n67), .Y(n1458) );
  OAI21X1 U1085 ( .A(n1254), .B(n1319), .C(n1458), .Y(n2293) );
  NAND2X1 U1086 ( .A(\mem<25><4> ), .B(n67), .Y(n1459) );
  OAI21X1 U1087 ( .A(n1254), .B(n1320), .C(n1459), .Y(n2292) );
  NAND2X1 U1088 ( .A(\mem<25><5> ), .B(n67), .Y(n1460) );
  OAI21X1 U1089 ( .A(n1254), .B(n1322), .C(n1460), .Y(n2291) );
  NAND2X1 U1090 ( .A(\mem<25><6> ), .B(n67), .Y(n1461) );
  OAI21X1 U1091 ( .A(n1254), .B(n1325), .C(n1461), .Y(n2290) );
  NAND2X1 U1092 ( .A(\mem<25><7> ), .B(n67), .Y(n1462) );
  OAI21X1 U1093 ( .A(n1254), .B(n1327), .C(n1462), .Y(n2289) );
  NAND2X1 U1094 ( .A(\mem<25><8> ), .B(n67), .Y(n1463) );
  OAI21X1 U1095 ( .A(n1255), .B(n1329), .C(n1463), .Y(n2288) );
  NAND2X1 U1096 ( .A(\mem<25><9> ), .B(n67), .Y(n1464) );
  OAI21X1 U1097 ( .A(n1255), .B(n1331), .C(n1464), .Y(n2287) );
  NAND2X1 U1098 ( .A(\mem<25><10> ), .B(n67), .Y(n1465) );
  OAI21X1 U1099 ( .A(n1255), .B(n1333), .C(n1465), .Y(n2286) );
  NAND2X1 U1100 ( .A(\mem<25><11> ), .B(n67), .Y(n1466) );
  OAI21X1 U1101 ( .A(n1255), .B(n1335), .C(n1466), .Y(n2285) );
  NAND2X1 U1102 ( .A(\mem<25><12> ), .B(n67), .Y(n1467) );
  OAI21X1 U1103 ( .A(n1255), .B(n1337), .C(n1467), .Y(n2284) );
  NAND2X1 U1104 ( .A(\mem<25><13> ), .B(n67), .Y(n1468) );
  OAI21X1 U1105 ( .A(n1255), .B(n1339), .C(n1468), .Y(n2283) );
  NAND2X1 U1106 ( .A(\mem<25><14> ), .B(n67), .Y(n1469) );
  OAI21X1 U1107 ( .A(n1255), .B(n1341), .C(n1469), .Y(n2282) );
  NAND2X1 U1108 ( .A(\mem<25><15> ), .B(n67), .Y(n1470) );
  OAI21X1 U1109 ( .A(n1255), .B(n1343), .C(n1470), .Y(n2281) );
  NOR3X1 U1110 ( .A(n1345), .B(n1347), .C(n1349), .Y(n1864) );
  NAND2X1 U1111 ( .A(\mem<24><0> ), .B(n15), .Y(n1471) );
  OAI21X1 U1112 ( .A(n1256), .B(n1312), .C(n1471), .Y(n2280) );
  NAND2X1 U1113 ( .A(\mem<24><1> ), .B(n15), .Y(n1472) );
  OAI21X1 U1114 ( .A(n1256), .B(n1314), .C(n1472), .Y(n2279) );
  NAND2X1 U1115 ( .A(\mem<24><2> ), .B(n52), .Y(n1473) );
  OAI21X1 U1116 ( .A(n1256), .B(n1316), .C(n1473), .Y(n2278) );
  NAND2X1 U1117 ( .A(\mem<24><3> ), .B(n15), .Y(n1474) );
  OAI21X1 U1118 ( .A(n1256), .B(n1319), .C(n1474), .Y(n2277) );
  NAND2X1 U1119 ( .A(\mem<24><4> ), .B(n52), .Y(n1475) );
  OAI21X1 U1120 ( .A(n1256), .B(n1320), .C(n1475), .Y(n2276) );
  NAND2X1 U1121 ( .A(\mem<24><5> ), .B(n14), .Y(n1476) );
  OAI21X1 U1122 ( .A(n1256), .B(n1322), .C(n1476), .Y(n2275) );
  NAND2X1 U1123 ( .A(\mem<24><6> ), .B(n180), .Y(n1477) );
  OAI21X1 U1124 ( .A(n1256), .B(n1325), .C(n1477), .Y(n2274) );
  NAND2X1 U1125 ( .A(\mem<24><7> ), .B(n14), .Y(n1478) );
  OAI21X1 U1126 ( .A(n1256), .B(n1327), .C(n1478), .Y(n2273) );
  NAND2X1 U1127 ( .A(\mem<24><8> ), .B(n180), .Y(n1479) );
  OAI21X1 U1128 ( .A(n1256), .B(n1328), .C(n1479), .Y(n2272) );
  NAND2X1 U1129 ( .A(\mem<24><9> ), .B(n180), .Y(n1480) );
  OAI21X1 U1130 ( .A(n1256), .B(n1330), .C(n1480), .Y(n2271) );
  NAND2X1 U1131 ( .A(\mem<24><10> ), .B(n52), .Y(n1481) );
  OAI21X1 U1132 ( .A(n1256), .B(n1332), .C(n1481), .Y(n2270) );
  NAND2X1 U1133 ( .A(\mem<24><11> ), .B(n14), .Y(n1482) );
  OAI21X1 U1134 ( .A(n1256), .B(n1334), .C(n1482), .Y(n2269) );
  NAND2X1 U1135 ( .A(\mem<24><12> ), .B(n52), .Y(n1483) );
  OAI21X1 U1136 ( .A(n1256), .B(n1336), .C(n1483), .Y(n2268) );
  NAND2X1 U1137 ( .A(\mem<24><13> ), .B(n14), .Y(n1484) );
  OAI21X1 U1138 ( .A(n1256), .B(n1338), .C(n1484), .Y(n2267) );
  NAND2X1 U1139 ( .A(\mem<24><14> ), .B(n15), .Y(n1485) );
  OAI21X1 U1140 ( .A(n1256), .B(n1340), .C(n1485), .Y(n2266) );
  NAND2X1 U1141 ( .A(\mem<24><15> ), .B(n180), .Y(n1486) );
  OAI21X1 U1142 ( .A(n1256), .B(n1342), .C(n1486), .Y(n2265) );
  NAND2X1 U1143 ( .A(\mem<23><0> ), .B(n11), .Y(n1487) );
  OAI21X1 U1144 ( .A(n1257), .B(n1312), .C(n1487), .Y(n2264) );
  NAND2X1 U1145 ( .A(\mem<23><1> ), .B(n69), .Y(n1488) );
  OAI21X1 U1146 ( .A(n1257), .B(n1315), .C(n1488), .Y(n2263) );
  NAND2X1 U1147 ( .A(\mem<23><2> ), .B(n1259), .Y(n1489) );
  OAI21X1 U1148 ( .A(n1257), .B(n1317), .C(n1489), .Y(n2262) );
  NAND2X1 U1149 ( .A(\mem<23><3> ), .B(n11), .Y(n1490) );
  OAI21X1 U1150 ( .A(n1257), .B(n1319), .C(n1490), .Y(n2261) );
  NAND2X1 U1151 ( .A(\mem<23><4> ), .B(n12), .Y(n1491) );
  OAI21X1 U1152 ( .A(n1257), .B(n1321), .C(n1491), .Y(n2260) );
  NAND2X1 U1153 ( .A(\mem<23><5> ), .B(n12), .Y(n1492) );
  OAI21X1 U1154 ( .A(n1257), .B(n1323), .C(n1492), .Y(n2259) );
  NAND2X1 U1155 ( .A(\mem<23><6> ), .B(n11), .Y(n1493) );
  OAI21X1 U1156 ( .A(n1257), .B(n1325), .C(n1493), .Y(n2258) );
  NAND2X1 U1157 ( .A(\mem<23><7> ), .B(n11), .Y(n1494) );
  OAI21X1 U1158 ( .A(n1257), .B(n1327), .C(n1494), .Y(n2257) );
  NAND2X1 U1159 ( .A(\mem<23><8> ), .B(n1259), .Y(n1495) );
  OAI21X1 U1160 ( .A(n1258), .B(n1329), .C(n1495), .Y(n2256) );
  NAND2X1 U1161 ( .A(\mem<23><9> ), .B(n69), .Y(n1496) );
  OAI21X1 U1162 ( .A(n1258), .B(n1331), .C(n1496), .Y(n2255) );
  NAND2X1 U1163 ( .A(\mem<23><10> ), .B(n1259), .Y(n1497) );
  OAI21X1 U1164 ( .A(n1258), .B(n1333), .C(n1497), .Y(n2254) );
  NAND2X1 U1165 ( .A(\mem<23><11> ), .B(n12), .Y(n1498) );
  OAI21X1 U1166 ( .A(n1258), .B(n1335), .C(n1498), .Y(n2253) );
  NAND2X1 U1167 ( .A(\mem<23><12> ), .B(n69), .Y(n1499) );
  OAI21X1 U1168 ( .A(n1258), .B(n1337), .C(n1499), .Y(n2252) );
  NAND2X1 U1169 ( .A(\mem<23><13> ), .B(n12), .Y(n1500) );
  OAI21X1 U1170 ( .A(n1258), .B(n1339), .C(n1500), .Y(n2251) );
  NAND2X1 U1171 ( .A(\mem<23><14> ), .B(n1259), .Y(n1501) );
  OAI21X1 U1172 ( .A(n1258), .B(n1341), .C(n1501), .Y(n2250) );
  NAND2X1 U1173 ( .A(\mem<23><15> ), .B(n69), .Y(n1502) );
  OAI21X1 U1174 ( .A(n1258), .B(n1343), .C(n1502), .Y(n2249) );
  NAND2X1 U1175 ( .A(\mem<22><0> ), .B(n9), .Y(n1503) );
  OAI21X1 U1177 ( .A(n1260), .B(n1312), .C(n1503), .Y(n2248) );
  NAND2X1 U1178 ( .A(\mem<22><1> ), .B(n72), .Y(n1504) );
  OAI21X1 U1179 ( .A(n1260), .B(n1315), .C(n1504), .Y(n2247) );
  NAND2X1 U1180 ( .A(\mem<22><2> ), .B(n1262), .Y(n1505) );
  OAI21X1 U1181 ( .A(n1260), .B(n1317), .C(n1505), .Y(n2246) );
  NAND2X1 U1182 ( .A(\mem<22><3> ), .B(n9), .Y(n1506) );
  OAI21X1 U1183 ( .A(n1260), .B(n1319), .C(n1506), .Y(n2245) );
  NAND2X1 U1184 ( .A(\mem<22><4> ), .B(n10), .Y(n1507) );
  OAI21X1 U1185 ( .A(n1260), .B(n1321), .C(n1507), .Y(n2244) );
  NAND2X1 U1186 ( .A(\mem<22><5> ), .B(n10), .Y(n1508) );
  OAI21X1 U1187 ( .A(n1260), .B(n1323), .C(n1508), .Y(n2243) );
  NAND2X1 U1188 ( .A(\mem<22><6> ), .B(n9), .Y(n1509) );
  OAI21X1 U1189 ( .A(n1260), .B(n1325), .C(n1509), .Y(n2242) );
  NAND2X1 U1190 ( .A(\mem<22><7> ), .B(n9), .Y(n1510) );
  OAI21X1 U1191 ( .A(n1260), .B(n1327), .C(n1510), .Y(n2241) );
  NAND2X1 U1192 ( .A(\mem<22><8> ), .B(n1262), .Y(n1511) );
  OAI21X1 U1193 ( .A(n1261), .B(n1329), .C(n1511), .Y(n2240) );
  NAND2X1 U1194 ( .A(\mem<22><9> ), .B(n72), .Y(n1512) );
  OAI21X1 U1195 ( .A(n1261), .B(n1331), .C(n1512), .Y(n2239) );
  NAND2X1 U1196 ( .A(\mem<22><10> ), .B(n1262), .Y(n1513) );
  OAI21X1 U1197 ( .A(n1261), .B(n1333), .C(n1513), .Y(n2238) );
  NAND2X1 U1198 ( .A(\mem<22><11> ), .B(n10), .Y(n1514) );
  OAI21X1 U1199 ( .A(n1261), .B(n1335), .C(n1514), .Y(n2237) );
  NAND2X1 U1200 ( .A(\mem<22><12> ), .B(n72), .Y(n1515) );
  OAI21X1 U1201 ( .A(n1261), .B(n1337), .C(n1515), .Y(n2236) );
  NAND2X1 U1202 ( .A(\mem<22><13> ), .B(n10), .Y(n1516) );
  OAI21X1 U1203 ( .A(n1261), .B(n1339), .C(n1516), .Y(n2235) );
  NAND2X1 U1204 ( .A(\mem<22><14> ), .B(n1262), .Y(n1517) );
  OAI21X1 U1205 ( .A(n1261), .B(n1341), .C(n1517), .Y(n2234) );
  NAND2X1 U1206 ( .A(\mem<22><15> ), .B(n72), .Y(n1518) );
  OAI21X1 U1207 ( .A(n1261), .B(n1343), .C(n1518), .Y(n2233) );
  NAND2X1 U1208 ( .A(\mem<21><0> ), .B(n8), .Y(n1519) );
  OAI21X1 U1209 ( .A(n1263), .B(n1312), .C(n1519), .Y(n2232) );
  NAND2X1 U1210 ( .A(\mem<21><1> ), .B(n7), .Y(n1520) );
  OAI21X1 U1211 ( .A(n1263), .B(n1315), .C(n1520), .Y(n2231) );
  NAND2X1 U1212 ( .A(\mem<21><2> ), .B(n1265), .Y(n1521) );
  OAI21X1 U1213 ( .A(n1263), .B(n1317), .C(n1521), .Y(n2230) );
  NAND2X1 U1214 ( .A(\mem<21><3> ), .B(n7), .Y(n1522) );
  OAI21X1 U1215 ( .A(n1263), .B(n1319), .C(n1522), .Y(n2229) );
  NAND2X1 U1216 ( .A(\mem<21><4> ), .B(n7), .Y(n1523) );
  OAI21X1 U1217 ( .A(n1263), .B(n1321), .C(n1523), .Y(n2228) );
  NAND2X1 U1218 ( .A(\mem<21><5> ), .B(n8), .Y(n1524) );
  OAI21X1 U1219 ( .A(n1263), .B(n1323), .C(n1524), .Y(n2227) );
  NAND2X1 U1220 ( .A(\mem<21><6> ), .B(n1265), .Y(n1525) );
  OAI21X1 U1221 ( .A(n1263), .B(n1325), .C(n1525), .Y(n2226) );
  NAND2X1 U1222 ( .A(\mem<21><7> ), .B(n7), .Y(n1526) );
  OAI21X1 U1223 ( .A(n1263), .B(n1327), .C(n1526), .Y(n2225) );
  NAND2X1 U1224 ( .A(\mem<21><8> ), .B(n8), .Y(n1527) );
  OAI21X1 U1225 ( .A(n1264), .B(n1329), .C(n1527), .Y(n2224) );
  NAND2X1 U1226 ( .A(\mem<21><9> ), .B(n46), .Y(n1528) );
  OAI21X1 U1227 ( .A(n1264), .B(n1331), .C(n1528), .Y(n2223) );
  NAND2X1 U1228 ( .A(\mem<21><10> ), .B(n46), .Y(n1529) );
  OAI21X1 U1229 ( .A(n1264), .B(n1333), .C(n1529), .Y(n2222) );
  NAND2X1 U1230 ( .A(\mem<21><11> ), .B(n1265), .Y(n1530) );
  OAI21X1 U1231 ( .A(n1264), .B(n1335), .C(n1530), .Y(n2221) );
  NAND2X1 U1232 ( .A(\mem<21><12> ), .B(n1265), .Y(n1531) );
  OAI21X1 U1233 ( .A(n1264), .B(n1337), .C(n1531), .Y(n2220) );
  NAND2X1 U1234 ( .A(\mem<21><13> ), .B(n46), .Y(n1532) );
  OAI21X1 U1235 ( .A(n1264), .B(n1339), .C(n1532), .Y(n2219) );
  NAND2X1 U1236 ( .A(\mem<21><14> ), .B(n8), .Y(n1533) );
  OAI21X1 U1237 ( .A(n1264), .B(n1341), .C(n1533), .Y(n2218) );
  NAND2X1 U1238 ( .A(\mem<21><15> ), .B(n46), .Y(n1534) );
  OAI21X1 U1239 ( .A(n1264), .B(n1343), .C(n1534), .Y(n2217) );
  NAND2X1 U1240 ( .A(\mem<20><0> ), .B(n6), .Y(n1535) );
  OAI21X1 U1241 ( .A(n1266), .B(n1312), .C(n1535), .Y(n2216) );
  NAND2X1 U1242 ( .A(\mem<20><1> ), .B(n5), .Y(n1536) );
  OAI21X1 U1243 ( .A(n1266), .B(n1315), .C(n1536), .Y(n2215) );
  NAND2X1 U1244 ( .A(\mem<20><2> ), .B(n1268), .Y(n1537) );
  OAI21X1 U1245 ( .A(n1266), .B(n1317), .C(n1537), .Y(n2214) );
  NAND2X1 U1246 ( .A(\mem<20><3> ), .B(n5), .Y(n1538) );
  OAI21X1 U1247 ( .A(n1266), .B(n1319), .C(n1538), .Y(n2213) );
  NAND2X1 U1248 ( .A(\mem<20><4> ), .B(n5), .Y(n1539) );
  OAI21X1 U1249 ( .A(n1266), .B(n1321), .C(n1539), .Y(n2212) );
  NAND2X1 U1250 ( .A(\mem<20><5> ), .B(n6), .Y(n1540) );
  OAI21X1 U1251 ( .A(n1266), .B(n1323), .C(n1540), .Y(n2211) );
  NAND2X1 U1252 ( .A(\mem<20><6> ), .B(n1268), .Y(n1541) );
  OAI21X1 U1253 ( .A(n1266), .B(n1325), .C(n1541), .Y(n2210) );
  NAND2X1 U1254 ( .A(\mem<20><7> ), .B(n5), .Y(n1542) );
  OAI21X1 U1255 ( .A(n1266), .B(n1327), .C(n1542), .Y(n2209) );
  NAND2X1 U1256 ( .A(\mem<20><8> ), .B(n6), .Y(n1543) );
  OAI21X1 U1257 ( .A(n1267), .B(n1329), .C(n1543), .Y(n2208) );
  NAND2X1 U1258 ( .A(\mem<20><9> ), .B(n49), .Y(n1544) );
  OAI21X1 U1259 ( .A(n1267), .B(n1331), .C(n1544), .Y(n2207) );
  NAND2X1 U1260 ( .A(\mem<20><10> ), .B(n49), .Y(n1545) );
  OAI21X1 U1261 ( .A(n1267), .B(n1333), .C(n1545), .Y(n2206) );
  NAND2X1 U1262 ( .A(\mem<20><11> ), .B(n1268), .Y(n1546) );
  OAI21X1 U1263 ( .A(n1267), .B(n1335), .C(n1546), .Y(n2205) );
  NAND2X1 U1264 ( .A(\mem<20><12> ), .B(n1268), .Y(n1547) );
  OAI21X1 U1265 ( .A(n1267), .B(n1337), .C(n1547), .Y(n2204) );
  NAND2X1 U1266 ( .A(\mem<20><13> ), .B(n49), .Y(n1548) );
  OAI21X1 U1267 ( .A(n1267), .B(n1339), .C(n1548), .Y(n2203) );
  NAND2X1 U1268 ( .A(\mem<20><14> ), .B(n6), .Y(n1549) );
  OAI21X1 U1269 ( .A(n1267), .B(n1341), .C(n1549), .Y(n2202) );
  NAND2X1 U1270 ( .A(\mem<20><15> ), .B(n49), .Y(n1550) );
  OAI21X1 U1271 ( .A(n1267), .B(n1343), .C(n1550), .Y(n2201) );
  NAND2X1 U1272 ( .A(\mem<19><0> ), .B(n75), .Y(n1551) );
  OAI21X1 U1273 ( .A(n1269), .B(n1313), .C(n1551), .Y(n2200) );
  NAND2X1 U1274 ( .A(\mem<19><1> ), .B(n75), .Y(n1552) );
  OAI21X1 U1275 ( .A(n1269), .B(n1315), .C(n1552), .Y(n2199) );
  NAND2X1 U1276 ( .A(\mem<19><2> ), .B(n75), .Y(n1553) );
  OAI21X1 U1277 ( .A(n1269), .B(n1317), .C(n1553), .Y(n2198) );
  NAND2X1 U1278 ( .A(\mem<19><3> ), .B(n75), .Y(n1554) );
  OAI21X1 U1279 ( .A(n1269), .B(n1319), .C(n1554), .Y(n2197) );
  NAND2X1 U1280 ( .A(\mem<19><4> ), .B(n75), .Y(n1555) );
  OAI21X1 U1281 ( .A(n1269), .B(n1321), .C(n1555), .Y(n2196) );
  NAND2X1 U1282 ( .A(\mem<19><5> ), .B(n75), .Y(n1556) );
  OAI21X1 U1283 ( .A(n1269), .B(n1323), .C(n1556), .Y(n2195) );
  NAND2X1 U1284 ( .A(\mem<19><6> ), .B(n75), .Y(n1557) );
  OAI21X1 U1285 ( .A(n1269), .B(n1325), .C(n1557), .Y(n2194) );
  NAND2X1 U1286 ( .A(\mem<19><7> ), .B(n75), .Y(n1558) );
  OAI21X1 U1287 ( .A(n1269), .B(n1326), .C(n1558), .Y(n2193) );
  NAND2X1 U1288 ( .A(\mem<19><8> ), .B(n75), .Y(n1559) );
  OAI21X1 U1289 ( .A(n1270), .B(n1329), .C(n1559), .Y(n2192) );
  NAND2X1 U1290 ( .A(\mem<19><9> ), .B(n75), .Y(n1560) );
  OAI21X1 U1291 ( .A(n1270), .B(n1331), .C(n1560), .Y(n2191) );
  NAND2X1 U1292 ( .A(\mem<19><10> ), .B(n75), .Y(n1561) );
  OAI21X1 U1293 ( .A(n1270), .B(n1333), .C(n1561), .Y(n2190) );
  NAND2X1 U1294 ( .A(\mem<19><11> ), .B(n75), .Y(n1562) );
  OAI21X1 U1295 ( .A(n1270), .B(n1335), .C(n1562), .Y(n2189) );
  NAND2X1 U1296 ( .A(\mem<19><12> ), .B(n75), .Y(n1563) );
  OAI21X1 U1297 ( .A(n1270), .B(n1337), .C(n1563), .Y(n2188) );
  NAND2X1 U1298 ( .A(\mem<19><13> ), .B(n75), .Y(n1564) );
  OAI21X1 U1299 ( .A(n1270), .B(n1339), .C(n1564), .Y(n2187) );
  NAND2X1 U1300 ( .A(\mem<19><14> ), .B(n75), .Y(n1565) );
  OAI21X1 U1301 ( .A(n1270), .B(n1341), .C(n1565), .Y(n2186) );
  NAND2X1 U1302 ( .A(\mem<19><15> ), .B(n75), .Y(n1566) );
  OAI21X1 U1303 ( .A(n1270), .B(n1343), .C(n1566), .Y(n2185) );
  NAND2X1 U1304 ( .A(\mem<18><0> ), .B(n77), .Y(n1567) );
  OAI21X1 U1305 ( .A(n1271), .B(n1313), .C(n1567), .Y(n2184) );
  NAND2X1 U1306 ( .A(\mem<18><1> ), .B(n77), .Y(n1568) );
  OAI21X1 U1307 ( .A(n1271), .B(n1315), .C(n1568), .Y(n2183) );
  NAND2X1 U1308 ( .A(\mem<18><2> ), .B(n77), .Y(n1569) );
  OAI21X1 U1309 ( .A(n1271), .B(n1317), .C(n1569), .Y(n2182) );
  NAND2X1 U1310 ( .A(\mem<18><3> ), .B(n77), .Y(n1570) );
  OAI21X1 U1311 ( .A(n1271), .B(n1319), .C(n1570), .Y(n2181) );
  NAND2X1 U1312 ( .A(\mem<18><4> ), .B(n77), .Y(n1571) );
  OAI21X1 U1313 ( .A(n1271), .B(n1321), .C(n1571), .Y(n2180) );
  NAND2X1 U1314 ( .A(\mem<18><5> ), .B(n77), .Y(n1572) );
  OAI21X1 U1315 ( .A(n1271), .B(n1323), .C(n1572), .Y(n2179) );
  NAND2X1 U1316 ( .A(\mem<18><6> ), .B(n77), .Y(n1573) );
  OAI21X1 U1317 ( .A(n1271), .B(n1325), .C(n1573), .Y(n2178) );
  NAND2X1 U1318 ( .A(\mem<18><7> ), .B(n77), .Y(n1574) );
  OAI21X1 U1319 ( .A(n1271), .B(n1327), .C(n1574), .Y(n2177) );
  NAND2X1 U1320 ( .A(\mem<18><8> ), .B(n77), .Y(n1575) );
  OAI21X1 U1321 ( .A(n1272), .B(n1329), .C(n1575), .Y(n2176) );
  NAND2X1 U1322 ( .A(\mem<18><9> ), .B(n77), .Y(n1576) );
  OAI21X1 U1323 ( .A(n1272), .B(n1331), .C(n1576), .Y(n2175) );
  NAND2X1 U1324 ( .A(\mem<18><10> ), .B(n77), .Y(n1577) );
  OAI21X1 U1325 ( .A(n1272), .B(n1333), .C(n1577), .Y(n2174) );
  NAND2X1 U1326 ( .A(\mem<18><11> ), .B(n77), .Y(n1578) );
  OAI21X1 U1327 ( .A(n1272), .B(n1335), .C(n1578), .Y(n2173) );
  NAND2X1 U1328 ( .A(\mem<18><12> ), .B(n77), .Y(n1579) );
  OAI21X1 U1329 ( .A(n1272), .B(n1337), .C(n1579), .Y(n2172) );
  NAND2X1 U1330 ( .A(\mem<18><13> ), .B(n77), .Y(n1580) );
  OAI21X1 U1331 ( .A(n1272), .B(n1339), .C(n1580), .Y(n2171) );
  NAND2X1 U1332 ( .A(\mem<18><14> ), .B(n77), .Y(n1581) );
  OAI21X1 U1333 ( .A(n1272), .B(n1341), .C(n1581), .Y(n2170) );
  NAND2X1 U1334 ( .A(\mem<18><15> ), .B(n77), .Y(n1582) );
  OAI21X1 U1335 ( .A(n1272), .B(n1343), .C(n1582), .Y(n2169) );
  NAND2X1 U1336 ( .A(\mem<17><0> ), .B(n79), .Y(n1583) );
  OAI21X1 U1337 ( .A(n1273), .B(n1313), .C(n1583), .Y(n2168) );
  NAND2X1 U1338 ( .A(\mem<17><1> ), .B(n79), .Y(n1584) );
  OAI21X1 U1339 ( .A(n1273), .B(n1315), .C(n1584), .Y(n2167) );
  NAND2X1 U1340 ( .A(\mem<17><2> ), .B(n79), .Y(n1585) );
  OAI21X1 U1341 ( .A(n1273), .B(n1317), .C(n1585), .Y(n2166) );
  NAND2X1 U1342 ( .A(\mem<17><3> ), .B(n79), .Y(n1586) );
  OAI21X1 U1343 ( .A(n1273), .B(n1319), .C(n1586), .Y(n2165) );
  NAND2X1 U1344 ( .A(\mem<17><4> ), .B(n79), .Y(n1587) );
  OAI21X1 U1345 ( .A(n1273), .B(n1321), .C(n1587), .Y(n2164) );
  NAND2X1 U1346 ( .A(\mem<17><5> ), .B(n79), .Y(n1588) );
  OAI21X1 U1347 ( .A(n1273), .B(n1323), .C(n1588), .Y(n2163) );
  NAND2X1 U1348 ( .A(\mem<17><6> ), .B(n79), .Y(n1589) );
  OAI21X1 U1349 ( .A(n1273), .B(n1325), .C(n1589), .Y(n2162) );
  NAND2X1 U1350 ( .A(\mem<17><7> ), .B(n79), .Y(n1590) );
  OAI21X1 U1351 ( .A(n1273), .B(n1326), .C(n1590), .Y(n2161) );
  NAND2X1 U1352 ( .A(\mem<17><8> ), .B(n79), .Y(n1591) );
  OAI21X1 U1353 ( .A(n1274), .B(n1329), .C(n1591), .Y(n2160) );
  NAND2X1 U1354 ( .A(\mem<17><9> ), .B(n79), .Y(n1592) );
  OAI21X1 U1355 ( .A(n1274), .B(n1331), .C(n1592), .Y(n2159) );
  NAND2X1 U1356 ( .A(\mem<17><10> ), .B(n79), .Y(n1593) );
  OAI21X1 U1357 ( .A(n1274), .B(n1333), .C(n1593), .Y(n2158) );
  NAND2X1 U1358 ( .A(\mem<17><11> ), .B(n79), .Y(n1594) );
  OAI21X1 U1359 ( .A(n1274), .B(n1335), .C(n1594), .Y(n2157) );
  NAND2X1 U1360 ( .A(\mem<17><12> ), .B(n79), .Y(n1595) );
  OAI21X1 U1361 ( .A(n1274), .B(n1337), .C(n1595), .Y(n2156) );
  NAND2X1 U1362 ( .A(\mem<17><13> ), .B(n79), .Y(n1596) );
  OAI21X1 U1363 ( .A(n1274), .B(n1339), .C(n1596), .Y(n2155) );
  NAND2X1 U1364 ( .A(\mem<17><14> ), .B(n79), .Y(n1597) );
  OAI21X1 U1365 ( .A(n1274), .B(n1341), .C(n1597), .Y(n2154) );
  NAND2X1 U1366 ( .A(\mem<17><15> ), .B(n79), .Y(n1598) );
  OAI21X1 U1367 ( .A(n1274), .B(n1343), .C(n1598), .Y(n2153) );
  NAND2X1 U1368 ( .A(\mem<16><0> ), .B(n3), .Y(n1599) );
  OAI21X1 U1369 ( .A(n1275), .B(n1313), .C(n1599), .Y(n2152) );
  NAND2X1 U1370 ( .A(\mem<16><1> ), .B(n3), .Y(n1600) );
  OAI21X1 U1371 ( .A(n1275), .B(n1315), .C(n1600), .Y(n2151) );
  NAND2X1 U1372 ( .A(\mem<16><2> ), .B(n1276), .Y(n1601) );
  OAI21X1 U1373 ( .A(n1275), .B(n1317), .C(n1601), .Y(n2150) );
  NAND2X1 U1374 ( .A(\mem<16><3> ), .B(n1276), .Y(n1602) );
  OAI21X1 U1375 ( .A(n1275), .B(n1319), .C(n1602), .Y(n2149) );
  NAND2X1 U1376 ( .A(\mem<16><4> ), .B(n3), .Y(n1603) );
  OAI21X1 U1377 ( .A(n1275), .B(n1321), .C(n1603), .Y(n2148) );
  NAND2X1 U1378 ( .A(\mem<16><5> ), .B(n3), .Y(n1604) );
  OAI21X1 U1379 ( .A(n1275), .B(n1323), .C(n1604), .Y(n2147) );
  NAND2X1 U1380 ( .A(\mem<16><6> ), .B(n1276), .Y(n1605) );
  OAI21X1 U1381 ( .A(n1275), .B(n1325), .C(n1605), .Y(n2146) );
  NAND2X1 U1382 ( .A(\mem<16><7> ), .B(n1276), .Y(n1606) );
  OAI21X1 U1383 ( .A(n1275), .B(n1327), .C(n1606), .Y(n2145) );
  NAND2X1 U1384 ( .A(\mem<16><8> ), .B(n82), .Y(n1607) );
  OAI21X1 U1385 ( .A(n1275), .B(n1329), .C(n1607), .Y(n2144) );
  NAND2X1 U1386 ( .A(\mem<16><9> ), .B(n2), .Y(n1608) );
  OAI21X1 U1387 ( .A(n1275), .B(n1331), .C(n1608), .Y(n2143) );
  NAND2X1 U1388 ( .A(\mem<16><10> ), .B(n82), .Y(n1609) );
  OAI21X1 U1389 ( .A(n1275), .B(n1333), .C(n1609), .Y(n2142) );
  NAND2X1 U1390 ( .A(\mem<16><11> ), .B(n2), .Y(n1610) );
  OAI21X1 U1391 ( .A(n1275), .B(n1335), .C(n1610), .Y(n2141) );
  NAND2X1 U1392 ( .A(\mem<16><12> ), .B(n82), .Y(n1611) );
  OAI21X1 U1393 ( .A(n1275), .B(n1337), .C(n1611), .Y(n2140) );
  NAND2X1 U1394 ( .A(\mem<16><13> ), .B(n2), .Y(n1612) );
  OAI21X1 U1395 ( .A(n1275), .B(n1339), .C(n1612), .Y(n2139) );
  NAND2X1 U1396 ( .A(\mem<16><14> ), .B(n82), .Y(n1613) );
  OAI21X1 U1397 ( .A(n1275), .B(n1341), .C(n1613), .Y(n2138) );
  NAND2X1 U1398 ( .A(\mem<16><15> ), .B(n2), .Y(n1614) );
  OAI21X1 U1399 ( .A(n1275), .B(n1343), .C(n1614), .Y(n2137) );
  NAND3X1 U1400 ( .A(n1351), .B(n2393), .C(n1353), .Y(n1615) );
  NAND2X1 U1401 ( .A(\mem<15><0> ), .B(n84), .Y(n1616) );
  OAI21X1 U1402 ( .A(n1277), .B(n1313), .C(n1616), .Y(n2136) );
  NAND2X1 U1403 ( .A(\mem<15><1> ), .B(n84), .Y(n1617) );
  OAI21X1 U1404 ( .A(n1277), .B(n1315), .C(n1617), .Y(n2135) );
  NAND2X1 U1405 ( .A(\mem<15><2> ), .B(n84), .Y(n1618) );
  OAI21X1 U1406 ( .A(n1277), .B(n1317), .C(n1618), .Y(n2134) );
  NAND2X1 U1407 ( .A(\mem<15><3> ), .B(n84), .Y(n1619) );
  OAI21X1 U1408 ( .A(n1277), .B(n1319), .C(n1619), .Y(n2133) );
  NAND2X1 U1409 ( .A(\mem<15><4> ), .B(n84), .Y(n1620) );
  OAI21X1 U1410 ( .A(n1277), .B(n1321), .C(n1620), .Y(n2132) );
  NAND2X1 U1411 ( .A(\mem<15><5> ), .B(n84), .Y(n1621) );
  OAI21X1 U1412 ( .A(n1277), .B(n1323), .C(n1621), .Y(n2131) );
  NAND2X1 U1413 ( .A(\mem<15><6> ), .B(n84), .Y(n1622) );
  OAI21X1 U1414 ( .A(n1277), .B(n1325), .C(n1622), .Y(n2130) );
  NAND2X1 U1415 ( .A(\mem<15><7> ), .B(n84), .Y(n1623) );
  OAI21X1 U1416 ( .A(n1277), .B(n1327), .C(n1623), .Y(n2129) );
  NAND2X1 U1417 ( .A(\mem<15><8> ), .B(n84), .Y(n1624) );
  OAI21X1 U1418 ( .A(n1278), .B(n1329), .C(n1624), .Y(n2128) );
  NAND2X1 U1419 ( .A(\mem<15><9> ), .B(n84), .Y(n1625) );
  OAI21X1 U1420 ( .A(n1278), .B(n1331), .C(n1625), .Y(n2127) );
  NAND2X1 U1421 ( .A(\mem<15><10> ), .B(n84), .Y(n1626) );
  OAI21X1 U1422 ( .A(n1278), .B(n1333), .C(n1626), .Y(n2126) );
  NAND2X1 U1423 ( .A(\mem<15><11> ), .B(n84), .Y(n1627) );
  OAI21X1 U1424 ( .A(n1278), .B(n1335), .C(n1627), .Y(n2125) );
  NAND2X1 U1425 ( .A(\mem<15><12> ), .B(n84), .Y(n1628) );
  OAI21X1 U1426 ( .A(n1278), .B(n1337), .C(n1628), .Y(n2124) );
  NAND2X1 U1427 ( .A(\mem<15><13> ), .B(n84), .Y(n1629) );
  OAI21X1 U1428 ( .A(n1278), .B(n1339), .C(n1629), .Y(n2123) );
  NAND2X1 U1429 ( .A(\mem<15><14> ), .B(n84), .Y(n1630) );
  OAI21X1 U1430 ( .A(n1278), .B(n1341), .C(n1630), .Y(n2122) );
  NAND2X1 U1431 ( .A(\mem<15><15> ), .B(n84), .Y(n1631) );
  OAI21X1 U1432 ( .A(n1278), .B(n1343), .C(n1631), .Y(n2121) );
  NAND2X1 U1433 ( .A(\mem<14><0> ), .B(n86), .Y(n1632) );
  OAI21X1 U1434 ( .A(n1279), .B(n1313), .C(n1632), .Y(n2120) );
  NAND2X1 U1435 ( .A(\mem<14><1> ), .B(n86), .Y(n1633) );
  OAI21X1 U1436 ( .A(n1279), .B(n1315), .C(n1633), .Y(n2119) );
  NAND2X1 U1437 ( .A(\mem<14><2> ), .B(n86), .Y(n1634) );
  OAI21X1 U1438 ( .A(n1279), .B(n1317), .C(n1634), .Y(n2118) );
  NAND2X1 U1439 ( .A(\mem<14><3> ), .B(n86), .Y(n1635) );
  OAI21X1 U1440 ( .A(n1279), .B(n1319), .C(n1635), .Y(n2117) );
  NAND2X1 U1441 ( .A(\mem<14><4> ), .B(n86), .Y(n1636) );
  OAI21X1 U1442 ( .A(n1279), .B(n1321), .C(n1636), .Y(n2116) );
  NAND2X1 U1443 ( .A(\mem<14><5> ), .B(n86), .Y(n1637) );
  OAI21X1 U1444 ( .A(n1279), .B(n1323), .C(n1637), .Y(n2115) );
  NAND2X1 U1445 ( .A(\mem<14><6> ), .B(n86), .Y(n1638) );
  OAI21X1 U1446 ( .A(n1279), .B(n1325), .C(n1638), .Y(n2114) );
  NAND2X1 U1447 ( .A(\mem<14><7> ), .B(n86), .Y(n1639) );
  OAI21X1 U1448 ( .A(n1279), .B(n1326), .C(n1639), .Y(n2113) );
  NAND2X1 U1449 ( .A(\mem<14><8> ), .B(n86), .Y(n1640) );
  OAI21X1 U1450 ( .A(n1280), .B(n1329), .C(n1640), .Y(n2112) );
  NAND2X1 U1451 ( .A(\mem<14><9> ), .B(n86), .Y(n1641) );
  OAI21X1 U1452 ( .A(n1280), .B(n1331), .C(n1641), .Y(n2111) );
  NAND2X1 U1453 ( .A(\mem<14><10> ), .B(n86), .Y(n1642) );
  OAI21X1 U1454 ( .A(n1280), .B(n1333), .C(n1642), .Y(n2110) );
  NAND2X1 U1455 ( .A(\mem<14><11> ), .B(n86), .Y(n1643) );
  OAI21X1 U1456 ( .A(n1280), .B(n1335), .C(n1643), .Y(n2109) );
  NAND2X1 U1457 ( .A(\mem<14><12> ), .B(n86), .Y(n1644) );
  OAI21X1 U1458 ( .A(n1280), .B(n1337), .C(n1644), .Y(n2108) );
  NAND2X1 U1459 ( .A(\mem<14><13> ), .B(n86), .Y(n1645) );
  OAI21X1 U1460 ( .A(n1280), .B(n1339), .C(n1645), .Y(n2107) );
  NAND2X1 U1461 ( .A(\mem<14><14> ), .B(n86), .Y(n1646) );
  OAI21X1 U1462 ( .A(n1280), .B(n1341), .C(n1646), .Y(n2106) );
  NAND2X1 U1463 ( .A(\mem<14><15> ), .B(n86), .Y(n1647) );
  OAI21X1 U1464 ( .A(n1280), .B(n1343), .C(n1647), .Y(n2105) );
  NAND2X1 U1465 ( .A(\mem<13><0> ), .B(n88), .Y(n1648) );
  OAI21X1 U1466 ( .A(n1281), .B(n1313), .C(n1648), .Y(n2104) );
  NAND2X1 U1467 ( .A(\mem<13><1> ), .B(n88), .Y(n1649) );
  OAI21X1 U1468 ( .A(n1281), .B(n1315), .C(n1649), .Y(n2103) );
  NAND2X1 U1469 ( .A(\mem<13><2> ), .B(n88), .Y(n1650) );
  OAI21X1 U1470 ( .A(n1281), .B(n1317), .C(n1650), .Y(n2102) );
  NAND2X1 U1471 ( .A(\mem<13><3> ), .B(n88), .Y(n1651) );
  OAI21X1 U1472 ( .A(n1281), .B(n1319), .C(n1651), .Y(n2101) );
  NAND2X1 U1473 ( .A(\mem<13><4> ), .B(n88), .Y(n1652) );
  OAI21X1 U1474 ( .A(n1281), .B(n1321), .C(n1652), .Y(n2100) );
  NAND2X1 U1475 ( .A(\mem<13><5> ), .B(n88), .Y(n1653) );
  OAI21X1 U1476 ( .A(n1281), .B(n1323), .C(n1653), .Y(n2099) );
  NAND2X1 U1477 ( .A(\mem<13><6> ), .B(n88), .Y(n1654) );
  OAI21X1 U1478 ( .A(n1281), .B(n1325), .C(n1654), .Y(n2098) );
  NAND2X1 U1479 ( .A(\mem<13><7> ), .B(n88), .Y(n1655) );
  OAI21X1 U1480 ( .A(n1281), .B(n1327), .C(n1655), .Y(n2097) );
  NAND2X1 U1481 ( .A(\mem<13><8> ), .B(n88), .Y(n1656) );
  OAI21X1 U1482 ( .A(n1282), .B(n1329), .C(n1656), .Y(n2096) );
  NAND2X1 U1483 ( .A(\mem<13><9> ), .B(n88), .Y(n1657) );
  OAI21X1 U1484 ( .A(n1282), .B(n1331), .C(n1657), .Y(n2095) );
  NAND2X1 U1485 ( .A(\mem<13><10> ), .B(n88), .Y(n1658) );
  OAI21X1 U1486 ( .A(n1282), .B(n1333), .C(n1658), .Y(n2094) );
  NAND2X1 U1487 ( .A(\mem<13><11> ), .B(n88), .Y(n1659) );
  OAI21X1 U1488 ( .A(n1282), .B(n1335), .C(n1659), .Y(n2093) );
  NAND2X1 U1489 ( .A(\mem<13><12> ), .B(n88), .Y(n1660) );
  OAI21X1 U1490 ( .A(n1282), .B(n1337), .C(n1660), .Y(n2092) );
  NAND2X1 U1491 ( .A(\mem<13><13> ), .B(n88), .Y(n1661) );
  OAI21X1 U1492 ( .A(n1282), .B(n1339), .C(n1661), .Y(n2091) );
  NAND2X1 U1493 ( .A(\mem<13><14> ), .B(n88), .Y(n1662) );
  OAI21X1 U1494 ( .A(n1282), .B(n1341), .C(n1662), .Y(n2090) );
  NAND2X1 U1495 ( .A(\mem<13><15> ), .B(n88), .Y(n1663) );
  OAI21X1 U1496 ( .A(n1282), .B(n1343), .C(n1663), .Y(n2089) );
  NAND2X1 U1497 ( .A(\mem<12><0> ), .B(n90), .Y(n1664) );
  OAI21X1 U1498 ( .A(n1283), .B(n1313), .C(n1664), .Y(n2088) );
  NAND2X1 U1499 ( .A(\mem<12><1> ), .B(n90), .Y(n1665) );
  OAI21X1 U1500 ( .A(n1283), .B(n1315), .C(n1665), .Y(n2087) );
  NAND2X1 U1501 ( .A(\mem<12><2> ), .B(n90), .Y(n1666) );
  OAI21X1 U1502 ( .A(n1283), .B(n1317), .C(n1666), .Y(n2086) );
  NAND2X1 U1503 ( .A(\mem<12><3> ), .B(n90), .Y(n1667) );
  OAI21X1 U1504 ( .A(n1283), .B(n1319), .C(n1667), .Y(n2085) );
  NAND2X1 U1505 ( .A(\mem<12><4> ), .B(n90), .Y(n1668) );
  OAI21X1 U1506 ( .A(n1283), .B(n1321), .C(n1668), .Y(n2084) );
  NAND2X1 U1507 ( .A(\mem<12><5> ), .B(n90), .Y(n1669) );
  OAI21X1 U1508 ( .A(n1283), .B(n1323), .C(n1669), .Y(n2083) );
  NAND2X1 U1509 ( .A(\mem<12><6> ), .B(n90), .Y(n1670) );
  OAI21X1 U1510 ( .A(n1283), .B(n1325), .C(n1670), .Y(n2082) );
  NAND2X1 U1511 ( .A(\mem<12><7> ), .B(n90), .Y(n1671) );
  OAI21X1 U1512 ( .A(n1283), .B(n1326), .C(n1671), .Y(n2081) );
  NAND2X1 U1513 ( .A(\mem<12><8> ), .B(n90), .Y(n1672) );
  OAI21X1 U1514 ( .A(n1284), .B(n1329), .C(n1672), .Y(n2080) );
  NAND2X1 U1515 ( .A(\mem<12><9> ), .B(n90), .Y(n1673) );
  OAI21X1 U1516 ( .A(n1284), .B(n1331), .C(n1673), .Y(n2079) );
  NAND2X1 U1517 ( .A(\mem<12><10> ), .B(n90), .Y(n1674) );
  OAI21X1 U1518 ( .A(n1284), .B(n1333), .C(n1674), .Y(n2078) );
  NAND2X1 U1519 ( .A(\mem<12><11> ), .B(n90), .Y(n1675) );
  OAI21X1 U1520 ( .A(n1284), .B(n1335), .C(n1675), .Y(n2077) );
  NAND2X1 U1521 ( .A(\mem<12><12> ), .B(n90), .Y(n1676) );
  OAI21X1 U1522 ( .A(n1284), .B(n1337), .C(n1676), .Y(n2076) );
  NAND2X1 U1523 ( .A(\mem<12><13> ), .B(n90), .Y(n1677) );
  OAI21X1 U1524 ( .A(n1284), .B(n1339), .C(n1677), .Y(n2075) );
  NAND2X1 U1525 ( .A(\mem<12><14> ), .B(n90), .Y(n1678) );
  OAI21X1 U1526 ( .A(n1284), .B(n1341), .C(n1678), .Y(n2074) );
  NAND2X1 U1527 ( .A(\mem<12><15> ), .B(n90), .Y(n1679) );
  OAI21X1 U1528 ( .A(n1284), .B(n1343), .C(n1679), .Y(n2073) );
  NAND2X1 U1529 ( .A(\mem<11><0> ), .B(n92), .Y(n1680) );
  OAI21X1 U1530 ( .A(n1285), .B(n1313), .C(n1680), .Y(n2072) );
  NAND2X1 U1531 ( .A(\mem<11><1> ), .B(n92), .Y(n1681) );
  OAI21X1 U1532 ( .A(n1285), .B(n1314), .C(n1681), .Y(n2071) );
  NAND2X1 U1533 ( .A(\mem<11><2> ), .B(n92), .Y(n1682) );
  OAI21X1 U1534 ( .A(n1285), .B(n1316), .C(n1682), .Y(n2070) );
  NAND2X1 U1535 ( .A(\mem<11><3> ), .B(n92), .Y(n1683) );
  OAI21X1 U1536 ( .A(n1285), .B(n1318), .C(n1683), .Y(n2069) );
  NAND2X1 U1537 ( .A(\mem<11><4> ), .B(n92), .Y(n1684) );
  OAI21X1 U1538 ( .A(n1285), .B(n1320), .C(n1684), .Y(n2068) );
  NAND2X1 U1539 ( .A(\mem<11><5> ), .B(n92), .Y(n1685) );
  OAI21X1 U1540 ( .A(n1285), .B(n1322), .C(n1685), .Y(n2067) );
  NAND2X1 U1541 ( .A(\mem<11><6> ), .B(n92), .Y(n1686) );
  OAI21X1 U1542 ( .A(n1285), .B(n1324), .C(n1686), .Y(n2066) );
  NAND2X1 U1543 ( .A(\mem<11><7> ), .B(n92), .Y(n1687) );
  OAI21X1 U1544 ( .A(n1285), .B(n1326), .C(n1687), .Y(n2065) );
  NAND2X1 U1545 ( .A(\mem<11><8> ), .B(n92), .Y(n1688) );
  OAI21X1 U1546 ( .A(n1286), .B(n1328), .C(n1688), .Y(n2064) );
  NAND2X1 U1547 ( .A(\mem<11><9> ), .B(n92), .Y(n1689) );
  OAI21X1 U1548 ( .A(n1286), .B(n1330), .C(n1689), .Y(n2063) );
  NAND2X1 U1549 ( .A(\mem<11><10> ), .B(n92), .Y(n1690) );
  OAI21X1 U1550 ( .A(n1286), .B(n1332), .C(n1690), .Y(n2062) );
  NAND2X1 U1551 ( .A(\mem<11><11> ), .B(n92), .Y(n1691) );
  OAI21X1 U1552 ( .A(n1286), .B(n1334), .C(n1691), .Y(n2061) );
  NAND2X1 U1553 ( .A(\mem<11><12> ), .B(n92), .Y(n1692) );
  OAI21X1 U1554 ( .A(n1286), .B(n1336), .C(n1692), .Y(n2060) );
  NAND2X1 U1555 ( .A(\mem<11><13> ), .B(n92), .Y(n1693) );
  OAI21X1 U1556 ( .A(n1286), .B(n1338), .C(n1693), .Y(n2059) );
  NAND2X1 U1557 ( .A(\mem<11><14> ), .B(n92), .Y(n1694) );
  OAI21X1 U1558 ( .A(n1286), .B(n1340), .C(n1694), .Y(n2058) );
  NAND2X1 U1559 ( .A(\mem<11><15> ), .B(n92), .Y(n1695) );
  OAI21X1 U1560 ( .A(n1286), .B(n1342), .C(n1695), .Y(n2057) );
  NAND2X1 U1561 ( .A(\mem<10><0> ), .B(n1), .Y(n1696) );
  OAI21X1 U1562 ( .A(n1287), .B(n1313), .C(n1696), .Y(n2056) );
  NAND2X1 U1563 ( .A(\mem<10><1> ), .B(n1), .Y(n1697) );
  OAI21X1 U1564 ( .A(n1287), .B(n1314), .C(n1697), .Y(n2055) );
  NAND2X1 U1565 ( .A(\mem<10><2> ), .B(n1), .Y(n1698) );
  OAI21X1 U1566 ( .A(n1287), .B(n1316), .C(n1698), .Y(n2054) );
  NAND2X1 U1567 ( .A(\mem<10><3> ), .B(n1), .Y(n1699) );
  OAI21X1 U1568 ( .A(n1287), .B(n1318), .C(n1699), .Y(n2053) );
  NAND2X1 U1569 ( .A(\mem<10><4> ), .B(n1), .Y(n1700) );
  OAI21X1 U1570 ( .A(n1287), .B(n1320), .C(n1700), .Y(n2052) );
  NAND2X1 U1571 ( .A(\mem<10><5> ), .B(n1), .Y(n1701) );
  OAI21X1 U1572 ( .A(n1287), .B(n1322), .C(n1701), .Y(n2051) );
  NAND2X1 U1573 ( .A(\mem<10><6> ), .B(n1), .Y(n1702) );
  OAI21X1 U1574 ( .A(n1287), .B(n1324), .C(n1702), .Y(n2050) );
  NAND2X1 U1575 ( .A(\mem<10><7> ), .B(n1), .Y(n1703) );
  OAI21X1 U1576 ( .A(n1287), .B(n1326), .C(n1703), .Y(n2049) );
  NAND2X1 U1577 ( .A(\mem<10><8> ), .B(n1), .Y(n1704) );
  OAI21X1 U1578 ( .A(n1288), .B(n1328), .C(n1704), .Y(n2048) );
  NAND2X1 U1579 ( .A(\mem<10><9> ), .B(n1), .Y(n1705) );
  OAI21X1 U1580 ( .A(n1288), .B(n1330), .C(n1705), .Y(n2047) );
  NAND2X1 U1581 ( .A(\mem<10><10> ), .B(n1), .Y(n1706) );
  OAI21X1 U1582 ( .A(n1288), .B(n1332), .C(n1706), .Y(n2046) );
  NAND2X1 U1583 ( .A(\mem<10><11> ), .B(n1), .Y(n1707) );
  OAI21X1 U1584 ( .A(n1288), .B(n1334), .C(n1707), .Y(n2045) );
  NAND2X1 U1585 ( .A(\mem<10><12> ), .B(n1), .Y(n1708) );
  OAI21X1 U1586 ( .A(n1288), .B(n1336), .C(n1708), .Y(n2044) );
  NAND2X1 U1587 ( .A(\mem<10><13> ), .B(n1), .Y(n1709) );
  OAI21X1 U1588 ( .A(n1288), .B(n1338), .C(n1709), .Y(n2043) );
  NAND2X1 U1589 ( .A(\mem<10><14> ), .B(n1), .Y(n1710) );
  OAI21X1 U1590 ( .A(n1288), .B(n1340), .C(n1710), .Y(n2042) );
  NAND2X1 U1591 ( .A(\mem<10><15> ), .B(n1), .Y(n1711) );
  OAI21X1 U1592 ( .A(n1288), .B(n1342), .C(n1711), .Y(n2041) );
  NAND2X1 U1593 ( .A(\mem<9><0> ), .B(n41), .Y(n1712) );
  OAI21X1 U1594 ( .A(n1289), .B(n1313), .C(n1712), .Y(n2040) );
  NAND2X1 U1595 ( .A(\mem<9><1> ), .B(n41), .Y(n1713) );
  OAI21X1 U1596 ( .A(n1289), .B(n1314), .C(n1713), .Y(n2039) );
  NAND2X1 U1597 ( .A(\mem<9><2> ), .B(n41), .Y(n1714) );
  OAI21X1 U1598 ( .A(n1289), .B(n1316), .C(n1714), .Y(n2038) );
  NAND2X1 U1599 ( .A(\mem<9><3> ), .B(n41), .Y(n1715) );
  OAI21X1 U1600 ( .A(n1289), .B(n1318), .C(n1715), .Y(n2037) );
  NAND2X1 U1601 ( .A(\mem<9><4> ), .B(n41), .Y(n1716) );
  OAI21X1 U1602 ( .A(n1289), .B(n1320), .C(n1716), .Y(n2036) );
  NAND2X1 U1603 ( .A(\mem<9><5> ), .B(n41), .Y(n1717) );
  OAI21X1 U1604 ( .A(n1289), .B(n1322), .C(n1717), .Y(n2035) );
  NAND2X1 U1605 ( .A(\mem<9><6> ), .B(n41), .Y(n1718) );
  OAI21X1 U1606 ( .A(n1289), .B(n1324), .C(n1718), .Y(n2034) );
  NAND2X1 U1607 ( .A(\mem<9><7> ), .B(n41), .Y(n1719) );
  OAI21X1 U1608 ( .A(n1289), .B(n1326), .C(n1719), .Y(n2033) );
  NAND2X1 U1609 ( .A(\mem<9><8> ), .B(n41), .Y(n1720) );
  OAI21X1 U1610 ( .A(n1290), .B(n1328), .C(n1720), .Y(n2032) );
  NAND2X1 U1611 ( .A(\mem<9><9> ), .B(n41), .Y(n1721) );
  OAI21X1 U1612 ( .A(n1290), .B(n1330), .C(n1721), .Y(n2031) );
  NAND2X1 U1613 ( .A(\mem<9><10> ), .B(n41), .Y(n1722) );
  OAI21X1 U1614 ( .A(n1290), .B(n1332), .C(n1722), .Y(n2030) );
  NAND2X1 U1615 ( .A(\mem<9><11> ), .B(n41), .Y(n1723) );
  OAI21X1 U1616 ( .A(n1290), .B(n1334), .C(n1723), .Y(n2029) );
  NAND2X1 U1617 ( .A(\mem<9><12> ), .B(n41), .Y(n1724) );
  OAI21X1 U1618 ( .A(n1290), .B(n1336), .C(n1724), .Y(n2028) );
  NAND2X1 U1619 ( .A(\mem<9><13> ), .B(n41), .Y(n1725) );
  OAI21X1 U1620 ( .A(n1290), .B(n1338), .C(n1725), .Y(n2027) );
  NAND2X1 U1621 ( .A(\mem<9><14> ), .B(n41), .Y(n1726) );
  OAI21X1 U1622 ( .A(n1290), .B(n1340), .C(n1726), .Y(n2026) );
  NAND2X1 U1623 ( .A(\mem<9><15> ), .B(n41), .Y(n1727) );
  OAI21X1 U1624 ( .A(n1290), .B(n1342), .C(n1727), .Y(n2025) );
  NAND2X1 U1625 ( .A(\mem<8><0> ), .B(n99), .Y(n1729) );
  OAI21X1 U1626 ( .A(n1291), .B(n1313), .C(n1729), .Y(n2024) );
  NAND2X1 U1627 ( .A(\mem<8><1> ), .B(n99), .Y(n1730) );
  OAI21X1 U1628 ( .A(n1291), .B(n1314), .C(n1730), .Y(n2023) );
  NAND2X1 U1629 ( .A(\mem<8><2> ), .B(n99), .Y(n1731) );
  OAI21X1 U1630 ( .A(n1291), .B(n1316), .C(n1731), .Y(n2022) );
  NAND2X1 U1631 ( .A(\mem<8><3> ), .B(n99), .Y(n1732) );
  OAI21X1 U1632 ( .A(n1291), .B(n1318), .C(n1732), .Y(n2021) );
  NAND2X1 U1633 ( .A(\mem<8><4> ), .B(n99), .Y(n1733) );
  OAI21X1 U1634 ( .A(n1291), .B(n1320), .C(n1733), .Y(n2020) );
  NAND2X1 U1635 ( .A(\mem<8><5> ), .B(n99), .Y(n1734) );
  OAI21X1 U1636 ( .A(n1291), .B(n1322), .C(n1734), .Y(n2019) );
  NAND2X1 U1637 ( .A(\mem<8><6> ), .B(n99), .Y(n1735) );
  OAI21X1 U1638 ( .A(n1291), .B(n1324), .C(n1735), .Y(n2018) );
  NAND2X1 U1639 ( .A(\mem<8><7> ), .B(n99), .Y(n1736) );
  OAI21X1 U1640 ( .A(n1291), .B(n1326), .C(n1736), .Y(n2017) );
  NAND2X1 U1641 ( .A(\mem<8><8> ), .B(n99), .Y(n1737) );
  OAI21X1 U1642 ( .A(n1291), .B(n1328), .C(n1737), .Y(n2016) );
  NAND2X1 U1643 ( .A(\mem<8><9> ), .B(n99), .Y(n1738) );
  OAI21X1 U1644 ( .A(n1291), .B(n1330), .C(n1738), .Y(n2015) );
  NAND2X1 U1645 ( .A(\mem<8><10> ), .B(n99), .Y(n1739) );
  OAI21X1 U1646 ( .A(n1291), .B(n1332), .C(n1739), .Y(n2014) );
  NAND2X1 U1647 ( .A(\mem<8><11> ), .B(n99), .Y(n1740) );
  OAI21X1 U1648 ( .A(n1291), .B(n1334), .C(n1740), .Y(n2013) );
  NAND2X1 U1649 ( .A(\mem<8><12> ), .B(n99), .Y(n1741) );
  OAI21X1 U1650 ( .A(n1291), .B(n1336), .C(n1741), .Y(n2012) );
  NAND2X1 U1651 ( .A(\mem<8><13> ), .B(n99), .Y(n1742) );
  OAI21X1 U1652 ( .A(n1291), .B(n1338), .C(n1742), .Y(n2011) );
  NAND2X1 U1653 ( .A(\mem<8><14> ), .B(n99), .Y(n1743) );
  OAI21X1 U1654 ( .A(n1291), .B(n1340), .C(n1743), .Y(n2010) );
  NAND2X1 U1655 ( .A(\mem<8><15> ), .B(n99), .Y(n1744) );
  OAI21X1 U1656 ( .A(n1291), .B(n1342), .C(n1744), .Y(n2009) );
  NAND3X1 U1657 ( .A(n1352), .B(n2393), .C(n1353), .Y(n1745) );
  NAND2X1 U1658 ( .A(\mem<7><0> ), .B(n100), .Y(n1746) );
  OAI21X1 U1659 ( .A(n1292), .B(n1312), .C(n1746), .Y(n2008) );
  NAND2X1 U1660 ( .A(\mem<7><1> ), .B(n100), .Y(n1747) );
  OAI21X1 U1661 ( .A(n1292), .B(n1314), .C(n1747), .Y(n2007) );
  NAND2X1 U1662 ( .A(\mem<7><2> ), .B(n100), .Y(n1748) );
  OAI21X1 U1663 ( .A(n1292), .B(n1316), .C(n1748), .Y(n2006) );
  NAND2X1 U1664 ( .A(\mem<7><3> ), .B(n100), .Y(n1749) );
  OAI21X1 U1665 ( .A(n1292), .B(n1318), .C(n1749), .Y(n2005) );
  NAND2X1 U1666 ( .A(\mem<7><4> ), .B(n100), .Y(n1750) );
  OAI21X1 U1667 ( .A(n1292), .B(n1320), .C(n1750), .Y(n2004) );
  NAND2X1 U1668 ( .A(\mem<7><5> ), .B(n100), .Y(n1751) );
  OAI21X1 U1669 ( .A(n1292), .B(n1322), .C(n1751), .Y(n2003) );
  NAND2X1 U1670 ( .A(\mem<7><6> ), .B(n100), .Y(n1752) );
  OAI21X1 U1671 ( .A(n1292), .B(n1324), .C(n1752), .Y(n2002) );
  NAND2X1 U1672 ( .A(\mem<7><7> ), .B(n100), .Y(n1753) );
  OAI21X1 U1673 ( .A(n1292), .B(n1326), .C(n1753), .Y(n2001) );
  NAND2X1 U1674 ( .A(\mem<7><8> ), .B(n100), .Y(n1754) );
  OAI21X1 U1675 ( .A(n1293), .B(n1328), .C(n1754), .Y(n2000) );
  NAND2X1 U1676 ( .A(\mem<7><9> ), .B(n100), .Y(n1755) );
  OAI21X1 U1677 ( .A(n1293), .B(n1330), .C(n1755), .Y(n1999) );
  NAND2X1 U1678 ( .A(\mem<7><10> ), .B(n100), .Y(n1756) );
  OAI21X1 U1679 ( .A(n1293), .B(n1332), .C(n1756), .Y(n1998) );
  NAND2X1 U1680 ( .A(\mem<7><11> ), .B(n100), .Y(n1757) );
  OAI21X1 U1681 ( .A(n1293), .B(n1334), .C(n1757), .Y(n1997) );
  NAND2X1 U1682 ( .A(\mem<7><12> ), .B(n100), .Y(n1758) );
  OAI21X1 U1683 ( .A(n1293), .B(n1336), .C(n1758), .Y(n1996) );
  NAND2X1 U1684 ( .A(\mem<7><13> ), .B(n100), .Y(n1759) );
  OAI21X1 U1685 ( .A(n1293), .B(n1338), .C(n1759), .Y(n1995) );
  NAND2X1 U1686 ( .A(\mem<7><14> ), .B(n100), .Y(n1760) );
  OAI21X1 U1687 ( .A(n1293), .B(n1340), .C(n1760), .Y(n1994) );
  NAND2X1 U1688 ( .A(\mem<7><15> ), .B(n100), .Y(n1761) );
  OAI21X1 U1689 ( .A(n1293), .B(n1342), .C(n1761), .Y(n1993) );
  NAND2X1 U1690 ( .A(\mem<6><0> ), .B(n101), .Y(n1762) );
  OAI21X1 U1691 ( .A(n1294), .B(n1313), .C(n1762), .Y(n1992) );
  NAND2X1 U1692 ( .A(\mem<6><1> ), .B(n101), .Y(n1763) );
  OAI21X1 U1693 ( .A(n1294), .B(n1314), .C(n1763), .Y(n1991) );
  NAND2X1 U1694 ( .A(\mem<6><2> ), .B(n101), .Y(n1764) );
  OAI21X1 U1695 ( .A(n1294), .B(n1316), .C(n1764), .Y(n1990) );
  NAND2X1 U1696 ( .A(\mem<6><3> ), .B(n101), .Y(n1765) );
  OAI21X1 U1697 ( .A(n1294), .B(n1318), .C(n1765), .Y(n1989) );
  NAND2X1 U1698 ( .A(\mem<6><4> ), .B(n101), .Y(n1766) );
  OAI21X1 U1699 ( .A(n1294), .B(n1320), .C(n1766), .Y(n1988) );
  NAND2X1 U1700 ( .A(\mem<6><5> ), .B(n101), .Y(n1767) );
  OAI21X1 U1701 ( .A(n1294), .B(n1322), .C(n1767), .Y(n1987) );
  NAND2X1 U1702 ( .A(\mem<6><6> ), .B(n101), .Y(n1768) );
  OAI21X1 U1703 ( .A(n1294), .B(n1324), .C(n1768), .Y(n1986) );
  NAND2X1 U1704 ( .A(\mem<6><7> ), .B(n101), .Y(n1769) );
  OAI21X1 U1705 ( .A(n1294), .B(n1326), .C(n1769), .Y(n1985) );
  NAND2X1 U1706 ( .A(\mem<6><8> ), .B(n101), .Y(n1770) );
  OAI21X1 U1707 ( .A(n1295), .B(n1328), .C(n1770), .Y(n1984) );
  NAND2X1 U1708 ( .A(\mem<6><9> ), .B(n101), .Y(n1771) );
  OAI21X1 U1709 ( .A(n1295), .B(n1330), .C(n1771), .Y(n1983) );
  NAND2X1 U1710 ( .A(\mem<6><10> ), .B(n101), .Y(n1772) );
  OAI21X1 U1711 ( .A(n1295), .B(n1332), .C(n1772), .Y(n1982) );
  NAND2X1 U1712 ( .A(\mem<6><11> ), .B(n101), .Y(n1773) );
  OAI21X1 U1713 ( .A(n1295), .B(n1334), .C(n1773), .Y(n1981) );
  NAND2X1 U1714 ( .A(\mem<6><12> ), .B(n101), .Y(n1774) );
  OAI21X1 U1715 ( .A(n1295), .B(n1336), .C(n1774), .Y(n1980) );
  NAND2X1 U1716 ( .A(\mem<6><13> ), .B(n101), .Y(n1775) );
  OAI21X1 U1717 ( .A(n1295), .B(n1338), .C(n1775), .Y(n1979) );
  NAND2X1 U1718 ( .A(\mem<6><14> ), .B(n101), .Y(n1776) );
  OAI21X1 U1719 ( .A(n1295), .B(n1340), .C(n1776), .Y(n1978) );
  NAND2X1 U1720 ( .A(\mem<6><15> ), .B(n101), .Y(n1777) );
  OAI21X1 U1721 ( .A(n1295), .B(n1342), .C(n1777), .Y(n1977) );
  NAND2X1 U1722 ( .A(\mem<5><0> ), .B(n102), .Y(n1779) );
  OAI21X1 U1723 ( .A(n1296), .B(n1312), .C(n1779), .Y(n1976) );
  NAND2X1 U1724 ( .A(\mem<5><1> ), .B(n102), .Y(n1780) );
  OAI21X1 U1725 ( .A(n1296), .B(n1314), .C(n1780), .Y(n1975) );
  NAND2X1 U1726 ( .A(\mem<5><2> ), .B(n102), .Y(n1781) );
  OAI21X1 U1727 ( .A(n1296), .B(n1316), .C(n1781), .Y(n1974) );
  NAND2X1 U1728 ( .A(\mem<5><3> ), .B(n102), .Y(n1782) );
  OAI21X1 U1729 ( .A(n1296), .B(n1318), .C(n1782), .Y(n1973) );
  NAND2X1 U1730 ( .A(\mem<5><4> ), .B(n102), .Y(n1783) );
  OAI21X1 U1731 ( .A(n1296), .B(n1320), .C(n1783), .Y(n1972) );
  NAND2X1 U1732 ( .A(\mem<5><5> ), .B(n102), .Y(n1784) );
  OAI21X1 U1733 ( .A(n1296), .B(n1322), .C(n1784), .Y(n1971) );
  NAND2X1 U1734 ( .A(\mem<5><6> ), .B(n102), .Y(n1785) );
  OAI21X1 U1735 ( .A(n1296), .B(n1324), .C(n1785), .Y(n1970) );
  NAND2X1 U1736 ( .A(\mem<5><7> ), .B(n102), .Y(n1786) );
  OAI21X1 U1737 ( .A(n1296), .B(n1326), .C(n1786), .Y(n1969) );
  NAND2X1 U1738 ( .A(\mem<5><8> ), .B(n102), .Y(n1787) );
  OAI21X1 U1739 ( .A(n1297), .B(n1328), .C(n1787), .Y(n1968) );
  NAND2X1 U1740 ( .A(\mem<5><9> ), .B(n102), .Y(n1788) );
  OAI21X1 U1741 ( .A(n1297), .B(n1330), .C(n1788), .Y(n1967) );
  NAND2X1 U1742 ( .A(\mem<5><10> ), .B(n102), .Y(n1789) );
  OAI21X1 U1743 ( .A(n1297), .B(n1332), .C(n1789), .Y(n1966) );
  NAND2X1 U1744 ( .A(\mem<5><11> ), .B(n102), .Y(n1790) );
  OAI21X1 U1745 ( .A(n1297), .B(n1334), .C(n1790), .Y(n1965) );
  NAND2X1 U1746 ( .A(\mem<5><12> ), .B(n102), .Y(n1791) );
  OAI21X1 U1747 ( .A(n1297), .B(n1336), .C(n1791), .Y(n1964) );
  NAND2X1 U1748 ( .A(\mem<5><13> ), .B(n102), .Y(n1792) );
  OAI21X1 U1749 ( .A(n1297), .B(n1338), .C(n1792), .Y(n1963) );
  NAND2X1 U1750 ( .A(\mem<5><14> ), .B(n102), .Y(n1793) );
  OAI21X1 U1751 ( .A(n1297), .B(n1340), .C(n1793), .Y(n1962) );
  NAND2X1 U1752 ( .A(\mem<5><15> ), .B(n102), .Y(n1794) );
  OAI21X1 U1753 ( .A(n1297), .B(n1342), .C(n1794), .Y(n1961) );
  NAND2X1 U1754 ( .A(\mem<4><0> ), .B(n103), .Y(n1796) );
  OAI21X1 U1755 ( .A(n1298), .B(n1313), .C(n1796), .Y(n1960) );
  NAND2X1 U1756 ( .A(\mem<4><1> ), .B(n103), .Y(n1797) );
  OAI21X1 U1757 ( .A(n1298), .B(n1314), .C(n1797), .Y(n1959) );
  NAND2X1 U1758 ( .A(\mem<4><2> ), .B(n103), .Y(n1798) );
  OAI21X1 U1759 ( .A(n1298), .B(n1316), .C(n1798), .Y(n1958) );
  NAND2X1 U1760 ( .A(\mem<4><3> ), .B(n103), .Y(n1799) );
  OAI21X1 U1761 ( .A(n1298), .B(n1318), .C(n1799), .Y(n1957) );
  NAND2X1 U1762 ( .A(\mem<4><4> ), .B(n103), .Y(n1800) );
  OAI21X1 U1763 ( .A(n1298), .B(n1320), .C(n1800), .Y(n1956) );
  NAND2X1 U1764 ( .A(\mem<4><5> ), .B(n103), .Y(n1801) );
  OAI21X1 U1765 ( .A(n1298), .B(n1322), .C(n1801), .Y(n1955) );
  NAND2X1 U1766 ( .A(\mem<4><6> ), .B(n103), .Y(n1802) );
  OAI21X1 U1767 ( .A(n1298), .B(n1324), .C(n1802), .Y(n1954) );
  NAND2X1 U1768 ( .A(\mem<4><7> ), .B(n103), .Y(n1803) );
  OAI21X1 U1769 ( .A(n1298), .B(n1326), .C(n1803), .Y(n1953) );
  NAND2X1 U1770 ( .A(\mem<4><8> ), .B(n103), .Y(n1804) );
  OAI21X1 U1771 ( .A(n1299), .B(n1328), .C(n1804), .Y(n1952) );
  NAND2X1 U1772 ( .A(\mem<4><9> ), .B(n103), .Y(n1805) );
  OAI21X1 U1773 ( .A(n1299), .B(n1330), .C(n1805), .Y(n1951) );
  NAND2X1 U1774 ( .A(\mem<4><10> ), .B(n103), .Y(n1806) );
  OAI21X1 U1775 ( .A(n1299), .B(n1332), .C(n1806), .Y(n1950) );
  NAND2X1 U1776 ( .A(\mem<4><11> ), .B(n103), .Y(n1807) );
  OAI21X1 U1777 ( .A(n1299), .B(n1334), .C(n1807), .Y(n1949) );
  NAND2X1 U1778 ( .A(\mem<4><12> ), .B(n103), .Y(n1808) );
  OAI21X1 U1779 ( .A(n1299), .B(n1336), .C(n1808), .Y(n1948) );
  NAND2X1 U1780 ( .A(\mem<4><13> ), .B(n103), .Y(n1809) );
  OAI21X1 U1781 ( .A(n1299), .B(n1338), .C(n1809), .Y(n1947) );
  NAND2X1 U1782 ( .A(\mem<4><14> ), .B(n103), .Y(n1810) );
  OAI21X1 U1783 ( .A(n1299), .B(n1340), .C(n1810), .Y(n1946) );
  NAND2X1 U1784 ( .A(\mem<4><15> ), .B(n103), .Y(n1811) );
  OAI21X1 U1785 ( .A(n1299), .B(n1342), .C(n1811), .Y(n1945) );
  NAND2X1 U1786 ( .A(\mem<3><0> ), .B(n104), .Y(n1813) );
  OAI21X1 U1787 ( .A(n1300), .B(n1312), .C(n1813), .Y(n1944) );
  NAND2X1 U1788 ( .A(\mem<3><1> ), .B(n104), .Y(n1814) );
  OAI21X1 U1789 ( .A(n1300), .B(n1314), .C(n1814), .Y(n1943) );
  NAND2X1 U1790 ( .A(\mem<3><2> ), .B(n104), .Y(n1815) );
  OAI21X1 U1791 ( .A(n1300), .B(n1316), .C(n1815), .Y(n1942) );
  NAND2X1 U1792 ( .A(\mem<3><3> ), .B(n104), .Y(n1816) );
  OAI21X1 U1793 ( .A(n1300), .B(n1318), .C(n1816), .Y(n1941) );
  NAND2X1 U1794 ( .A(\mem<3><4> ), .B(n104), .Y(n1817) );
  OAI21X1 U1795 ( .A(n1300), .B(n1320), .C(n1817), .Y(n1940) );
  NAND2X1 U1796 ( .A(\mem<3><5> ), .B(n104), .Y(n1818) );
  OAI21X1 U1797 ( .A(n1300), .B(n1322), .C(n1818), .Y(n1939) );
  NAND2X1 U1798 ( .A(\mem<3><6> ), .B(n104), .Y(n1819) );
  OAI21X1 U1799 ( .A(n1300), .B(n1324), .C(n1819), .Y(n1938) );
  NAND2X1 U1800 ( .A(\mem<3><7> ), .B(n104), .Y(n1820) );
  OAI21X1 U1801 ( .A(n1300), .B(n1326), .C(n1820), .Y(n1937) );
  NAND2X1 U1802 ( .A(\mem<3><8> ), .B(n104), .Y(n1821) );
  OAI21X1 U1803 ( .A(n1301), .B(n1328), .C(n1821), .Y(n1936) );
  NAND2X1 U1804 ( .A(\mem<3><9> ), .B(n104), .Y(n1822) );
  OAI21X1 U1805 ( .A(n1301), .B(n1330), .C(n1822), .Y(n1935) );
  NAND2X1 U1806 ( .A(\mem<3><10> ), .B(n104), .Y(n1823) );
  OAI21X1 U1807 ( .A(n1301), .B(n1332), .C(n1823), .Y(n1934) );
  NAND2X1 U1808 ( .A(\mem<3><11> ), .B(n104), .Y(n1824) );
  OAI21X1 U1809 ( .A(n1301), .B(n1334), .C(n1824), .Y(n1933) );
  NAND2X1 U1810 ( .A(\mem<3><12> ), .B(n104), .Y(n1825) );
  OAI21X1 U1811 ( .A(n1301), .B(n1336), .C(n1825), .Y(n1932) );
  NAND2X1 U1812 ( .A(\mem<3><13> ), .B(n104), .Y(n1826) );
  OAI21X1 U1813 ( .A(n1301), .B(n1338), .C(n1826), .Y(n1931) );
  NAND2X1 U1814 ( .A(\mem<3><14> ), .B(n104), .Y(n1827) );
  OAI21X1 U1815 ( .A(n1301), .B(n1340), .C(n1827), .Y(n1930) );
  NAND2X1 U1816 ( .A(\mem<3><15> ), .B(n104), .Y(n1828) );
  OAI21X1 U1817 ( .A(n1301), .B(n1342), .C(n1828), .Y(n1929) );
  NAND2X1 U1818 ( .A(\mem<2><0> ), .B(n105), .Y(n1830) );
  OAI21X1 U1819 ( .A(n1302), .B(n1313), .C(n1830), .Y(n1928) );
  NAND2X1 U1820 ( .A(\mem<2><1> ), .B(n105), .Y(n1831) );
  OAI21X1 U1821 ( .A(n1302), .B(n1314), .C(n1831), .Y(n1927) );
  NAND2X1 U1822 ( .A(\mem<2><2> ), .B(n105), .Y(n1832) );
  OAI21X1 U1823 ( .A(n1302), .B(n1316), .C(n1832), .Y(n1926) );
  NAND2X1 U1824 ( .A(\mem<2><3> ), .B(n105), .Y(n1833) );
  OAI21X1 U1825 ( .A(n1302), .B(n1318), .C(n1833), .Y(n1925) );
  NAND2X1 U1826 ( .A(\mem<2><4> ), .B(n105), .Y(n1834) );
  OAI21X1 U1827 ( .A(n1302), .B(n1320), .C(n1834), .Y(n1924) );
  NAND2X1 U1828 ( .A(\mem<2><5> ), .B(n105), .Y(n1835) );
  OAI21X1 U1829 ( .A(n1302), .B(n1322), .C(n1835), .Y(n1923) );
  NAND2X1 U1830 ( .A(\mem<2><6> ), .B(n105), .Y(n1836) );
  OAI21X1 U1831 ( .A(n1302), .B(n1324), .C(n1836), .Y(n1922) );
  NAND2X1 U1832 ( .A(\mem<2><7> ), .B(n105), .Y(n1837) );
  OAI21X1 U1833 ( .A(n1302), .B(n1326), .C(n1837), .Y(n1921) );
  NAND2X1 U1834 ( .A(\mem<2><8> ), .B(n105), .Y(n1838) );
  OAI21X1 U1835 ( .A(n1303), .B(n1328), .C(n1838), .Y(n1920) );
  NAND2X1 U1836 ( .A(\mem<2><9> ), .B(n105), .Y(n1839) );
  OAI21X1 U1837 ( .A(n1303), .B(n1330), .C(n1839), .Y(n1919) );
  NAND2X1 U1838 ( .A(\mem<2><10> ), .B(n105), .Y(n1840) );
  OAI21X1 U1839 ( .A(n1303), .B(n1332), .C(n1840), .Y(n1918) );
  NAND2X1 U1840 ( .A(\mem<2><11> ), .B(n105), .Y(n1841) );
  OAI21X1 U1841 ( .A(n1303), .B(n1334), .C(n1841), .Y(n1917) );
  NAND2X1 U1842 ( .A(\mem<2><12> ), .B(n105), .Y(n1842) );
  OAI21X1 U1843 ( .A(n1303), .B(n1336), .C(n1842), .Y(n1916) );
  NAND2X1 U1844 ( .A(\mem<2><13> ), .B(n105), .Y(n1843) );
  OAI21X1 U1845 ( .A(n1303), .B(n1338), .C(n1843), .Y(n1915) );
  NAND2X1 U1846 ( .A(\mem<2><14> ), .B(n105), .Y(n1844) );
  OAI21X1 U1847 ( .A(n1303), .B(n1340), .C(n1844), .Y(n1914) );
  NAND2X1 U1848 ( .A(\mem<2><15> ), .B(n105), .Y(n1845) );
  OAI21X1 U1849 ( .A(n1303), .B(n1342), .C(n1845), .Y(n1913) );
  NAND2X1 U1850 ( .A(\mem<1><0> ), .B(n106), .Y(n1847) );
  OAI21X1 U1851 ( .A(n1304), .B(n1312), .C(n1847), .Y(n1912) );
  NAND2X1 U1852 ( .A(\mem<1><1> ), .B(n106), .Y(n1848) );
  OAI21X1 U1853 ( .A(n1304), .B(n1314), .C(n1848), .Y(n1911) );
  NAND2X1 U1854 ( .A(\mem<1><2> ), .B(n106), .Y(n1849) );
  OAI21X1 U1855 ( .A(n1304), .B(n1316), .C(n1849), .Y(n1910) );
  NAND2X1 U1856 ( .A(\mem<1><3> ), .B(n106), .Y(n1850) );
  OAI21X1 U1857 ( .A(n1304), .B(n1318), .C(n1850), .Y(n1909) );
  NAND2X1 U1858 ( .A(\mem<1><4> ), .B(n106), .Y(n1851) );
  OAI21X1 U1859 ( .A(n1304), .B(n1320), .C(n1851), .Y(n1908) );
  NAND2X1 U1860 ( .A(\mem<1><5> ), .B(n106), .Y(n1852) );
  OAI21X1 U1861 ( .A(n1304), .B(n1322), .C(n1852), .Y(n1907) );
  NAND2X1 U1862 ( .A(\mem<1><6> ), .B(n106), .Y(n1853) );
  OAI21X1 U1863 ( .A(n1304), .B(n1324), .C(n1853), .Y(n1906) );
  NAND2X1 U1864 ( .A(\mem<1><7> ), .B(n106), .Y(n1854) );
  OAI21X1 U1865 ( .A(n1304), .B(n1326), .C(n1854), .Y(n1905) );
  NAND2X1 U1866 ( .A(\mem<1><8> ), .B(n106), .Y(n1855) );
  OAI21X1 U1867 ( .A(n1305), .B(n1328), .C(n1855), .Y(n1904) );
  NAND2X1 U1868 ( .A(\mem<1><9> ), .B(n106), .Y(n1856) );
  OAI21X1 U1869 ( .A(n1305), .B(n1330), .C(n1856), .Y(n1903) );
  NAND2X1 U1870 ( .A(\mem<1><10> ), .B(n106), .Y(n1857) );
  OAI21X1 U1871 ( .A(n1305), .B(n1332), .C(n1857), .Y(n1902) );
  NAND2X1 U1872 ( .A(\mem<1><11> ), .B(n106), .Y(n1858) );
  OAI21X1 U1873 ( .A(n1305), .B(n1334), .C(n1858), .Y(n1901) );
  NAND2X1 U1874 ( .A(\mem<1><12> ), .B(n106), .Y(n1859) );
  OAI21X1 U1875 ( .A(n1305), .B(n1336), .C(n1859), .Y(n1900) );
  NAND2X1 U1876 ( .A(\mem<1><13> ), .B(n106), .Y(n1860) );
  OAI21X1 U1877 ( .A(n1305), .B(n1338), .C(n1860), .Y(n1899) );
  NAND2X1 U1878 ( .A(\mem<1><14> ), .B(n106), .Y(n1861) );
  OAI21X1 U1879 ( .A(n1305), .B(n1340), .C(n1861), .Y(n1898) );
  NAND2X1 U1880 ( .A(\mem<1><15> ), .B(n106), .Y(n1862) );
  OAI21X1 U1881 ( .A(n1305), .B(n1342), .C(n1862), .Y(n1897) );
  NAND2X1 U1882 ( .A(\mem<0><0> ), .B(n43), .Y(n1865) );
  OAI21X1 U1883 ( .A(n1306), .B(n1313), .C(n1865), .Y(n1896) );
  NAND2X1 U1884 ( .A(\mem<0><1> ), .B(n43), .Y(n1866) );
  OAI21X1 U1885 ( .A(n1306), .B(n1314), .C(n1866), .Y(n1895) );
  NAND2X1 U1886 ( .A(\mem<0><2> ), .B(n43), .Y(n1867) );
  OAI21X1 U1887 ( .A(n1306), .B(n1316), .C(n1867), .Y(n1894) );
  NAND2X1 U1888 ( .A(\mem<0><3> ), .B(n43), .Y(n1868) );
  OAI21X1 U1889 ( .A(n1306), .B(n1318), .C(n1868), .Y(n1893) );
  NAND2X1 U1890 ( .A(\mem<0><4> ), .B(n43), .Y(n1869) );
  OAI21X1 U1891 ( .A(n1306), .B(n1320), .C(n1869), .Y(n1892) );
  NAND2X1 U1892 ( .A(\mem<0><5> ), .B(n43), .Y(n1870) );
  OAI21X1 U1893 ( .A(n1306), .B(n1322), .C(n1870), .Y(n1891) );
  NAND2X1 U1894 ( .A(\mem<0><6> ), .B(n43), .Y(n1871) );
  OAI21X1 U1895 ( .A(n1306), .B(n1324), .C(n1871), .Y(n1890) );
  NAND2X1 U1896 ( .A(\mem<0><7> ), .B(n43), .Y(n1872) );
  OAI21X1 U1897 ( .A(n1306), .B(n1326), .C(n1872), .Y(n1889) );
  NAND2X1 U1898 ( .A(\mem<0><8> ), .B(n43), .Y(n1873) );
  OAI21X1 U1899 ( .A(n1306), .B(n1328), .C(n1873), .Y(n1888) );
  NAND2X1 U1900 ( .A(\mem<0><9> ), .B(n43), .Y(n1874) );
  OAI21X1 U1901 ( .A(n1306), .B(n1330), .C(n1874), .Y(n1887) );
  NAND2X1 U1902 ( .A(\mem<0><10> ), .B(n43), .Y(n1875) );
  OAI21X1 U1903 ( .A(n1306), .B(n1332), .C(n1875), .Y(n1886) );
  NAND2X1 U1904 ( .A(\mem<0><11> ), .B(n43), .Y(n1876) );
  OAI21X1 U1905 ( .A(n1306), .B(n1334), .C(n1876), .Y(n1885) );
  NAND2X1 U1906 ( .A(\mem<0><12> ), .B(n43), .Y(n1877) );
  OAI21X1 U1907 ( .A(n1306), .B(n1336), .C(n1877), .Y(n1884) );
  NAND2X1 U1908 ( .A(\mem<0><13> ), .B(n43), .Y(n1878) );
  OAI21X1 U1909 ( .A(n1306), .B(n1338), .C(n1878), .Y(n1883) );
  NAND2X1 U1910 ( .A(\mem<0><14> ), .B(n43), .Y(n1879) );
  OAI21X1 U1911 ( .A(n1306), .B(n1340), .C(n1879), .Y(n1882) );
  NAND2X1 U1912 ( .A(\mem<0><15> ), .B(n43), .Y(n1880) );
  OAI21X1 U1913 ( .A(n1306), .B(n1342), .C(n1880), .Y(n1881) );
endmodule


module memc_Size16_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1895), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1896), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1897), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1898), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1899), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1900), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1901), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1902), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1903), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1904), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1905), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1906), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1907), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1908), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1909), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1910), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1911), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1912), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1913), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1914), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1915), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1916), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1917), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1918), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1919), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1920), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1921), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1922), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1923), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1924), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1925), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1926), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1927), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1928), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1929), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1930), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1931), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1932), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1933), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1934), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1935), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1936), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1937), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1938), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1939), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1940), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1941), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1942), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1943), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1944), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1945), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1946), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1947), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1948), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1949), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1950), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1951), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1952), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1953), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1954), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1955), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1956), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1957), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1958), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1959), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1960), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1961), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1962), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1963), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1964), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1965), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1966), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1967), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1968), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1969), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1970), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1971), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1972), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1973), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1974), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1975), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1976), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1977), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1978), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1979), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1980), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1981), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1982), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1983), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1984), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1985), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1986), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1987), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1988), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1989), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1990), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1991), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1992), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1993), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1994), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1995), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1996), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1997), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1998), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1999), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2000), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2001), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2002), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2003), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2004), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2005), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2006), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2007), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2008), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2009), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2010), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2011), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2012), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2013), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2014), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2015), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2016), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2017), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2018), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2019), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2020), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2021), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2022), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2023), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2024), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2025), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2026), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2027), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2028), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2029), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2030), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2031), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2032), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2033), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2034), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2035), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2036), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2037), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2038), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2039), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2040), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2041), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2042), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2043), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2044), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2045), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2046), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2047), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2048), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2049), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2050), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2051), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2052), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2053), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2054), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2055), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2056), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2057), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2058), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2059), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2060), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2061), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2062), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2063), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2064), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2065), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2066), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2067), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2068), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2069), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2070), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2071), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2072), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2073), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2074), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2075), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2076), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2077), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2078), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2079), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2080), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2081), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2082), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2083), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2084), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2085), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2086), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2087), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2088), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2089), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2090), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2091), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2092), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2093), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2094), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2095), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2096), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2097), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2098), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2099), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2100), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2101), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2102), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2103), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2104), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2105), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2106), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2107), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2108), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2109), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2110), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2111), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2112), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2113), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2114), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2115), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2116), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2117), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2118), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2119), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2120), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2121), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2122), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2123), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2124), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2125), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2126), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2127), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2128), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2129), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2130), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2131), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2132), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2133), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2134), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2135), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2136), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2137), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2138), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2139), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2140), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2141), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2142), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2143), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2144), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2145), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2146), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2147), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2148), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2149), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2150), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2151), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2152), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2153), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2154), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2155), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2156), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2157), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2158), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2159), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2160), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2161), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2162), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2163), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2164), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2165), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2166), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2167), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2168), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2169), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2170), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2171), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2172), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2173), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2174), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2175), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2176), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2177), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2178), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2179), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2180), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2181), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2182), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2183), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2184), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2185), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2186), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2187), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2188), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2189), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2190), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2191), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2192), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2193), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2194), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2195), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2196), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2197), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2198), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2199), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2200), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2201), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2202), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2203), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2204), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2205), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2206), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2207), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2208), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2209), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2210), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2211), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2212), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2213), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2214), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2215), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2216), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2217), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2218), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2219), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2220), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2221), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2222), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2223), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2224), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2225), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2226), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2227), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2228), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2229), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2230), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2231), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2232), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2233), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2234), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2235), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2236), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2237), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2238), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2239), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2240), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2241), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2242), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2243), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2244), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2245), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2246), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2247), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2248), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2249), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2250), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2251), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2252), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2253), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2254), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2255), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2256), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2257), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2258), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2259), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2260), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2261), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2262), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2263), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2264), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2265), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2266), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2267), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2268), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2269), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2270), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2271), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2272), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2273), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2274), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2275), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2276), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2277), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2278), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2279), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2280), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2281), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2282), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2283), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2284), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2285), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2286), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2287), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2288), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2289), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2290), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2291), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2292), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2293), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2294), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2295), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2296), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2297), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2298), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2299), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2300), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2301), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2302), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2303), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2304), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2305), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2306), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2307), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2308), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2309), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2310), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2311), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2312), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2313), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2314), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2315), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2316), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2317), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2318), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2319), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2320), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2321), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2322), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2323), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2324), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2325), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2326), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2327), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2328), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2329), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2330), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2331), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2332), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2333), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2334), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2335), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2336), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2337), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2338), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2339), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2340), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2341), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2342), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2343), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2344), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2345), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2346), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2347), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2348), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2349), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2350), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2351), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2352), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2353), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2354), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2355), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2356), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2357), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2358), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2359), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2360), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2361), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2362), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2363), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2364), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2365), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2366), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2367), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2368), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2369), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2370), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2371), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2372), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2373), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2374), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2375), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2376), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2377), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2378), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2379), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2380), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2381), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2382), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2383), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2384), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2385), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2386), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2387), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2388), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2389), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2390), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2391), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2392), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2393), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2394), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2395), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2396), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2397), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2398), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2399), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2400), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2401), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2402), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2403), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2404), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2405), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2406), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2407) );
  INVX1 U2 ( .A(n1168), .Y(N32) );
  INVX1 U3 ( .A(n1170), .Y(N30) );
  INVX1 U4 ( .A(n1171), .Y(N29) );
  INVX1 U5 ( .A(n1173), .Y(N27) );
  INVX1 U6 ( .A(n1176), .Y(N24) );
  INVX1 U7 ( .A(n1178), .Y(N22) );
  INVX1 U8 ( .A(n1179), .Y(N21) );
  INVX1 U9 ( .A(n1180), .Y(N20) );
  INVX1 U10 ( .A(n1183), .Y(N17) );
  INVX1 U11 ( .A(n1207), .Y(n1208) );
  INVX1 U12 ( .A(n1207), .Y(n1209) );
  INVX1 U13 ( .A(n1191), .Y(n1192) );
  INVX1 U14 ( .A(n1207), .Y(n1210) );
  INVX1 U15 ( .A(n1206), .Y(n1211) );
  INVX1 U16 ( .A(n1191), .Y(n1193) );
  INVX1 U17 ( .A(n1206), .Y(n1212) );
  INVX1 U18 ( .A(n1206), .Y(n1213) );
  INVX1 U19 ( .A(n1191), .Y(n1194) );
  INVX2 U20 ( .A(n1206), .Y(n1214) );
  INVX2 U21 ( .A(n1206), .Y(n1215) );
  INVX1 U22 ( .A(n1190), .Y(n1195) );
  INVX2 U23 ( .A(n1206), .Y(n1216) );
  INVX1 U24 ( .A(n1205), .Y(n1217) );
  INVX1 U25 ( .A(n1190), .Y(n1196) );
  INVX1 U26 ( .A(n1205), .Y(n1218) );
  INVX1 U27 ( .A(n1205), .Y(n1219) );
  INVX1 U28 ( .A(n1190), .Y(n1197) );
  INVX1 U29 ( .A(n1204), .Y(n1220) );
  INVX1 U30 ( .A(n1204), .Y(n1221) );
  INVX1 U31 ( .A(n1204), .Y(n1222) );
  INVX1 U32 ( .A(n1205), .Y(n1223) );
  INVX1 U33 ( .A(n1205), .Y(n1224) );
  INVX1 U34 ( .A(n1204), .Y(n1225) );
  INVX1 U35 ( .A(n1203), .Y(n1226) );
  INVX1 U36 ( .A(n1203), .Y(n1227) );
  INVX2 U37 ( .A(n1190), .Y(n1200) );
  INVX1 U38 ( .A(n1207), .Y(n1228) );
  INVX1 U39 ( .A(n1203), .Y(n1229) );
  INVX1 U40 ( .A(n1191), .Y(n1201) );
  INVX1 U41 ( .A(n1177), .Y(N23) );
  INVX1 U42 ( .A(n1169), .Y(N31) );
  INVX1 U43 ( .A(n1172), .Y(N28) );
  INVX1 U44 ( .A(n1174), .Y(N26) );
  INVX1 U45 ( .A(n1175), .Y(N25) );
  INVX1 U46 ( .A(n1181), .Y(N19) );
  INVX1 U47 ( .A(n1182), .Y(N18) );
  BUFX2 U48 ( .A(n102), .Y(n1231) );
  BUFX2 U49 ( .A(n104), .Y(n1233) );
  BUFX2 U50 ( .A(n106), .Y(n1235) );
  BUFX2 U51 ( .A(n108), .Y(n1237) );
  BUFX2 U52 ( .A(n110), .Y(n1239) );
  BUFX2 U53 ( .A(n112), .Y(n1241) );
  BUFX2 U54 ( .A(n114), .Y(n1243) );
  BUFX2 U55 ( .A(n116), .Y(n1248) );
  BUFX2 U56 ( .A(n118), .Y(n1250) );
  BUFX2 U57 ( .A(n120), .Y(n1254) );
  BUFX2 U58 ( .A(n122), .Y(n1258) );
  BUFX2 U59 ( .A(n124), .Y(n1262) );
  BUFX2 U60 ( .A(n127), .Y(n1264) );
  BUFX2 U61 ( .A(n130), .Y(n1266) );
  BUFX2 U62 ( .A(n133), .Y(n1271) );
  BUFX2 U63 ( .A(n135), .Y(n1275) );
  BUFX2 U64 ( .A(n137), .Y(n1279) );
  BUFX2 U65 ( .A(n139), .Y(n1283) );
  BUFX2 U66 ( .A(n141), .Y(n1287) );
  BUFX2 U67 ( .A(n143), .Y(n1291) );
  BUFX2 U68 ( .A(n145), .Y(n1295) );
  BUFX2 U69 ( .A(n147), .Y(n1302) );
  BUFX2 U70 ( .A(n149), .Y(n1306) );
  BUFX2 U71 ( .A(n152), .Y(n1308) );
  BUFX2 U72 ( .A(n155), .Y(n1310) );
  BUFX2 U73 ( .A(n158), .Y(n1312) );
  BUFX2 U74 ( .A(n161), .Y(n1314) );
  BUFX2 U75 ( .A(n164), .Y(n1316) );
  INVX2 U76 ( .A(n1202), .Y(n1198) );
  INVX1 U77 ( .A(n1202), .Y(n1199) );
  INVX1 U78 ( .A(n1358), .Y(n1186) );
  INVX1 U79 ( .A(n1358), .Y(n1185) );
  INVX1 U80 ( .A(N12), .Y(n1356) );
  INVX2 U81 ( .A(n1356), .Y(n1188) );
  INVX1 U82 ( .A(n1230), .Y(n1205) );
  INVX1 U83 ( .A(n1230), .Y(n1204) );
  INVX1 U84 ( .A(n1354), .Y(n1202) );
  INVX1 U85 ( .A(n1356), .Y(n1189) );
  INVX1 U86 ( .A(n1356), .Y(n1187) );
  INVX1 U87 ( .A(n1352), .Y(n1206) );
  INVX1 U88 ( .A(n99), .Y(n1299) );
  INVX1 U89 ( .A(n100), .Y(n1318) );
  BUFX2 U90 ( .A(n120), .Y(n1255) );
  BUFX2 U91 ( .A(n122), .Y(n1259) );
  BUFX2 U92 ( .A(n130), .Y(n1267) );
  BUFX2 U93 ( .A(n112), .Y(n1242) );
  BUFX2 U94 ( .A(n110), .Y(n1240) );
  BUFX2 U95 ( .A(n106), .Y(n1236) );
  BUFX2 U96 ( .A(n133), .Y(n1272) );
  BUFX2 U97 ( .A(n137), .Y(n1280) );
  BUFX2 U98 ( .A(n139), .Y(n1284) );
  BUFX2 U99 ( .A(n141), .Y(n1288) );
  BUFX2 U100 ( .A(n143), .Y(n1292) );
  BUFX2 U101 ( .A(n145), .Y(n1296) );
  BUFX2 U102 ( .A(n147), .Y(n1303) );
  INVX1 U103 ( .A(n1358), .Y(n1357) );
  INVX1 U104 ( .A(N13), .Y(n1358) );
  INVX1 U105 ( .A(N14), .Y(n1359) );
  INVX1 U106 ( .A(n1353), .Y(n1230) );
  INVX1 U107 ( .A(n1230), .Y(n1203) );
  INVX1 U108 ( .A(n1230), .Y(n1207) );
  BUFX2 U109 ( .A(n102), .Y(n1232) );
  BUFX2 U110 ( .A(n118), .Y(n1251) );
  BUFX2 U111 ( .A(n124), .Y(n1263) );
  BUFX2 U112 ( .A(n127), .Y(n1265) );
  BUFX2 U113 ( .A(n135), .Y(n1276) );
  BUFX2 U114 ( .A(n149), .Y(n1307) );
  BUFX2 U115 ( .A(n152), .Y(n1309) );
  BUFX2 U116 ( .A(n155), .Y(n1311) );
  BUFX2 U117 ( .A(n158), .Y(n1313) );
  BUFX2 U118 ( .A(n161), .Y(n1315) );
  BUFX2 U119 ( .A(n164), .Y(n1317) );
  BUFX2 U120 ( .A(n116), .Y(n1249) );
  BUFX2 U121 ( .A(n114), .Y(n1244) );
  BUFX2 U122 ( .A(n108), .Y(n1238) );
  BUFX2 U123 ( .A(n104), .Y(n1234) );
  INVX1 U124 ( .A(n97), .Y(n1245) );
  INVX1 U125 ( .A(n98), .Y(n1270) );
  INVX1 U126 ( .A(n1354), .Y(n1190) );
  INVX1 U127 ( .A(n1354), .Y(n1191) );
  INVX1 U128 ( .A(n1359), .Y(n1184) );
  INVX1 U129 ( .A(rst), .Y(n1351) );
  INVX4 U130 ( .A(n66), .Y(n166) );
  INVX4 U131 ( .A(n41), .Y(n131) );
  INVX4 U132 ( .A(n65), .Y(n165) );
  INVX4 U133 ( .A(n64), .Y(n162) );
  INVX4 U134 ( .A(n63), .Y(n159) );
  INVX4 U135 ( .A(n62), .Y(n156) );
  INVX4 U136 ( .A(n38), .Y(n128) );
  INVX4 U137 ( .A(n37), .Y(n125) );
  INVX4 U138 ( .A(n61), .Y(n153) );
  INVX4 U139 ( .A(n60), .Y(n150) );
  INVX1 U140 ( .A(n67), .Y(n1) );
  INVX1 U141 ( .A(n67), .Y(n2) );
  INVX1 U142 ( .A(n67), .Y(n3) );
  INVX1 U143 ( .A(n67), .Y(n4) );
  INVX1 U144 ( .A(n67), .Y(n5) );
  INVX1 U145 ( .A(n67), .Y(n6) );
  INVX1 U146 ( .A(n2), .Y(n7) );
  INVX1 U147 ( .A(n2), .Y(n8) );
  INVX1 U148 ( .A(n2), .Y(n9) );
  INVX1 U149 ( .A(n1), .Y(n10) );
  INVX1 U150 ( .A(n1), .Y(n11) );
  INVX1 U151 ( .A(n1), .Y(n12) );
  INVX1 U152 ( .A(n3), .Y(n13) );
  INVX1 U153 ( .A(n3), .Y(n14) );
  INVX1 U154 ( .A(n3), .Y(n15) );
  INVX1 U155 ( .A(n4), .Y(n16) );
  INVX1 U156 ( .A(n4), .Y(n17) );
  INVX1 U157 ( .A(n4), .Y(n18) );
  INVX1 U158 ( .A(n5), .Y(n19) );
  INVX1 U159 ( .A(n5), .Y(n20) );
  INVX1 U160 ( .A(n5), .Y(n21) );
  INVX1 U161 ( .A(n6), .Y(n22) );
  INVX1 U162 ( .A(n6), .Y(n23) );
  INVX1 U163 ( .A(n6), .Y(n24) );
  INVX1 U164 ( .A(n27), .Y(n25) );
  INVX2 U165 ( .A(n27), .Y(n26) );
  INVX2 U166 ( .A(n27), .Y(n28) );
  OR2X2 U167 ( .A(write), .B(rst), .Y(n27) );
  AND2X2 U168 ( .A(n19), .B(n97), .Y(n29) );
  INVX1 U169 ( .A(n29), .Y(n30) );
  AND2X2 U170 ( .A(n20), .B(n117), .Y(n31) );
  INVX1 U171 ( .A(n31), .Y(n32) );
  AND2X2 U172 ( .A(n21), .B(n119), .Y(n33) );
  INVX1 U173 ( .A(n33), .Y(n34) );
  AND2X2 U174 ( .A(n22), .B(n121), .Y(n35) );
  INVX1 U175 ( .A(n35), .Y(n36) );
  AND2X2 U176 ( .A(n14), .B(n123), .Y(n37) );
  AND2X2 U177 ( .A(n17), .B(n126), .Y(n38) );
  AND2X2 U178 ( .A(n7), .B(n129), .Y(n39) );
  INVX1 U179 ( .A(n39), .Y(n40) );
  AND2X2 U180 ( .A(n13), .B(n98), .Y(n41) );
  AND2X2 U181 ( .A(n8), .B(n132), .Y(n42) );
  INVX1 U182 ( .A(n42), .Y(n43) );
  AND2X2 U183 ( .A(n7), .B(n134), .Y(n44) );
  INVX1 U184 ( .A(n44), .Y(n45) );
  AND2X2 U185 ( .A(n8), .B(n136), .Y(n46) );
  INVX1 U186 ( .A(n46), .Y(n47) );
  AND2X2 U187 ( .A(n9), .B(n138), .Y(n48) );
  INVX1 U188 ( .A(n48), .Y(n49) );
  AND2X2 U189 ( .A(n10), .B(n140), .Y(n50) );
  INVX1 U190 ( .A(n50), .Y(n51) );
  AND2X2 U191 ( .A(n11), .B(n142), .Y(n52) );
  INVX1 U192 ( .A(n52), .Y(n53) );
  AND2X2 U193 ( .A(n12), .B(n144), .Y(n54) );
  INVX1 U194 ( .A(n54), .Y(n55) );
  AND2X2 U195 ( .A(n23), .B(n99), .Y(n56) );
  INVX1 U196 ( .A(n56), .Y(n57) );
  AND2X2 U197 ( .A(n24), .B(n146), .Y(n58) );
  INVX1 U198 ( .A(n58), .Y(n59) );
  AND2X2 U199 ( .A(n18), .B(n148), .Y(n60) );
  AND2X2 U200 ( .A(n14), .B(n151), .Y(n61) );
  AND2X2 U201 ( .A(n18), .B(n154), .Y(n62) );
  AND2X2 U202 ( .A(n17), .B(n157), .Y(n63) );
  AND2X2 U203 ( .A(n16), .B(n160), .Y(n64) );
  AND2X2 U204 ( .A(n18), .B(n163), .Y(n65) );
  AND2X2 U205 ( .A(n13), .B(n100), .Y(n66) );
  BUFX2 U206 ( .A(n40), .Y(n1268) );
  BUFX2 U207 ( .A(n40), .Y(n1269) );
  BUFX2 U208 ( .A(n43), .Y(n1273) );
  BUFX2 U209 ( .A(n43), .Y(n1274) );
  BUFX2 U210 ( .A(n45), .Y(n1277) );
  BUFX2 U211 ( .A(n45), .Y(n1278) );
  BUFX2 U212 ( .A(n47), .Y(n1281) );
  BUFX2 U213 ( .A(n47), .Y(n1282) );
  BUFX2 U214 ( .A(n49), .Y(n1285) );
  BUFX2 U215 ( .A(n49), .Y(n1286) );
  BUFX2 U216 ( .A(n51), .Y(n1289) );
  BUFX2 U217 ( .A(n51), .Y(n1290) );
  BUFX2 U218 ( .A(n53), .Y(n1293) );
  BUFX2 U219 ( .A(n53), .Y(n1294) );
  BUFX2 U220 ( .A(n55), .Y(n1297) );
  BUFX2 U221 ( .A(n55), .Y(n1298) );
  BUFX2 U222 ( .A(n57), .Y(n1300) );
  BUFX2 U223 ( .A(n57), .Y(n1301) );
  BUFX2 U224 ( .A(n59), .Y(n1304) );
  BUFX2 U225 ( .A(n59), .Y(n1305) );
  AND2X2 U226 ( .A(write), .B(n1351), .Y(n67) );
  AND2X2 U227 ( .A(\data_in<0> ), .B(n21), .Y(n68) );
  AND2X2 U228 ( .A(\data_in<1> ), .B(n18), .Y(n69) );
  AND2X2 U229 ( .A(\data_in<2> ), .B(n24), .Y(n70) );
  AND2X2 U230 ( .A(\data_in<3> ), .B(n18), .Y(n71) );
  AND2X2 U231 ( .A(\data_in<4> ), .B(n15), .Y(n72) );
  AND2X2 U232 ( .A(\data_in<5> ), .B(n19), .Y(n73) );
  AND2X2 U233 ( .A(\data_in<6> ), .B(n17), .Y(n74) );
  AND2X2 U234 ( .A(\data_in<7> ), .B(n20), .Y(n75) );
  AND2X2 U235 ( .A(\data_in<8> ), .B(n22), .Y(n76) );
  AND2X2 U236 ( .A(\data_in<9> ), .B(n23), .Y(n77) );
  AND2X2 U237 ( .A(\data_in<10> ), .B(n17), .Y(n78) );
  AND2X2 U238 ( .A(\data_in<11> ), .B(n14), .Y(n79) );
  AND2X2 U239 ( .A(\data_in<12> ), .B(n13), .Y(n80) );
  AND2X2 U240 ( .A(\data_in<13> ), .B(n15), .Y(n81) );
  AND2X2 U241 ( .A(\data_in<14> ), .B(n16), .Y(n82) );
  AND2X2 U242 ( .A(\data_in<15> ), .B(n17), .Y(n83) );
  INVX1 U243 ( .A(n1353), .Y(n1352) );
  AND2X1 U244 ( .A(n1187), .B(n1354), .Y(n84) );
  INVX1 U245 ( .A(n1355), .Y(n1354) );
  AND2X1 U246 ( .A(n2407), .B(N14), .Y(n85) );
  INVX2 U247 ( .A(n174), .Y(n1375) );
  INVX2 U248 ( .A(n173), .Y(n1392) );
  INVX2 U249 ( .A(n171), .Y(n1410) );
  INVX2 U250 ( .A(n172), .Y(n1428) );
  INVX2 U251 ( .A(n170), .Y(n1446) );
  INVX2 U252 ( .A(n169), .Y(n1464) );
  INVX2 U253 ( .A(n168), .Y(n1482) );
  INVX2 U254 ( .A(n167), .Y(n1515) );
  BUFX2 U255 ( .A(n1394), .Y(n86) );
  INVX1 U256 ( .A(n86), .Y(n1792) );
  BUFX2 U257 ( .A(n1412), .Y(n87) );
  INVX1 U258 ( .A(n87), .Y(n1809) );
  BUFX2 U259 ( .A(n1430), .Y(n88) );
  INVX1 U260 ( .A(n88), .Y(n1826) );
  BUFX2 U261 ( .A(n1448), .Y(n89) );
  INVX1 U262 ( .A(n89), .Y(n1843) );
  BUFX2 U263 ( .A(n1466), .Y(n90) );
  INVX1 U264 ( .A(n90), .Y(n1860) );
  BUFX2 U265 ( .A(n1629), .Y(n91) );
  INVX1 U266 ( .A(n91), .Y(n1742) );
  BUFX2 U267 ( .A(n1759), .Y(n92) );
  INVX1 U268 ( .A(n92), .Y(n1877) );
  AND2X1 U269 ( .A(n1352), .B(n84), .Y(n93) );
  AND2X1 U270 ( .A(n1357), .B(n85), .Y(n94) );
  AND2X1 U271 ( .A(n1353), .B(n84), .Y(n95) );
  AND2X1 U272 ( .A(n1358), .B(n85), .Y(n96) );
  AND2X1 U273 ( .A(n94), .B(n1878), .Y(n97) );
  AND2X1 U274 ( .A(n1878), .B(n96), .Y(n98) );
  AND2X1 U275 ( .A(n1878), .B(n1742), .Y(n99) );
  AND2X1 U276 ( .A(n1878), .B(n1877), .Y(n100) );
  AND2X1 U277 ( .A(n93), .B(n94), .Y(n101) );
  INVX1 U278 ( .A(n101), .Y(n102) );
  AND2X1 U279 ( .A(n94), .B(n95), .Y(n103) );
  INVX1 U280 ( .A(n103), .Y(n104) );
  AND2X1 U281 ( .A(n94), .B(n1792), .Y(n105) );
  INVX1 U282 ( .A(n105), .Y(n106) );
  AND2X1 U283 ( .A(n94), .B(n1809), .Y(n107) );
  INVX1 U284 ( .A(n107), .Y(n108) );
  AND2X1 U285 ( .A(n94), .B(n1826), .Y(n109) );
  INVX1 U286 ( .A(n109), .Y(n110) );
  AND2X1 U287 ( .A(n94), .B(n1843), .Y(n111) );
  INVX1 U288 ( .A(n111), .Y(n112) );
  AND2X1 U289 ( .A(n94), .B(n1860), .Y(n113) );
  INVX1 U290 ( .A(n113), .Y(n114) );
  AND2X1 U291 ( .A(n93), .B(n96), .Y(n115) );
  INVX1 U292 ( .A(n115), .Y(n116) );
  AND2X1 U293 ( .A(n95), .B(n96), .Y(n117) );
  INVX1 U294 ( .A(n117), .Y(n118) );
  AND2X1 U295 ( .A(n1792), .B(n96), .Y(n119) );
  INVX1 U296 ( .A(n119), .Y(n120) );
  AND2X1 U297 ( .A(n1809), .B(n96), .Y(n121) );
  INVX1 U298 ( .A(n121), .Y(n122) );
  AND2X1 U299 ( .A(n1826), .B(n96), .Y(n123) );
  INVX1 U300 ( .A(n123), .Y(n124) );
  AND2X1 U301 ( .A(n1843), .B(n96), .Y(n126) );
  INVX1 U302 ( .A(n126), .Y(n127) );
  AND2X1 U303 ( .A(n1860), .B(n96), .Y(n129) );
  INVX1 U304 ( .A(n129), .Y(n130) );
  AND2X1 U305 ( .A(n93), .B(n1742), .Y(n132) );
  INVX1 U306 ( .A(n132), .Y(n133) );
  AND2X1 U307 ( .A(n95), .B(n1742), .Y(n134) );
  INVX1 U308 ( .A(n134), .Y(n135) );
  AND2X1 U309 ( .A(n1792), .B(n1742), .Y(n136) );
  INVX1 U310 ( .A(n136), .Y(n137) );
  AND2X1 U311 ( .A(n1809), .B(n1742), .Y(n138) );
  INVX1 U312 ( .A(n138), .Y(n139) );
  AND2X1 U313 ( .A(n1826), .B(n1742), .Y(n140) );
  INVX1 U314 ( .A(n140), .Y(n141) );
  AND2X1 U315 ( .A(n1843), .B(n1742), .Y(n142) );
  INVX1 U316 ( .A(n142), .Y(n143) );
  AND2X1 U317 ( .A(n1860), .B(n1742), .Y(n144) );
  INVX1 U318 ( .A(n144), .Y(n145) );
  AND2X1 U319 ( .A(n93), .B(n1877), .Y(n146) );
  INVX1 U320 ( .A(n146), .Y(n147) );
  AND2X1 U321 ( .A(n95), .B(n1877), .Y(n148) );
  INVX1 U322 ( .A(n148), .Y(n149) );
  AND2X1 U323 ( .A(n1792), .B(n1877), .Y(n151) );
  INVX1 U324 ( .A(n151), .Y(n152) );
  AND2X1 U325 ( .A(n1809), .B(n1877), .Y(n154) );
  INVX1 U326 ( .A(n154), .Y(n155) );
  AND2X1 U327 ( .A(n1826), .B(n1877), .Y(n157) );
  INVX1 U328 ( .A(n157), .Y(n158) );
  AND2X1 U329 ( .A(n1843), .B(n1877), .Y(n160) );
  INVX1 U330 ( .A(n160), .Y(n161) );
  AND2X1 U331 ( .A(n1860), .B(n1877), .Y(n163) );
  INVX1 U332 ( .A(n163), .Y(n164) );
  BUFX2 U333 ( .A(n30), .Y(n1246) );
  BUFX2 U334 ( .A(n30), .Y(n1247) );
  BUFX2 U335 ( .A(n36), .Y(n1260) );
  BUFX2 U336 ( .A(n36), .Y(n1261) );
  BUFX2 U337 ( .A(n34), .Y(n1256) );
  BUFX2 U338 ( .A(n34), .Y(n1257) );
  BUFX2 U339 ( .A(n32), .Y(n1252) );
  BUFX2 U340 ( .A(n32), .Y(n1253) );
  AND2X2 U341 ( .A(n14), .B(n115), .Y(n167) );
  AND2X2 U342 ( .A(n15), .B(n113), .Y(n168) );
  AND2X2 U343 ( .A(n16), .B(n111), .Y(n169) );
  AND2X2 U344 ( .A(n9), .B(n109), .Y(n170) );
  AND2X2 U345 ( .A(n10), .B(n105), .Y(n171) );
  AND2X2 U346 ( .A(n11), .B(n107), .Y(n172) );
  AND2X2 U347 ( .A(n12), .B(n103), .Y(n173) );
  AND2X2 U348 ( .A(n13), .B(n101), .Y(n174) );
  INVX1 U349 ( .A(N11), .Y(n1355) );
  MUX2X1 U350 ( .B(n176), .A(n177), .S(n1192), .Y(n175) );
  MUX2X1 U351 ( .B(n179), .A(n180), .S(n1192), .Y(n178) );
  MUX2X1 U352 ( .B(n182), .A(n183), .S(n1192), .Y(n181) );
  MUX2X1 U353 ( .B(n185), .A(n186), .S(n1192), .Y(n184) );
  MUX2X1 U354 ( .B(n188), .A(n189), .S(n1186), .Y(n187) );
  MUX2X1 U355 ( .B(n191), .A(n192), .S(n1192), .Y(n190) );
  MUX2X1 U356 ( .B(n194), .A(n195), .S(n1192), .Y(n193) );
  MUX2X1 U357 ( .B(n197), .A(n198), .S(n1192), .Y(n196) );
  MUX2X1 U358 ( .B(n200), .A(n201), .S(n1192), .Y(n199) );
  MUX2X1 U359 ( .B(n203), .A(n204), .S(n1186), .Y(n202) );
  MUX2X1 U360 ( .B(n206), .A(n207), .S(n1193), .Y(n205) );
  MUX2X1 U361 ( .B(n209), .A(n210), .S(n1193), .Y(n208) );
  MUX2X1 U362 ( .B(n212), .A(n213), .S(n1193), .Y(n211) );
  MUX2X1 U363 ( .B(n216), .A(n217), .S(n1193), .Y(n215) );
  MUX2X1 U364 ( .B(n219), .A(n220), .S(n1186), .Y(n218) );
  MUX2X1 U365 ( .B(n222), .A(n223), .S(n1193), .Y(n221) );
  MUX2X1 U366 ( .B(n225), .A(n226), .S(n1193), .Y(n224) );
  MUX2X1 U367 ( .B(n228), .A(n229), .S(n1193), .Y(n227) );
  MUX2X1 U368 ( .B(n231), .A(n232), .S(n1193), .Y(n230) );
  MUX2X1 U369 ( .B(n234), .A(n235), .S(n1186), .Y(n233) );
  MUX2X1 U370 ( .B(n237), .A(n238), .S(n1193), .Y(n236) );
  MUX2X1 U371 ( .B(n240), .A(n241), .S(n1193), .Y(n239) );
  MUX2X1 U372 ( .B(n243), .A(n244), .S(n1193), .Y(n242) );
  MUX2X1 U373 ( .B(n246), .A(n247), .S(n1193), .Y(n245) );
  MUX2X1 U374 ( .B(n249), .A(n250), .S(n1186), .Y(n248) );
  MUX2X1 U375 ( .B(n252), .A(n253), .S(n1194), .Y(n251) );
  MUX2X1 U376 ( .B(n255), .A(n256), .S(n1194), .Y(n254) );
  MUX2X1 U377 ( .B(n258), .A(n259), .S(n1194), .Y(n257) );
  MUX2X1 U378 ( .B(n261), .A(n262), .S(n1194), .Y(n260) );
  MUX2X1 U379 ( .B(n264), .A(n265), .S(n1186), .Y(n263) );
  MUX2X1 U380 ( .B(n267), .A(n268), .S(n1194), .Y(n266) );
  MUX2X1 U381 ( .B(n270), .A(n271), .S(n1194), .Y(n269) );
  MUX2X1 U382 ( .B(n273), .A(n274), .S(n1194), .Y(n272) );
  MUX2X1 U383 ( .B(n276), .A(n277), .S(n1194), .Y(n275) );
  MUX2X1 U384 ( .B(n279), .A(n280), .S(n1186), .Y(n278) );
  MUX2X1 U385 ( .B(n282), .A(n283), .S(n1194), .Y(n281) );
  MUX2X1 U386 ( .B(n285), .A(n286), .S(n1194), .Y(n284) );
  MUX2X1 U387 ( .B(n288), .A(n289), .S(n1194), .Y(n287) );
  MUX2X1 U388 ( .B(n291), .A(n292), .S(n1194), .Y(n290) );
  MUX2X1 U389 ( .B(n294), .A(n295), .S(n1186), .Y(n293) );
  MUX2X1 U390 ( .B(n297), .A(n298), .S(n1195), .Y(n296) );
  MUX2X1 U391 ( .B(n300), .A(n301), .S(n1195), .Y(n299) );
  MUX2X1 U392 ( .B(n303), .A(n304), .S(n1195), .Y(n302) );
  MUX2X1 U393 ( .B(n306), .A(n307), .S(n1195), .Y(n305) );
  MUX2X1 U394 ( .B(n309), .A(n310), .S(n1186), .Y(n308) );
  MUX2X1 U395 ( .B(n312), .A(n313), .S(n1195), .Y(n311) );
  MUX2X1 U396 ( .B(n315), .A(n316), .S(n1195), .Y(n314) );
  MUX2X1 U397 ( .B(n318), .A(n319), .S(n1195), .Y(n317) );
  MUX2X1 U398 ( .B(n321), .A(n322), .S(n1195), .Y(n320) );
  MUX2X1 U399 ( .B(n324), .A(n325), .S(n1186), .Y(n323) );
  MUX2X1 U400 ( .B(n327), .A(n328), .S(n1195), .Y(n326) );
  MUX2X1 U401 ( .B(n330), .A(n331), .S(n1195), .Y(n329) );
  MUX2X1 U402 ( .B(n333), .A(n334), .S(n1195), .Y(n332) );
  MUX2X1 U403 ( .B(n336), .A(n337), .S(n1195), .Y(n335) );
  MUX2X1 U404 ( .B(n339), .A(n340), .S(n1186), .Y(n338) );
  MUX2X1 U405 ( .B(n342), .A(n343), .S(n1196), .Y(n341) );
  MUX2X1 U406 ( .B(n345), .A(n346), .S(n1196), .Y(n344) );
  MUX2X1 U407 ( .B(n348), .A(n349), .S(n1196), .Y(n347) );
  MUX2X1 U408 ( .B(n351), .A(n352), .S(n1196), .Y(n350) );
  MUX2X1 U409 ( .B(n354), .A(n355), .S(n1186), .Y(n353) );
  MUX2X1 U410 ( .B(n357), .A(n358), .S(n1196), .Y(n356) );
  MUX2X1 U411 ( .B(n360), .A(n361), .S(n1196), .Y(n359) );
  MUX2X1 U412 ( .B(n363), .A(n364), .S(n1196), .Y(n362) );
  MUX2X1 U413 ( .B(n366), .A(n367), .S(n1196), .Y(n365) );
  MUX2X1 U414 ( .B(n369), .A(n370), .S(n1185), .Y(n368) );
  MUX2X1 U415 ( .B(n372), .A(n373), .S(n1196), .Y(n371) );
  MUX2X1 U416 ( .B(n375), .A(n376), .S(n1196), .Y(n374) );
  MUX2X1 U417 ( .B(n378), .A(n379), .S(n1196), .Y(n377) );
  MUX2X1 U418 ( .B(n381), .A(n382), .S(n1196), .Y(n380) );
  MUX2X1 U419 ( .B(n384), .A(n385), .S(n1185), .Y(n383) );
  MUX2X1 U420 ( .B(n387), .A(n388), .S(n1197), .Y(n386) );
  MUX2X1 U421 ( .B(n390), .A(n391), .S(n1197), .Y(n389) );
  MUX2X1 U422 ( .B(n393), .A(n394), .S(n1197), .Y(n392) );
  MUX2X1 U423 ( .B(n396), .A(n397), .S(n1197), .Y(n395) );
  MUX2X1 U424 ( .B(n399), .A(n400), .S(n1185), .Y(n398) );
  MUX2X1 U425 ( .B(n402), .A(n403), .S(n1197), .Y(n401) );
  MUX2X1 U426 ( .B(n405), .A(n406), .S(n1197), .Y(n404) );
  MUX2X1 U427 ( .B(n408), .A(n409), .S(n1197), .Y(n407) );
  MUX2X1 U428 ( .B(n411), .A(n412), .S(n1197), .Y(n410) );
  MUX2X1 U429 ( .B(n414), .A(n415), .S(n1185), .Y(n413) );
  MUX2X1 U430 ( .B(n417), .A(n418), .S(n1197), .Y(n416) );
  MUX2X1 U431 ( .B(n420), .A(n421), .S(n1197), .Y(n419) );
  MUX2X1 U432 ( .B(n423), .A(n424), .S(n1197), .Y(n422) );
  MUX2X1 U433 ( .B(n426), .A(n427), .S(n1197), .Y(n425) );
  MUX2X1 U434 ( .B(n429), .A(n430), .S(n1185), .Y(n428) );
  MUX2X1 U435 ( .B(n432), .A(n433), .S(n1198), .Y(n431) );
  MUX2X1 U436 ( .B(n435), .A(n436), .S(n1198), .Y(n434) );
  MUX2X1 U437 ( .B(n438), .A(n439), .S(n1198), .Y(n437) );
  MUX2X1 U438 ( .B(n441), .A(n442), .S(n1198), .Y(n440) );
  MUX2X1 U439 ( .B(n444), .A(n445), .S(n1185), .Y(n443) );
  MUX2X1 U440 ( .B(n447), .A(n448), .S(n1198), .Y(n446) );
  MUX2X1 U441 ( .B(n450), .A(n451), .S(n1198), .Y(n449) );
  MUX2X1 U442 ( .B(n453), .A(n454), .S(n1198), .Y(n452) );
  MUX2X1 U443 ( .B(n456), .A(n457), .S(n1198), .Y(n455) );
  MUX2X1 U444 ( .B(n459), .A(n460), .S(n1185), .Y(n458) );
  MUX2X1 U445 ( .B(n462), .A(n463), .S(n1198), .Y(n461) );
  MUX2X1 U446 ( .B(n465), .A(n466), .S(n1198), .Y(n464) );
  MUX2X1 U447 ( .B(n468), .A(n469), .S(n1198), .Y(n467) );
  MUX2X1 U448 ( .B(n471), .A(n472), .S(n1198), .Y(n470) );
  MUX2X1 U449 ( .B(n474), .A(n475), .S(n1185), .Y(n473) );
  MUX2X1 U450 ( .B(n477), .A(n478), .S(n1199), .Y(n476) );
  MUX2X1 U451 ( .B(n480), .A(n481), .S(n1199), .Y(n479) );
  MUX2X1 U452 ( .B(n483), .A(n484), .S(n1199), .Y(n482) );
  MUX2X1 U453 ( .B(n486), .A(n487), .S(n1199), .Y(n485) );
  MUX2X1 U454 ( .B(n489), .A(n490), .S(n1185), .Y(n488) );
  MUX2X1 U455 ( .B(n492), .A(n493), .S(n1199), .Y(n491) );
  MUX2X1 U456 ( .B(n495), .A(n496), .S(n1199), .Y(n494) );
  MUX2X1 U457 ( .B(n498), .A(n499), .S(n1199), .Y(n497) );
  MUX2X1 U458 ( .B(n501), .A(n502), .S(n1199), .Y(n500) );
  MUX2X1 U459 ( .B(n504), .A(n505), .S(n1185), .Y(n503) );
  MUX2X1 U460 ( .B(n507), .A(n508), .S(n1199), .Y(n506) );
  MUX2X1 U461 ( .B(n510), .A(n511), .S(n1199), .Y(n509) );
  MUX2X1 U462 ( .B(n513), .A(n514), .S(n1199), .Y(n512) );
  MUX2X1 U463 ( .B(n516), .A(n517), .S(n1199), .Y(n515) );
  MUX2X1 U464 ( .B(n519), .A(n520), .S(n1185), .Y(n518) );
  MUX2X1 U465 ( .B(n522), .A(n523), .S(n1198), .Y(n521) );
  MUX2X1 U466 ( .B(n525), .A(n526), .S(n1198), .Y(n524) );
  MUX2X1 U467 ( .B(n528), .A(n529), .S(n1198), .Y(n527) );
  MUX2X1 U468 ( .B(n531), .A(n532), .S(n1198), .Y(n530) );
  MUX2X1 U469 ( .B(n534), .A(n535), .S(n1185), .Y(n533) );
  MUX2X1 U470 ( .B(n537), .A(n538), .S(n1199), .Y(n536) );
  MUX2X1 U471 ( .B(n540), .A(n541), .S(n1198), .Y(n539) );
  MUX2X1 U472 ( .B(n543), .A(n544), .S(n1198), .Y(n542) );
  MUX2X1 U473 ( .B(n546), .A(n547), .S(n1199), .Y(n545) );
  MUX2X1 U474 ( .B(n549), .A(n550), .S(n1185), .Y(n548) );
  MUX2X1 U475 ( .B(n552), .A(n553), .S(n1198), .Y(n551) );
  MUX2X1 U476 ( .B(n555), .A(n556), .S(n1198), .Y(n554) );
  MUX2X1 U477 ( .B(n558), .A(n559), .S(n1198), .Y(n557) );
  MUX2X1 U478 ( .B(n561), .A(n562), .S(n1198), .Y(n560) );
  MUX2X1 U479 ( .B(n564), .A(n565), .S(n1186), .Y(n563) );
  MUX2X1 U480 ( .B(n567), .A(n568), .S(n1200), .Y(n566) );
  MUX2X1 U481 ( .B(n570), .A(n571), .S(n1200), .Y(n569) );
  MUX2X1 U482 ( .B(n573), .A(n574), .S(n1200), .Y(n572) );
  MUX2X1 U483 ( .B(n576), .A(n577), .S(n1200), .Y(n575) );
  MUX2X1 U484 ( .B(n579), .A(n580), .S(n1185), .Y(n578) );
  MUX2X1 U485 ( .B(n582), .A(n583), .S(n1200), .Y(n581) );
  MUX2X1 U486 ( .B(n585), .A(n586), .S(n1200), .Y(n584) );
  MUX2X1 U487 ( .B(n588), .A(n589), .S(n1200), .Y(n587) );
  MUX2X1 U488 ( .B(n591), .A(n592), .S(n1200), .Y(n590) );
  MUX2X1 U489 ( .B(n594), .A(n595), .S(n1186), .Y(n593) );
  MUX2X1 U490 ( .B(n597), .A(n598), .S(n1200), .Y(n596) );
  MUX2X1 U491 ( .B(n600), .A(n601), .S(n1200), .Y(n599) );
  MUX2X1 U492 ( .B(n603), .A(n604), .S(n1200), .Y(n602) );
  MUX2X1 U493 ( .B(n606), .A(n607), .S(n1200), .Y(n605) );
  MUX2X1 U494 ( .B(n609), .A(n610), .S(n1186), .Y(n608) );
  MUX2X1 U495 ( .B(n612), .A(n613), .S(n1201), .Y(n611) );
  MUX2X1 U496 ( .B(n615), .A(n616), .S(n1201), .Y(n614) );
  MUX2X1 U497 ( .B(n618), .A(n619), .S(n1201), .Y(n617) );
  MUX2X1 U498 ( .B(n621), .A(n622), .S(n1201), .Y(n620) );
  MUX2X1 U499 ( .B(n624), .A(n625), .S(n1185), .Y(n623) );
  MUX2X1 U500 ( .B(n627), .A(n628), .S(n1201), .Y(n626) );
  MUX2X1 U501 ( .B(n630), .A(n631), .S(n1201), .Y(n629) );
  MUX2X1 U502 ( .B(n633), .A(n634), .S(n1201), .Y(n632) );
  MUX2X1 U503 ( .B(n636), .A(n637), .S(n1201), .Y(n635) );
  MUX2X1 U504 ( .B(n639), .A(n640), .S(n1185), .Y(n638) );
  MUX2X1 U505 ( .B(n642), .A(n643), .S(n1201), .Y(n641) );
  MUX2X1 U506 ( .B(n645), .A(n646), .S(n1201), .Y(n644) );
  MUX2X1 U507 ( .B(n648), .A(n649), .S(n1201), .Y(n647) );
  MUX2X1 U508 ( .B(n1163), .A(n1164), .S(n1201), .Y(n650) );
  MUX2X1 U509 ( .B(n1166), .A(n1167), .S(n1186), .Y(n1165) );
  MUX2X1 U510 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1208), .Y(n177) );
  MUX2X1 U511 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1208), .Y(n176) );
  MUX2X1 U512 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1208), .Y(n180) );
  MUX2X1 U513 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1208), .Y(n179) );
  MUX2X1 U514 ( .B(n178), .A(n175), .S(n1189), .Y(n189) );
  MUX2X1 U515 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1209), .Y(n183) );
  MUX2X1 U516 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1209), .Y(n182) );
  MUX2X1 U517 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1209), .Y(n186) );
  MUX2X1 U518 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1209), .Y(n185) );
  MUX2X1 U519 ( .B(n184), .A(n181), .S(n1189), .Y(n188) );
  MUX2X1 U520 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1209), .Y(n192) );
  MUX2X1 U521 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1209), .Y(n191) );
  MUX2X1 U522 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1209), .Y(n195) );
  MUX2X1 U523 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1209), .Y(n194) );
  MUX2X1 U524 ( .B(n193), .A(n190), .S(n1189), .Y(n204) );
  MUX2X1 U525 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1209), .Y(n198) );
  MUX2X1 U526 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1209), .Y(n197) );
  MUX2X1 U527 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1209), .Y(n201) );
  MUX2X1 U528 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1209), .Y(n200) );
  MUX2X1 U529 ( .B(n199), .A(n196), .S(n1189), .Y(n203) );
  MUX2X1 U530 ( .B(n202), .A(n187), .S(n1184), .Y(n1168) );
  MUX2X1 U531 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1210), .Y(n207) );
  MUX2X1 U532 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1210), .Y(n206) );
  MUX2X1 U533 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1210), .Y(n210) );
  MUX2X1 U534 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1210), .Y(n209) );
  MUX2X1 U535 ( .B(n208), .A(n205), .S(n1189), .Y(n220) );
  MUX2X1 U536 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1210), .Y(n213) );
  MUX2X1 U537 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1210), .Y(n212) );
  MUX2X1 U538 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1210), .Y(n217) );
  MUX2X1 U539 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1210), .Y(n216) );
  MUX2X1 U540 ( .B(n215), .A(n211), .S(n1189), .Y(n219) );
  MUX2X1 U541 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1210), .Y(n223) );
  MUX2X1 U542 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1210), .Y(n222) );
  MUX2X1 U543 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1210), .Y(n226) );
  MUX2X1 U544 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1210), .Y(n225) );
  MUX2X1 U545 ( .B(n224), .A(n221), .S(n1189), .Y(n235) );
  MUX2X1 U546 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1211), .Y(n229) );
  MUX2X1 U547 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1211), .Y(n228) );
  MUX2X1 U548 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1211), .Y(n232) );
  MUX2X1 U549 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1211), .Y(n231) );
  MUX2X1 U550 ( .B(n230), .A(n227), .S(n1189), .Y(n234) );
  MUX2X1 U551 ( .B(n233), .A(n218), .S(n1184), .Y(n1169) );
  MUX2X1 U552 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1211), .Y(n238) );
  MUX2X1 U553 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1211), .Y(n237) );
  MUX2X1 U554 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1211), .Y(n241) );
  MUX2X1 U555 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1211), .Y(n240) );
  MUX2X1 U556 ( .B(n239), .A(n236), .S(n1189), .Y(n250) );
  MUX2X1 U557 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1211), .Y(n244) );
  MUX2X1 U558 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1211), .Y(n243) );
  MUX2X1 U559 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1211), .Y(n247) );
  MUX2X1 U560 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1211), .Y(n246) );
  MUX2X1 U561 ( .B(n245), .A(n242), .S(n1189), .Y(n249) );
  MUX2X1 U562 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1212), .Y(n253) );
  MUX2X1 U563 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1212), .Y(n252) );
  MUX2X1 U564 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1212), .Y(n256) );
  MUX2X1 U565 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1212), .Y(n255) );
  MUX2X1 U566 ( .B(n254), .A(n251), .S(n1189), .Y(n265) );
  MUX2X1 U567 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1212), .Y(n259) );
  MUX2X1 U568 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1212), .Y(n258) );
  MUX2X1 U569 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1212), .Y(n262) );
  MUX2X1 U570 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1212), .Y(n261) );
  MUX2X1 U571 ( .B(n260), .A(n257), .S(n1189), .Y(n264) );
  MUX2X1 U572 ( .B(n263), .A(n248), .S(n1184), .Y(n1170) );
  MUX2X1 U573 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1212), .Y(n268) );
  MUX2X1 U574 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1212), .Y(n267) );
  MUX2X1 U575 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1212), .Y(n271) );
  MUX2X1 U576 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1212), .Y(n270) );
  MUX2X1 U577 ( .B(n269), .A(n266), .S(n1188), .Y(n280) );
  MUX2X1 U578 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1213), .Y(n274) );
  MUX2X1 U579 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1213), .Y(n273) );
  MUX2X1 U580 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1213), .Y(n277) );
  MUX2X1 U581 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1213), .Y(n276) );
  MUX2X1 U582 ( .B(n275), .A(n272), .S(n1188), .Y(n279) );
  MUX2X1 U583 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1213), .Y(n283) );
  MUX2X1 U584 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1213), .Y(n282) );
  MUX2X1 U585 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1213), .Y(n286) );
  MUX2X1 U586 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1213), .Y(n285) );
  MUX2X1 U587 ( .B(n284), .A(n281), .S(n1188), .Y(n295) );
  MUX2X1 U588 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1213), .Y(n289) );
  MUX2X1 U589 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1213), .Y(n288) );
  MUX2X1 U590 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1213), .Y(n292) );
  MUX2X1 U591 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1213), .Y(n291) );
  MUX2X1 U592 ( .B(n290), .A(n287), .S(n1188), .Y(n294) );
  MUX2X1 U593 ( .B(n293), .A(n278), .S(n1184), .Y(n1171) );
  MUX2X1 U594 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1214), .Y(n298) );
  MUX2X1 U595 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1214), .Y(n297) );
  MUX2X1 U596 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1214), .Y(n301) );
  MUX2X1 U597 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1214), .Y(n300) );
  MUX2X1 U598 ( .B(n299), .A(n296), .S(n1188), .Y(n310) );
  MUX2X1 U599 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1214), .Y(n304) );
  MUX2X1 U600 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1214), .Y(n303) );
  MUX2X1 U601 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1214), .Y(n307) );
  MUX2X1 U602 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1214), .Y(n306) );
  MUX2X1 U603 ( .B(n305), .A(n302), .S(n1188), .Y(n309) );
  MUX2X1 U604 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1214), .Y(n313) );
  MUX2X1 U605 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1214), .Y(n312) );
  MUX2X1 U606 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1214), .Y(n316) );
  MUX2X1 U607 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1214), .Y(n315) );
  MUX2X1 U608 ( .B(n314), .A(n311), .S(n1188), .Y(n325) );
  MUX2X1 U609 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1215), .Y(n319) );
  MUX2X1 U610 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1215), .Y(n318) );
  MUX2X1 U611 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1215), .Y(n322) );
  MUX2X1 U612 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1215), .Y(n321) );
  MUX2X1 U613 ( .B(n320), .A(n317), .S(n1188), .Y(n324) );
  MUX2X1 U614 ( .B(n323), .A(n308), .S(n1184), .Y(n1172) );
  MUX2X1 U615 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1215), .Y(n328) );
  MUX2X1 U616 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1215), .Y(n327) );
  MUX2X1 U617 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1215), .Y(n331) );
  MUX2X1 U618 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1215), .Y(n330) );
  MUX2X1 U619 ( .B(n329), .A(n326), .S(n1188), .Y(n340) );
  MUX2X1 U620 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1215), .Y(n334) );
  MUX2X1 U621 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1215), .Y(n333) );
  MUX2X1 U622 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1215), .Y(n337) );
  MUX2X1 U623 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1215), .Y(n336) );
  MUX2X1 U624 ( .B(n335), .A(n332), .S(n1188), .Y(n339) );
  MUX2X1 U625 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1216), .Y(n343) );
  MUX2X1 U626 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1216), .Y(n342) );
  MUX2X1 U627 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1216), .Y(n346) );
  MUX2X1 U628 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1216), .Y(n345) );
  MUX2X1 U629 ( .B(n344), .A(n341), .S(n1188), .Y(n355) );
  MUX2X1 U630 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1216), .Y(n349) );
  MUX2X1 U631 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1216), .Y(n348) );
  MUX2X1 U632 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1216), .Y(n352) );
  MUX2X1 U633 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1216), .Y(n351) );
  MUX2X1 U634 ( .B(n350), .A(n347), .S(n1188), .Y(n354) );
  MUX2X1 U635 ( .B(n353), .A(n338), .S(n1184), .Y(n1173) );
  MUX2X1 U636 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1216), .Y(n358) );
  MUX2X1 U637 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1216), .Y(n357) );
  MUX2X1 U638 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1216), .Y(n361) );
  MUX2X1 U639 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1216), .Y(n360) );
  MUX2X1 U640 ( .B(n359), .A(n356), .S(n1188), .Y(n370) );
  MUX2X1 U641 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1217), .Y(n364) );
  MUX2X1 U642 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1217), .Y(n363) );
  MUX2X1 U643 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1217), .Y(n367) );
  MUX2X1 U644 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1217), .Y(n366) );
  MUX2X1 U645 ( .B(n365), .A(n362), .S(n1188), .Y(n369) );
  MUX2X1 U646 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1217), .Y(n373) );
  MUX2X1 U647 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1217), .Y(n372) );
  MUX2X1 U648 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1217), .Y(n376) );
  MUX2X1 U649 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1217), .Y(n375) );
  MUX2X1 U650 ( .B(n374), .A(n371), .S(n1188), .Y(n385) );
  MUX2X1 U651 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1217), .Y(n379) );
  MUX2X1 U652 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1217), .Y(n378) );
  MUX2X1 U653 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1217), .Y(n382) );
  MUX2X1 U654 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1217), .Y(n381) );
  MUX2X1 U655 ( .B(n380), .A(n377), .S(n1188), .Y(n384) );
  MUX2X1 U656 ( .B(n383), .A(n368), .S(n1184), .Y(n1174) );
  MUX2X1 U657 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1218), .Y(n388) );
  MUX2X1 U658 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1218), .Y(n387) );
  MUX2X1 U659 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1218), .Y(n391) );
  MUX2X1 U660 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1218), .Y(n390) );
  MUX2X1 U661 ( .B(n389), .A(n386), .S(n1188), .Y(n400) );
  MUX2X1 U662 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1218), .Y(n394) );
  MUX2X1 U663 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1218), .Y(n393) );
  MUX2X1 U664 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1218), .Y(n397) );
  MUX2X1 U665 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1218), .Y(n396) );
  MUX2X1 U666 ( .B(n395), .A(n392), .S(n1188), .Y(n399) );
  MUX2X1 U667 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1218), .Y(n403) );
  MUX2X1 U668 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1218), .Y(n402) );
  MUX2X1 U669 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1218), .Y(n406) );
  MUX2X1 U670 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1218), .Y(n405) );
  MUX2X1 U671 ( .B(n404), .A(n401), .S(n1188), .Y(n415) );
  MUX2X1 U672 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1219), .Y(n409) );
  MUX2X1 U673 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1219), .Y(n408) );
  MUX2X1 U674 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1219), .Y(n412) );
  MUX2X1 U675 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1219), .Y(n411) );
  MUX2X1 U676 ( .B(n410), .A(n407), .S(n1188), .Y(n414) );
  MUX2X1 U677 ( .B(n413), .A(n398), .S(n1184), .Y(n1175) );
  MUX2X1 U678 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1219), .Y(n418) );
  MUX2X1 U679 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1219), .Y(n417) );
  MUX2X1 U680 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1219), .Y(n421) );
  MUX2X1 U681 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1219), .Y(n420) );
  MUX2X1 U682 ( .B(n419), .A(n416), .S(n1188), .Y(n430) );
  MUX2X1 U683 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1219), .Y(n424) );
  MUX2X1 U684 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1219), .Y(n423) );
  MUX2X1 U685 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1219), .Y(n427) );
  MUX2X1 U686 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1219), .Y(n426) );
  MUX2X1 U687 ( .B(n425), .A(n422), .S(n1188), .Y(n429) );
  MUX2X1 U688 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1220), .Y(n433) );
  MUX2X1 U689 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1220), .Y(n432) );
  MUX2X1 U690 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1220), .Y(n436) );
  MUX2X1 U691 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1220), .Y(n435) );
  MUX2X1 U692 ( .B(n434), .A(n431), .S(n1188), .Y(n445) );
  MUX2X1 U693 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1220), .Y(n439) );
  MUX2X1 U694 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1220), .Y(n438) );
  MUX2X1 U695 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1220), .Y(n442) );
  MUX2X1 U696 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1220), .Y(n441) );
  MUX2X1 U697 ( .B(n440), .A(n437), .S(n1188), .Y(n444) );
  MUX2X1 U698 ( .B(n443), .A(n428), .S(n1184), .Y(n1176) );
  MUX2X1 U699 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1220), .Y(n448) );
  MUX2X1 U700 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1220), .Y(n447) );
  MUX2X1 U701 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1220), .Y(n451) );
  MUX2X1 U702 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1220), .Y(n450) );
  MUX2X1 U703 ( .B(n449), .A(n446), .S(n1188), .Y(n460) );
  MUX2X1 U704 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1221), .Y(n454) );
  MUX2X1 U705 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1221), .Y(n453) );
  MUX2X1 U706 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1221), .Y(n457) );
  MUX2X1 U707 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1221), .Y(n456) );
  MUX2X1 U708 ( .B(n455), .A(n452), .S(n1188), .Y(n459) );
  MUX2X1 U709 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1221), .Y(n463) );
  MUX2X1 U710 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1221), .Y(n462) );
  MUX2X1 U711 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1221), .Y(n466) );
  MUX2X1 U712 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1221), .Y(n465) );
  MUX2X1 U713 ( .B(n464), .A(n461), .S(n1188), .Y(n475) );
  MUX2X1 U714 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1221), .Y(n469) );
  MUX2X1 U715 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1221), .Y(n468) );
  MUX2X1 U716 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1221), .Y(n472) );
  MUX2X1 U717 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1221), .Y(n471) );
  MUX2X1 U718 ( .B(n470), .A(n467), .S(n1189), .Y(n474) );
  MUX2X1 U719 ( .B(n473), .A(n458), .S(n1184), .Y(n1177) );
  MUX2X1 U720 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1222), .Y(n478) );
  MUX2X1 U721 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1222), .Y(n477) );
  MUX2X1 U722 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1222), .Y(n481) );
  MUX2X1 U723 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1222), .Y(n480) );
  MUX2X1 U724 ( .B(n479), .A(n476), .S(n1188), .Y(n490) );
  MUX2X1 U725 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1222), .Y(n484) );
  MUX2X1 U726 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1222), .Y(n483) );
  MUX2X1 U727 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1222), .Y(n487) );
  MUX2X1 U728 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1222), .Y(n486) );
  MUX2X1 U729 ( .B(n485), .A(n482), .S(n1188), .Y(n489) );
  MUX2X1 U730 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1222), .Y(n493) );
  MUX2X1 U731 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1222), .Y(n492) );
  MUX2X1 U732 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1222), .Y(n496) );
  MUX2X1 U733 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1222), .Y(n495) );
  MUX2X1 U734 ( .B(n494), .A(n491), .S(n1188), .Y(n505) );
  MUX2X1 U735 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1223), .Y(n499) );
  MUX2X1 U736 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1223), .Y(n498) );
  MUX2X1 U737 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1223), .Y(n502) );
  MUX2X1 U738 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1223), .Y(n501) );
  MUX2X1 U739 ( .B(n500), .A(n497), .S(n1188), .Y(n504) );
  MUX2X1 U740 ( .B(n503), .A(n488), .S(n1184), .Y(n1178) );
  MUX2X1 U741 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1223), .Y(n508) );
  MUX2X1 U742 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1223), .Y(n507) );
  MUX2X1 U743 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1223), .Y(n511) );
  MUX2X1 U744 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1223), .Y(n510) );
  MUX2X1 U745 ( .B(n509), .A(n506), .S(n1188), .Y(n520) );
  MUX2X1 U746 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1223), .Y(n514) );
  MUX2X1 U747 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1223), .Y(n513) );
  MUX2X1 U748 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1223), .Y(n517) );
  MUX2X1 U749 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1223), .Y(n516) );
  MUX2X1 U750 ( .B(n515), .A(n512), .S(n1189), .Y(n519) );
  MUX2X1 U751 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1224), .Y(n523) );
  MUX2X1 U752 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1224), .Y(n522) );
  MUX2X1 U753 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1224), .Y(n526) );
  MUX2X1 U754 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1224), .Y(n525) );
  MUX2X1 U755 ( .B(n524), .A(n521), .S(n1188), .Y(n535) );
  MUX2X1 U756 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1224), .Y(n529) );
  MUX2X1 U757 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1224), .Y(n528) );
  MUX2X1 U758 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1224), .Y(n532) );
  MUX2X1 U759 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1224), .Y(n531) );
  MUX2X1 U760 ( .B(n530), .A(n527), .S(n1188), .Y(n534) );
  MUX2X1 U761 ( .B(n533), .A(n518), .S(n1184), .Y(n1179) );
  MUX2X1 U762 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1224), .Y(n538) );
  MUX2X1 U763 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1224), .Y(n537) );
  MUX2X1 U764 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1224), .Y(n541) );
  MUX2X1 U765 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1224), .Y(n540) );
  MUX2X1 U766 ( .B(n539), .A(n536), .S(n1187), .Y(n550) );
  MUX2X1 U767 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1225), .Y(n544) );
  MUX2X1 U768 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1225), .Y(n543) );
  MUX2X1 U769 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1225), .Y(n547) );
  MUX2X1 U770 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1225), .Y(n546) );
  MUX2X1 U771 ( .B(n545), .A(n542), .S(n1187), .Y(n549) );
  MUX2X1 U772 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1225), .Y(n553) );
  MUX2X1 U773 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1225), .Y(n552) );
  MUX2X1 U774 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1225), .Y(n556) );
  MUX2X1 U775 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1225), .Y(n555) );
  MUX2X1 U776 ( .B(n554), .A(n551), .S(n1187), .Y(n565) );
  MUX2X1 U777 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1225), .Y(n559) );
  MUX2X1 U778 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1225), .Y(n558) );
  MUX2X1 U779 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1225), .Y(n562) );
  MUX2X1 U780 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1225), .Y(n561) );
  MUX2X1 U781 ( .B(n560), .A(n557), .S(n1187), .Y(n564) );
  MUX2X1 U782 ( .B(n563), .A(n548), .S(n1184), .Y(n1180) );
  MUX2X1 U783 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1226), .Y(n568) );
  MUX2X1 U784 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1226), .Y(n567) );
  MUX2X1 U785 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1226), .Y(n571) );
  MUX2X1 U786 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1226), .Y(n570) );
  MUX2X1 U787 ( .B(n569), .A(n566), .S(n1187), .Y(n580) );
  MUX2X1 U788 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1226), .Y(n574) );
  MUX2X1 U789 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1226), .Y(n573) );
  MUX2X1 U790 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1226), .Y(n577) );
  MUX2X1 U791 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1226), .Y(n576) );
  MUX2X1 U792 ( .B(n575), .A(n572), .S(n1187), .Y(n579) );
  MUX2X1 U793 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1226), .Y(n583) );
  MUX2X1 U794 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1226), .Y(n582) );
  MUX2X1 U795 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1226), .Y(n586) );
  MUX2X1 U796 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1226), .Y(n585) );
  MUX2X1 U797 ( .B(n584), .A(n581), .S(n1187), .Y(n595) );
  MUX2X1 U798 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1227), .Y(n589) );
  MUX2X1 U799 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1227), .Y(n588) );
  MUX2X1 U800 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1227), .Y(n592) );
  MUX2X1 U801 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1227), .Y(n591) );
  MUX2X1 U802 ( .B(n590), .A(n587), .S(n1187), .Y(n594) );
  MUX2X1 U803 ( .B(n593), .A(n578), .S(n1184), .Y(n1181) );
  MUX2X1 U804 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1227), .Y(n598) );
  MUX2X1 U805 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1227), .Y(n597) );
  MUX2X1 U806 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1227), .Y(n601) );
  MUX2X1 U807 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1227), .Y(n600) );
  MUX2X1 U808 ( .B(n599), .A(n596), .S(n1187), .Y(n610) );
  MUX2X1 U809 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1227), .Y(n604) );
  MUX2X1 U810 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1227), .Y(n603) );
  MUX2X1 U811 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1227), .Y(n607) );
  MUX2X1 U812 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1227), .Y(n606) );
  MUX2X1 U813 ( .B(n605), .A(n602), .S(n1187), .Y(n609) );
  MUX2X1 U814 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1228), .Y(n613) );
  MUX2X1 U815 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1228), .Y(n612) );
  MUX2X1 U816 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1228), .Y(n616) );
  MUX2X1 U817 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1228), .Y(n615) );
  MUX2X1 U818 ( .B(n614), .A(n611), .S(n1187), .Y(n625) );
  MUX2X1 U819 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1228), .Y(n619) );
  MUX2X1 U820 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1228), .Y(n618) );
  MUX2X1 U821 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1228), .Y(n622) );
  MUX2X1 U822 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1228), .Y(n621) );
  MUX2X1 U823 ( .B(n620), .A(n617), .S(n1187), .Y(n624) );
  MUX2X1 U824 ( .B(n623), .A(n608), .S(n1184), .Y(n1182) );
  MUX2X1 U825 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1228), .Y(n628) );
  MUX2X1 U826 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1228), .Y(n627) );
  MUX2X1 U827 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1228), .Y(n631) );
  MUX2X1 U828 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1228), .Y(n630) );
  MUX2X1 U829 ( .B(n629), .A(n626), .S(n1189), .Y(n640) );
  MUX2X1 U830 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1229), .Y(n634) );
  MUX2X1 U831 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1229), .Y(n633) );
  MUX2X1 U832 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1229), .Y(n637) );
  MUX2X1 U833 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1229), .Y(n636) );
  MUX2X1 U834 ( .B(n635), .A(n632), .S(n1187), .Y(n639) );
  MUX2X1 U835 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1229), .Y(n643) );
  MUX2X1 U836 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1229), .Y(n642) );
  MUX2X1 U837 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1229), .Y(n646) );
  MUX2X1 U838 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1229), .Y(n645) );
  MUX2X1 U839 ( .B(n644), .A(n641), .S(n1189), .Y(n1167) );
  MUX2X1 U840 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1229), .Y(n649) );
  MUX2X1 U841 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1229), .Y(n648) );
  MUX2X1 U842 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1229), .Y(n1164) );
  MUX2X1 U843 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1229), .Y(n1163) );
  MUX2X1 U844 ( .B(n650), .A(n647), .S(n1189), .Y(n1166) );
  MUX2X1 U845 ( .B(n1165), .A(n638), .S(n1184), .Y(n1183) );
  INVX1 U846 ( .A(N10), .Y(n1353) );
  INVX8 U847 ( .A(n68), .Y(n1319) );
  INVX8 U848 ( .A(n68), .Y(n1320) );
  INVX8 U849 ( .A(n69), .Y(n1321) );
  INVX8 U850 ( .A(n69), .Y(n1322) );
  INVX8 U851 ( .A(n70), .Y(n1323) );
  INVX8 U852 ( .A(n70), .Y(n1324) );
  INVX8 U853 ( .A(n71), .Y(n1325) );
  INVX8 U854 ( .A(n71), .Y(n1326) );
  INVX8 U855 ( .A(n72), .Y(n1327) );
  INVX8 U856 ( .A(n72), .Y(n1328) );
  INVX8 U857 ( .A(n73), .Y(n1329) );
  INVX8 U858 ( .A(n73), .Y(n1330) );
  INVX8 U859 ( .A(n74), .Y(n1331) );
  INVX8 U860 ( .A(n74), .Y(n1332) );
  INVX8 U861 ( .A(n75), .Y(n1333) );
  INVX8 U862 ( .A(n75), .Y(n1334) );
  INVX8 U863 ( .A(n76), .Y(n1335) );
  INVX8 U864 ( .A(n76), .Y(n1336) );
  INVX8 U865 ( .A(n77), .Y(n1337) );
  INVX8 U866 ( .A(n77), .Y(n1338) );
  INVX8 U867 ( .A(n78), .Y(n1339) );
  INVX8 U868 ( .A(n78), .Y(n1340) );
  INVX8 U869 ( .A(n79), .Y(n1341) );
  INVX8 U870 ( .A(n79), .Y(n1342) );
  INVX8 U871 ( .A(n80), .Y(n1343) );
  INVX8 U872 ( .A(n80), .Y(n1344) );
  INVX8 U873 ( .A(n81), .Y(n1345) );
  INVX8 U874 ( .A(n81), .Y(n1346) );
  INVX8 U875 ( .A(n82), .Y(n1347) );
  INVX8 U876 ( .A(n82), .Y(n1348) );
  INVX8 U877 ( .A(n83), .Y(n1349) );
  INVX8 U878 ( .A(n83), .Y(n1350) );
  AND2X2 U879 ( .A(N32), .B(n26), .Y(\data_out<0> ) );
  AND2X2 U880 ( .A(N31), .B(n28), .Y(\data_out<1> ) );
  AND2X2 U881 ( .A(n26), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U882 ( .A(N29), .B(n28), .Y(\data_out<3> ) );
  AND2X2 U883 ( .A(n25), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U884 ( .A(N27), .B(n28), .Y(\data_out<5> ) );
  AND2X2 U885 ( .A(n26), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U886 ( .A(n26), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U887 ( .A(N24), .B(n26), .Y(\data_out<8> ) );
  AND2X2 U888 ( .A(N23), .B(n28), .Y(\data_out<9> ) );
  AND2X2 U889 ( .A(n25), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U890 ( .A(N21), .B(n28), .Y(\data_out<11> ) );
  AND2X2 U891 ( .A(N20), .B(n26), .Y(\data_out<12> ) );
  AND2X2 U892 ( .A(n25), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U893 ( .A(N18), .B(n28), .Y(\data_out<14> ) );
  AND2X2 U894 ( .A(n26), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U895 ( .A(\mem<31><0> ), .B(n1375), .Y(n1360) );
  OAI21X1 U896 ( .A(n1232), .B(n1319), .C(n1360), .Y(n2406) );
  NAND2X1 U897 ( .A(\mem<31><1> ), .B(n1375), .Y(n1361) );
  OAI21X1 U898 ( .A(n1322), .B(n1231), .C(n1361), .Y(n2405) );
  NAND2X1 U899 ( .A(\mem<31><2> ), .B(n1375), .Y(n1362) );
  OAI21X1 U900 ( .A(n1324), .B(n1231), .C(n1362), .Y(n2404) );
  NAND2X1 U901 ( .A(\mem<31><3> ), .B(n1375), .Y(n1363) );
  OAI21X1 U902 ( .A(n1326), .B(n1231), .C(n1363), .Y(n2403) );
  NAND2X1 U903 ( .A(\mem<31><4> ), .B(n1375), .Y(n1364) );
  OAI21X1 U904 ( .A(n1328), .B(n1231), .C(n1364), .Y(n2402) );
  NAND2X1 U905 ( .A(\mem<31><5> ), .B(n1375), .Y(n1365) );
  OAI21X1 U906 ( .A(n1330), .B(n1231), .C(n1365), .Y(n2401) );
  NAND2X1 U907 ( .A(\mem<31><6> ), .B(n1375), .Y(n1366) );
  OAI21X1 U908 ( .A(n1332), .B(n1231), .C(n1366), .Y(n2400) );
  NAND2X1 U909 ( .A(\mem<31><7> ), .B(n1375), .Y(n1367) );
  OAI21X1 U910 ( .A(n1334), .B(n1231), .C(n1367), .Y(n2399) );
  NAND2X1 U911 ( .A(\mem<31><8> ), .B(n1375), .Y(n1368) );
  OAI21X1 U912 ( .A(n1336), .B(n1231), .C(n1368), .Y(n2398) );
  NAND2X1 U913 ( .A(\mem<31><9> ), .B(n1375), .Y(n1369) );
  OAI21X1 U914 ( .A(n1338), .B(n1232), .C(n1369), .Y(n2397) );
  NAND2X1 U915 ( .A(\mem<31><10> ), .B(n1375), .Y(n1370) );
  OAI21X1 U916 ( .A(n1340), .B(n1232), .C(n1370), .Y(n2396) );
  NAND2X1 U917 ( .A(\mem<31><11> ), .B(n1375), .Y(n1371) );
  OAI21X1 U918 ( .A(n1342), .B(n1232), .C(n1371), .Y(n2395) );
  NAND2X1 U919 ( .A(\mem<31><12> ), .B(n1375), .Y(n1372) );
  OAI21X1 U920 ( .A(n1344), .B(n1232), .C(n1372), .Y(n2394) );
  NAND2X1 U921 ( .A(\mem<31><13> ), .B(n1375), .Y(n1373) );
  OAI21X1 U922 ( .A(n1346), .B(n1232), .C(n1373), .Y(n2393) );
  NAND2X1 U923 ( .A(\mem<31><14> ), .B(n1375), .Y(n1374) );
  OAI21X1 U924 ( .A(n1348), .B(n1232), .C(n1374), .Y(n2392) );
  NAND2X1 U925 ( .A(\mem<31><15> ), .B(n1375), .Y(n1376) );
  OAI21X1 U926 ( .A(n1350), .B(n1232), .C(n1376), .Y(n2391) );
  NAND2X1 U927 ( .A(\mem<30><0> ), .B(n1392), .Y(n1377) );
  OAI21X1 U928 ( .A(n1233), .B(n1319), .C(n1377), .Y(n2390) );
  NAND2X1 U929 ( .A(\mem<30><1> ), .B(n1392), .Y(n1378) );
  OAI21X1 U930 ( .A(n1233), .B(n1322), .C(n1378), .Y(n2389) );
  NAND2X1 U931 ( .A(\mem<30><2> ), .B(n1392), .Y(n1379) );
  OAI21X1 U932 ( .A(n1233), .B(n1324), .C(n1379), .Y(n2388) );
  NAND2X1 U933 ( .A(\mem<30><3> ), .B(n1392), .Y(n1380) );
  OAI21X1 U934 ( .A(n1233), .B(n1326), .C(n1380), .Y(n2387) );
  NAND2X1 U935 ( .A(\mem<30><4> ), .B(n1392), .Y(n1381) );
  OAI21X1 U936 ( .A(n1233), .B(n1328), .C(n1381), .Y(n2386) );
  NAND2X1 U937 ( .A(\mem<30><5> ), .B(n1392), .Y(n1382) );
  OAI21X1 U938 ( .A(n1233), .B(n1330), .C(n1382), .Y(n2385) );
  NAND2X1 U939 ( .A(\mem<30><6> ), .B(n1392), .Y(n1383) );
  OAI21X1 U940 ( .A(n1233), .B(n1332), .C(n1383), .Y(n2384) );
  NAND2X1 U941 ( .A(\mem<30><7> ), .B(n1392), .Y(n1384) );
  OAI21X1 U942 ( .A(n1233), .B(n1334), .C(n1384), .Y(n2383) );
  NAND2X1 U943 ( .A(\mem<30><8> ), .B(n1392), .Y(n1385) );
  OAI21X1 U944 ( .A(n1234), .B(n1336), .C(n1385), .Y(n2382) );
  NAND2X1 U945 ( .A(\mem<30><9> ), .B(n1392), .Y(n1386) );
  OAI21X1 U946 ( .A(n1234), .B(n1338), .C(n1386), .Y(n2381) );
  NAND2X1 U947 ( .A(\mem<30><10> ), .B(n1392), .Y(n1387) );
  OAI21X1 U948 ( .A(n1234), .B(n1340), .C(n1387), .Y(n2380) );
  NAND2X1 U949 ( .A(\mem<30><11> ), .B(n1392), .Y(n1388) );
  OAI21X1 U950 ( .A(n1234), .B(n1342), .C(n1388), .Y(n2379) );
  NAND2X1 U951 ( .A(\mem<30><12> ), .B(n1392), .Y(n1389) );
  OAI21X1 U952 ( .A(n1234), .B(n1344), .C(n1389), .Y(n2378) );
  NAND2X1 U953 ( .A(\mem<30><13> ), .B(n1392), .Y(n1390) );
  OAI21X1 U954 ( .A(n1234), .B(n1346), .C(n1390), .Y(n2377) );
  NAND2X1 U955 ( .A(\mem<30><14> ), .B(n1392), .Y(n1391) );
  OAI21X1 U956 ( .A(n1234), .B(n1348), .C(n1391), .Y(n2376) );
  NAND2X1 U957 ( .A(\mem<30><15> ), .B(n1392), .Y(n1393) );
  OAI21X1 U958 ( .A(n1234), .B(n1350), .C(n1393), .Y(n2375) );
  NAND3X1 U959 ( .A(n1352), .B(n1187), .C(n1355), .Y(n1394) );
  NAND2X1 U960 ( .A(\mem<29><0> ), .B(n1410), .Y(n1395) );
  OAI21X1 U961 ( .A(n1235), .B(n1319), .C(n1395), .Y(n2374) );
  NAND2X1 U962 ( .A(\mem<29><1> ), .B(n1410), .Y(n1396) );
  OAI21X1 U963 ( .A(n1235), .B(n1322), .C(n1396), .Y(n2373) );
  NAND2X1 U964 ( .A(\mem<29><2> ), .B(n1410), .Y(n1397) );
  OAI21X1 U965 ( .A(n1235), .B(n1324), .C(n1397), .Y(n2372) );
  NAND2X1 U966 ( .A(\mem<29><3> ), .B(n1410), .Y(n1398) );
  OAI21X1 U967 ( .A(n1235), .B(n1326), .C(n1398), .Y(n2371) );
  NAND2X1 U968 ( .A(\mem<29><4> ), .B(n1410), .Y(n1399) );
  OAI21X1 U969 ( .A(n1235), .B(n1328), .C(n1399), .Y(n2370) );
  NAND2X1 U970 ( .A(\mem<29><5> ), .B(n1410), .Y(n1400) );
  OAI21X1 U971 ( .A(n1235), .B(n1330), .C(n1400), .Y(n2369) );
  NAND2X1 U972 ( .A(\mem<29><6> ), .B(n1410), .Y(n1401) );
  OAI21X1 U973 ( .A(n1235), .B(n1332), .C(n1401), .Y(n2368) );
  NAND2X1 U974 ( .A(\mem<29><7> ), .B(n1410), .Y(n1402) );
  OAI21X1 U975 ( .A(n1235), .B(n1334), .C(n1402), .Y(n2367) );
  NAND2X1 U976 ( .A(\mem<29><8> ), .B(n1410), .Y(n1403) );
  OAI21X1 U977 ( .A(n1236), .B(n1336), .C(n1403), .Y(n2366) );
  NAND2X1 U978 ( .A(\mem<29><9> ), .B(n1410), .Y(n1404) );
  OAI21X1 U979 ( .A(n1236), .B(n1338), .C(n1404), .Y(n2365) );
  NAND2X1 U980 ( .A(\mem<29><10> ), .B(n1410), .Y(n1405) );
  OAI21X1 U981 ( .A(n1236), .B(n1340), .C(n1405), .Y(n2364) );
  NAND2X1 U982 ( .A(\mem<29><11> ), .B(n1410), .Y(n1406) );
  OAI21X1 U983 ( .A(n1236), .B(n1342), .C(n1406), .Y(n2363) );
  NAND2X1 U984 ( .A(\mem<29><12> ), .B(n1410), .Y(n1407) );
  OAI21X1 U985 ( .A(n1236), .B(n1344), .C(n1407), .Y(n2362) );
  NAND2X1 U986 ( .A(\mem<29><13> ), .B(n1410), .Y(n1408) );
  OAI21X1 U987 ( .A(n1236), .B(n1346), .C(n1408), .Y(n2361) );
  NAND2X1 U988 ( .A(\mem<29><14> ), .B(n1410), .Y(n1409) );
  OAI21X1 U989 ( .A(n1236), .B(n1348), .C(n1409), .Y(n2360) );
  NAND2X1 U990 ( .A(\mem<29><15> ), .B(n1410), .Y(n1411) );
  OAI21X1 U991 ( .A(n1236), .B(n1350), .C(n1411), .Y(n2359) );
  NAND3X1 U992 ( .A(n1187), .B(n1355), .C(n1353), .Y(n1412) );
  NAND2X1 U993 ( .A(\mem<28><0> ), .B(n1428), .Y(n1413) );
  OAI21X1 U994 ( .A(n1237), .B(n1319), .C(n1413), .Y(n2358) );
  NAND2X1 U995 ( .A(\mem<28><1> ), .B(n1428), .Y(n1414) );
  OAI21X1 U996 ( .A(n1237), .B(n1322), .C(n1414), .Y(n2357) );
  NAND2X1 U997 ( .A(\mem<28><2> ), .B(n1428), .Y(n1415) );
  OAI21X1 U998 ( .A(n1237), .B(n1324), .C(n1415), .Y(n2356) );
  NAND2X1 U999 ( .A(\mem<28><3> ), .B(n1428), .Y(n1416) );
  OAI21X1 U1000 ( .A(n1237), .B(n1326), .C(n1416), .Y(n2355) );
  NAND2X1 U1001 ( .A(\mem<28><4> ), .B(n1428), .Y(n1417) );
  OAI21X1 U1002 ( .A(n1237), .B(n1328), .C(n1417), .Y(n2354) );
  NAND2X1 U1003 ( .A(\mem<28><5> ), .B(n1428), .Y(n1418) );
  OAI21X1 U1004 ( .A(n1237), .B(n1330), .C(n1418), .Y(n2353) );
  NAND2X1 U1005 ( .A(\mem<28><6> ), .B(n1428), .Y(n1419) );
  OAI21X1 U1006 ( .A(n1237), .B(n1332), .C(n1419), .Y(n2352) );
  NAND2X1 U1007 ( .A(\mem<28><7> ), .B(n1428), .Y(n1420) );
  OAI21X1 U1008 ( .A(n1237), .B(n1334), .C(n1420), .Y(n2351) );
  NAND2X1 U1009 ( .A(\mem<28><8> ), .B(n1428), .Y(n1421) );
  OAI21X1 U1010 ( .A(n1238), .B(n1336), .C(n1421), .Y(n2350) );
  NAND2X1 U1011 ( .A(\mem<28><9> ), .B(n1428), .Y(n1422) );
  OAI21X1 U1012 ( .A(n1238), .B(n1338), .C(n1422), .Y(n2349) );
  NAND2X1 U1013 ( .A(\mem<28><10> ), .B(n1428), .Y(n1423) );
  OAI21X1 U1014 ( .A(n1238), .B(n1340), .C(n1423), .Y(n2348) );
  NAND2X1 U1015 ( .A(\mem<28><11> ), .B(n1428), .Y(n1424) );
  OAI21X1 U1016 ( .A(n1238), .B(n1342), .C(n1424), .Y(n2347) );
  NAND2X1 U1017 ( .A(\mem<28><12> ), .B(n1428), .Y(n1425) );
  OAI21X1 U1018 ( .A(n1238), .B(n1344), .C(n1425), .Y(n2346) );
  NAND2X1 U1019 ( .A(\mem<28><13> ), .B(n1428), .Y(n1426) );
  OAI21X1 U1020 ( .A(n1238), .B(n1346), .C(n1426), .Y(n2345) );
  NAND2X1 U1021 ( .A(\mem<28><14> ), .B(n1428), .Y(n1427) );
  OAI21X1 U1022 ( .A(n1238), .B(n1348), .C(n1427), .Y(n2344) );
  NAND2X1 U1023 ( .A(\mem<28><15> ), .B(n1428), .Y(n1429) );
  OAI21X1 U1024 ( .A(n1238), .B(n1350), .C(n1429), .Y(n2343) );
  NAND3X1 U1025 ( .A(n1352), .B(n1354), .C(n1356), .Y(n1430) );
  NAND2X1 U1026 ( .A(\mem<27><0> ), .B(n1446), .Y(n1431) );
  OAI21X1 U1027 ( .A(n1239), .B(n1319), .C(n1431), .Y(n2342) );
  NAND2X1 U1028 ( .A(\mem<27><1> ), .B(n1446), .Y(n1432) );
  OAI21X1 U1029 ( .A(n1239), .B(n1322), .C(n1432), .Y(n2341) );
  NAND2X1 U1030 ( .A(\mem<27><2> ), .B(n1446), .Y(n1433) );
  OAI21X1 U1031 ( .A(n1239), .B(n1324), .C(n1433), .Y(n2340) );
  NAND2X1 U1032 ( .A(\mem<27><3> ), .B(n1446), .Y(n1434) );
  OAI21X1 U1033 ( .A(n1239), .B(n1326), .C(n1434), .Y(n2339) );
  NAND2X1 U1034 ( .A(\mem<27><4> ), .B(n1446), .Y(n1435) );
  OAI21X1 U1035 ( .A(n1239), .B(n1328), .C(n1435), .Y(n2338) );
  NAND2X1 U1036 ( .A(\mem<27><5> ), .B(n1446), .Y(n1436) );
  OAI21X1 U1037 ( .A(n1239), .B(n1330), .C(n1436), .Y(n2337) );
  NAND2X1 U1038 ( .A(\mem<27><6> ), .B(n1446), .Y(n1437) );
  OAI21X1 U1039 ( .A(n1239), .B(n1332), .C(n1437), .Y(n2336) );
  NAND2X1 U1040 ( .A(\mem<27><7> ), .B(n1446), .Y(n1438) );
  OAI21X1 U1041 ( .A(n1239), .B(n1334), .C(n1438), .Y(n2335) );
  NAND2X1 U1042 ( .A(\mem<27><8> ), .B(n1446), .Y(n1439) );
  OAI21X1 U1043 ( .A(n1240), .B(n1336), .C(n1439), .Y(n2334) );
  NAND2X1 U1044 ( .A(\mem<27><9> ), .B(n1446), .Y(n1440) );
  OAI21X1 U1045 ( .A(n1240), .B(n1338), .C(n1440), .Y(n2333) );
  NAND2X1 U1046 ( .A(\mem<27><10> ), .B(n1446), .Y(n1441) );
  OAI21X1 U1047 ( .A(n1240), .B(n1340), .C(n1441), .Y(n2332) );
  NAND2X1 U1048 ( .A(\mem<27><11> ), .B(n1446), .Y(n1442) );
  OAI21X1 U1049 ( .A(n1240), .B(n1342), .C(n1442), .Y(n2331) );
  NAND2X1 U1050 ( .A(\mem<27><12> ), .B(n1446), .Y(n1443) );
  OAI21X1 U1051 ( .A(n1240), .B(n1344), .C(n1443), .Y(n2330) );
  NAND2X1 U1052 ( .A(\mem<27><13> ), .B(n1446), .Y(n1444) );
  OAI21X1 U1053 ( .A(n1240), .B(n1346), .C(n1444), .Y(n2329) );
  NAND2X1 U1054 ( .A(\mem<27><14> ), .B(n1446), .Y(n1445) );
  OAI21X1 U1055 ( .A(n1240), .B(n1348), .C(n1445), .Y(n2328) );
  NAND2X1 U1056 ( .A(\mem<27><15> ), .B(n1446), .Y(n1447) );
  OAI21X1 U1057 ( .A(n1240), .B(n1350), .C(n1447), .Y(n2327) );
  NAND3X1 U1058 ( .A(n1356), .B(n1354), .C(n1353), .Y(n1448) );
  NAND2X1 U1059 ( .A(\mem<26><0> ), .B(n1464), .Y(n1449) );
  OAI21X1 U1060 ( .A(n1241), .B(n1319), .C(n1449), .Y(n2326) );
  NAND2X1 U1061 ( .A(\mem<26><1> ), .B(n1464), .Y(n1450) );
  OAI21X1 U1062 ( .A(n1241), .B(n1322), .C(n1450), .Y(n2325) );
  NAND2X1 U1063 ( .A(\mem<26><2> ), .B(n1464), .Y(n1451) );
  OAI21X1 U1064 ( .A(n1241), .B(n1324), .C(n1451), .Y(n2324) );
  NAND2X1 U1065 ( .A(\mem<26><3> ), .B(n1464), .Y(n1452) );
  OAI21X1 U1066 ( .A(n1241), .B(n1326), .C(n1452), .Y(n2323) );
  NAND2X1 U1067 ( .A(\mem<26><4> ), .B(n1464), .Y(n1453) );
  OAI21X1 U1068 ( .A(n1241), .B(n1328), .C(n1453), .Y(n2322) );
  NAND2X1 U1069 ( .A(\mem<26><5> ), .B(n1464), .Y(n1454) );
  OAI21X1 U1070 ( .A(n1241), .B(n1330), .C(n1454), .Y(n2321) );
  NAND2X1 U1071 ( .A(\mem<26><6> ), .B(n1464), .Y(n1455) );
  OAI21X1 U1072 ( .A(n1241), .B(n1332), .C(n1455), .Y(n2320) );
  NAND2X1 U1073 ( .A(\mem<26><7> ), .B(n1464), .Y(n1456) );
  OAI21X1 U1074 ( .A(n1241), .B(n1334), .C(n1456), .Y(n2319) );
  NAND2X1 U1075 ( .A(\mem<26><8> ), .B(n1464), .Y(n1457) );
  OAI21X1 U1076 ( .A(n1242), .B(n1336), .C(n1457), .Y(n2318) );
  NAND2X1 U1077 ( .A(\mem<26><9> ), .B(n1464), .Y(n1458) );
  OAI21X1 U1078 ( .A(n1242), .B(n1338), .C(n1458), .Y(n2317) );
  NAND2X1 U1079 ( .A(\mem<26><10> ), .B(n1464), .Y(n1459) );
  OAI21X1 U1080 ( .A(n1242), .B(n1340), .C(n1459), .Y(n2316) );
  NAND2X1 U1081 ( .A(\mem<26><11> ), .B(n1464), .Y(n1460) );
  OAI21X1 U1082 ( .A(n1242), .B(n1342), .C(n1460), .Y(n2315) );
  NAND2X1 U1083 ( .A(\mem<26><12> ), .B(n1464), .Y(n1461) );
  OAI21X1 U1084 ( .A(n1242), .B(n1344), .C(n1461), .Y(n2314) );
  NAND2X1 U1085 ( .A(\mem<26><13> ), .B(n1464), .Y(n1462) );
  OAI21X1 U1086 ( .A(n1242), .B(n1346), .C(n1462), .Y(n2313) );
  NAND2X1 U1087 ( .A(\mem<26><14> ), .B(n1464), .Y(n1463) );
  OAI21X1 U1088 ( .A(n1242), .B(n1348), .C(n1463), .Y(n2312) );
  NAND2X1 U1089 ( .A(\mem<26><15> ), .B(n1464), .Y(n1465) );
  OAI21X1 U1090 ( .A(n1242), .B(n1350), .C(n1465), .Y(n2311) );
  NAND3X1 U1091 ( .A(n1352), .B(n1356), .C(n1355), .Y(n1466) );
  NAND2X1 U1092 ( .A(\mem<25><0> ), .B(n1482), .Y(n1467) );
  OAI21X1 U1093 ( .A(n1243), .B(n1319), .C(n1467), .Y(n2310) );
  NAND2X1 U1094 ( .A(\mem<25><1> ), .B(n1482), .Y(n1468) );
  OAI21X1 U1095 ( .A(n1243), .B(n1322), .C(n1468), .Y(n2309) );
  NAND2X1 U1096 ( .A(\mem<25><2> ), .B(n1482), .Y(n1469) );
  OAI21X1 U1097 ( .A(n1243), .B(n1324), .C(n1469), .Y(n2308) );
  NAND2X1 U1098 ( .A(\mem<25><3> ), .B(n1482), .Y(n1470) );
  OAI21X1 U1099 ( .A(n1243), .B(n1326), .C(n1470), .Y(n2307) );
  NAND2X1 U1100 ( .A(\mem<25><4> ), .B(n1482), .Y(n1471) );
  OAI21X1 U1101 ( .A(n1243), .B(n1328), .C(n1471), .Y(n2306) );
  NAND2X1 U1102 ( .A(\mem<25><5> ), .B(n1482), .Y(n1472) );
  OAI21X1 U1103 ( .A(n1243), .B(n1330), .C(n1472), .Y(n2305) );
  NAND2X1 U1104 ( .A(\mem<25><6> ), .B(n1482), .Y(n1473) );
  OAI21X1 U1105 ( .A(n1243), .B(n1332), .C(n1473), .Y(n2304) );
  NAND2X1 U1106 ( .A(\mem<25><7> ), .B(n1482), .Y(n1474) );
  OAI21X1 U1107 ( .A(n1243), .B(n1334), .C(n1474), .Y(n2303) );
  NAND2X1 U1108 ( .A(\mem<25><8> ), .B(n1482), .Y(n1475) );
  OAI21X1 U1109 ( .A(n1244), .B(n1336), .C(n1475), .Y(n2302) );
  NAND2X1 U1110 ( .A(\mem<25><9> ), .B(n1482), .Y(n1476) );
  OAI21X1 U1111 ( .A(n1244), .B(n1338), .C(n1476), .Y(n2301) );
  NAND2X1 U1112 ( .A(\mem<25><10> ), .B(n1482), .Y(n1477) );
  OAI21X1 U1113 ( .A(n1244), .B(n1340), .C(n1477), .Y(n2300) );
  NAND2X1 U1114 ( .A(\mem<25><11> ), .B(n1482), .Y(n1478) );
  OAI21X1 U1115 ( .A(n1244), .B(n1342), .C(n1478), .Y(n2299) );
  NAND2X1 U1116 ( .A(\mem<25><12> ), .B(n1482), .Y(n1479) );
  OAI21X1 U1117 ( .A(n1244), .B(n1344), .C(n1479), .Y(n2298) );
  NAND2X1 U1118 ( .A(\mem<25><13> ), .B(n1482), .Y(n1480) );
  OAI21X1 U1119 ( .A(n1244), .B(n1346), .C(n1480), .Y(n2297) );
  NAND2X1 U1120 ( .A(\mem<25><14> ), .B(n1482), .Y(n1481) );
  OAI21X1 U1121 ( .A(n1244), .B(n1348), .C(n1481), .Y(n2296) );
  NAND2X1 U1122 ( .A(\mem<25><15> ), .B(n1482), .Y(n1483) );
  OAI21X1 U1123 ( .A(n1244), .B(n1350), .C(n1483), .Y(n2295) );
  NOR3X1 U1124 ( .A(n1352), .B(n1354), .C(n1187), .Y(n1878) );
  NAND2X1 U1125 ( .A(\mem<24><0> ), .B(n1246), .Y(n1484) );
  OAI21X1 U1126 ( .A(n1245), .B(n1319), .C(n1484), .Y(n2294) );
  NAND2X1 U1127 ( .A(\mem<24><1> ), .B(n1246), .Y(n1485) );
  OAI21X1 U1128 ( .A(n1245), .B(n1322), .C(n1485), .Y(n2293) );
  NAND2X1 U1129 ( .A(\mem<24><2> ), .B(n1246), .Y(n1486) );
  OAI21X1 U1130 ( .A(n1245), .B(n1324), .C(n1486), .Y(n2292) );
  NAND2X1 U1131 ( .A(\mem<24><3> ), .B(n1246), .Y(n1487) );
  OAI21X1 U1132 ( .A(n1245), .B(n1326), .C(n1487), .Y(n2291) );
  NAND2X1 U1133 ( .A(\mem<24><4> ), .B(n1246), .Y(n1488) );
  OAI21X1 U1134 ( .A(n1245), .B(n1328), .C(n1488), .Y(n2290) );
  NAND2X1 U1135 ( .A(\mem<24><5> ), .B(n1246), .Y(n1489) );
  OAI21X1 U1136 ( .A(n1245), .B(n1330), .C(n1489), .Y(n2289) );
  NAND2X1 U1137 ( .A(\mem<24><6> ), .B(n1246), .Y(n1490) );
  OAI21X1 U1138 ( .A(n1245), .B(n1332), .C(n1490), .Y(n2288) );
  NAND2X1 U1139 ( .A(\mem<24><7> ), .B(n1246), .Y(n1491) );
  OAI21X1 U1140 ( .A(n1245), .B(n1334), .C(n1491), .Y(n2287) );
  NAND2X1 U1141 ( .A(\mem<24><8> ), .B(n1247), .Y(n1492) );
  OAI21X1 U1142 ( .A(n1245), .B(n1336), .C(n1492), .Y(n2286) );
  NAND2X1 U1143 ( .A(\mem<24><9> ), .B(n1247), .Y(n1493) );
  OAI21X1 U1144 ( .A(n1245), .B(n1338), .C(n1493), .Y(n2285) );
  NAND2X1 U1145 ( .A(\mem<24><10> ), .B(n1247), .Y(n1494) );
  OAI21X1 U1146 ( .A(n1245), .B(n1340), .C(n1494), .Y(n2284) );
  NAND2X1 U1147 ( .A(\mem<24><11> ), .B(n1247), .Y(n1495) );
  OAI21X1 U1148 ( .A(n1245), .B(n1342), .C(n1495), .Y(n2283) );
  NAND2X1 U1149 ( .A(\mem<24><12> ), .B(n1247), .Y(n1496) );
  OAI21X1 U1150 ( .A(n1245), .B(n1344), .C(n1496), .Y(n2282) );
  NAND2X1 U1151 ( .A(\mem<24><13> ), .B(n1247), .Y(n1497) );
  OAI21X1 U1152 ( .A(n1245), .B(n1346), .C(n1497), .Y(n2281) );
  NAND2X1 U1153 ( .A(\mem<24><14> ), .B(n1247), .Y(n1498) );
  OAI21X1 U1154 ( .A(n1245), .B(n1348), .C(n1498), .Y(n2280) );
  NAND2X1 U1155 ( .A(\mem<24><15> ), .B(n1247), .Y(n1499) );
  OAI21X1 U1156 ( .A(n1245), .B(n1350), .C(n1499), .Y(n2279) );
  NAND2X1 U1157 ( .A(\mem<23><0> ), .B(n1515), .Y(n1500) );
  OAI21X1 U1158 ( .A(n1248), .B(n1319), .C(n1500), .Y(n2278) );
  NAND2X1 U1159 ( .A(\mem<23><1> ), .B(n1515), .Y(n1501) );
  OAI21X1 U1160 ( .A(n1248), .B(n1322), .C(n1501), .Y(n2277) );
  NAND2X1 U1161 ( .A(\mem<23><2> ), .B(n1515), .Y(n1502) );
  OAI21X1 U1162 ( .A(n1248), .B(n1324), .C(n1502), .Y(n2276) );
  NAND2X1 U1163 ( .A(\mem<23><3> ), .B(n1515), .Y(n1503) );
  OAI21X1 U1164 ( .A(n1248), .B(n1326), .C(n1503), .Y(n2275) );
  NAND2X1 U1165 ( .A(\mem<23><4> ), .B(n1515), .Y(n1504) );
  OAI21X1 U1166 ( .A(n1248), .B(n1328), .C(n1504), .Y(n2274) );
  NAND2X1 U1167 ( .A(\mem<23><5> ), .B(n1515), .Y(n1505) );
  OAI21X1 U1168 ( .A(n1248), .B(n1330), .C(n1505), .Y(n2273) );
  NAND2X1 U1169 ( .A(\mem<23><6> ), .B(n1515), .Y(n1506) );
  OAI21X1 U1170 ( .A(n1248), .B(n1332), .C(n1506), .Y(n2272) );
  NAND2X1 U1171 ( .A(\mem<23><7> ), .B(n1515), .Y(n1507) );
  OAI21X1 U1172 ( .A(n1248), .B(n1334), .C(n1507), .Y(n2271) );
  NAND2X1 U1173 ( .A(\mem<23><8> ), .B(n1515), .Y(n1508) );
  OAI21X1 U1174 ( .A(n1249), .B(n1336), .C(n1508), .Y(n2270) );
  NAND2X1 U1175 ( .A(\mem<23><9> ), .B(n1515), .Y(n1509) );
  OAI21X1 U1177 ( .A(n1249), .B(n1338), .C(n1509), .Y(n2269) );
  NAND2X1 U1178 ( .A(\mem<23><10> ), .B(n1515), .Y(n1510) );
  OAI21X1 U1179 ( .A(n1249), .B(n1340), .C(n1510), .Y(n2268) );
  NAND2X1 U1180 ( .A(\mem<23><11> ), .B(n1515), .Y(n1511) );
  OAI21X1 U1181 ( .A(n1249), .B(n1342), .C(n1511), .Y(n2267) );
  NAND2X1 U1182 ( .A(\mem<23><12> ), .B(n1515), .Y(n1512) );
  OAI21X1 U1183 ( .A(n1249), .B(n1344), .C(n1512), .Y(n2266) );
  NAND2X1 U1184 ( .A(\mem<23><13> ), .B(n1515), .Y(n1513) );
  OAI21X1 U1185 ( .A(n1249), .B(n1346), .C(n1513), .Y(n2265) );
  NAND2X1 U1186 ( .A(\mem<23><14> ), .B(n1515), .Y(n1514) );
  OAI21X1 U1187 ( .A(n1249), .B(n1348), .C(n1514), .Y(n2264) );
  NAND2X1 U1188 ( .A(\mem<23><15> ), .B(n1515), .Y(n1516) );
  OAI21X1 U1189 ( .A(n1249), .B(n1350), .C(n1516), .Y(n2263) );
  NAND2X1 U1190 ( .A(\mem<22><0> ), .B(n1252), .Y(n1517) );
  OAI21X1 U1191 ( .A(n1250), .B(n1319), .C(n1517), .Y(n2262) );
  NAND2X1 U1192 ( .A(\mem<22><1> ), .B(n1252), .Y(n1518) );
  OAI21X1 U1193 ( .A(n1250), .B(n1322), .C(n1518), .Y(n2261) );
  NAND2X1 U1194 ( .A(\mem<22><2> ), .B(n1252), .Y(n1519) );
  OAI21X1 U1195 ( .A(n1250), .B(n1324), .C(n1519), .Y(n2260) );
  NAND2X1 U1196 ( .A(\mem<22><3> ), .B(n1252), .Y(n1520) );
  OAI21X1 U1197 ( .A(n1250), .B(n1326), .C(n1520), .Y(n2259) );
  NAND2X1 U1198 ( .A(\mem<22><4> ), .B(n1252), .Y(n1521) );
  OAI21X1 U1199 ( .A(n1250), .B(n1328), .C(n1521), .Y(n2258) );
  NAND2X1 U1200 ( .A(\mem<22><5> ), .B(n1252), .Y(n1522) );
  OAI21X1 U1201 ( .A(n1250), .B(n1330), .C(n1522), .Y(n2257) );
  NAND2X1 U1202 ( .A(\mem<22><6> ), .B(n1252), .Y(n1523) );
  OAI21X1 U1203 ( .A(n1250), .B(n1332), .C(n1523), .Y(n2256) );
  NAND2X1 U1204 ( .A(\mem<22><7> ), .B(n1252), .Y(n1524) );
  OAI21X1 U1205 ( .A(n1250), .B(n1334), .C(n1524), .Y(n2255) );
  NAND2X1 U1206 ( .A(\mem<22><8> ), .B(n1253), .Y(n1525) );
  OAI21X1 U1207 ( .A(n1251), .B(n1336), .C(n1525), .Y(n2254) );
  NAND2X1 U1208 ( .A(\mem<22><9> ), .B(n1253), .Y(n1526) );
  OAI21X1 U1209 ( .A(n1251), .B(n1338), .C(n1526), .Y(n2253) );
  NAND2X1 U1210 ( .A(\mem<22><10> ), .B(n1253), .Y(n1527) );
  OAI21X1 U1211 ( .A(n1251), .B(n1340), .C(n1527), .Y(n2252) );
  NAND2X1 U1212 ( .A(\mem<22><11> ), .B(n1253), .Y(n1528) );
  OAI21X1 U1213 ( .A(n1251), .B(n1342), .C(n1528), .Y(n2251) );
  NAND2X1 U1214 ( .A(\mem<22><12> ), .B(n1253), .Y(n1529) );
  OAI21X1 U1215 ( .A(n1251), .B(n1344), .C(n1529), .Y(n2250) );
  NAND2X1 U1216 ( .A(\mem<22><13> ), .B(n1253), .Y(n1530) );
  OAI21X1 U1217 ( .A(n1251), .B(n1346), .C(n1530), .Y(n2249) );
  NAND2X1 U1218 ( .A(\mem<22><14> ), .B(n1253), .Y(n1531) );
  OAI21X1 U1219 ( .A(n1251), .B(n1348), .C(n1531), .Y(n2248) );
  NAND2X1 U1220 ( .A(\mem<22><15> ), .B(n1253), .Y(n1532) );
  OAI21X1 U1221 ( .A(n1251), .B(n1350), .C(n1532), .Y(n2247) );
  NAND2X1 U1222 ( .A(\mem<21><0> ), .B(n1256), .Y(n1533) );
  OAI21X1 U1223 ( .A(n1254), .B(n1319), .C(n1533), .Y(n2246) );
  NAND2X1 U1224 ( .A(\mem<21><1> ), .B(n1256), .Y(n1534) );
  OAI21X1 U1225 ( .A(n1254), .B(n1322), .C(n1534), .Y(n2245) );
  NAND2X1 U1226 ( .A(\mem<21><2> ), .B(n1256), .Y(n1535) );
  OAI21X1 U1227 ( .A(n1254), .B(n1324), .C(n1535), .Y(n2244) );
  NAND2X1 U1228 ( .A(\mem<21><3> ), .B(n1256), .Y(n1536) );
  OAI21X1 U1229 ( .A(n1254), .B(n1326), .C(n1536), .Y(n2243) );
  NAND2X1 U1230 ( .A(\mem<21><4> ), .B(n1256), .Y(n1537) );
  OAI21X1 U1231 ( .A(n1254), .B(n1328), .C(n1537), .Y(n2242) );
  NAND2X1 U1232 ( .A(\mem<21><5> ), .B(n1256), .Y(n1538) );
  OAI21X1 U1233 ( .A(n1254), .B(n1330), .C(n1538), .Y(n2241) );
  NAND2X1 U1234 ( .A(\mem<21><6> ), .B(n1256), .Y(n1539) );
  OAI21X1 U1235 ( .A(n1254), .B(n1332), .C(n1539), .Y(n2240) );
  NAND2X1 U1236 ( .A(\mem<21><7> ), .B(n1256), .Y(n1540) );
  OAI21X1 U1237 ( .A(n1254), .B(n1334), .C(n1540), .Y(n2239) );
  NAND2X1 U1238 ( .A(\mem<21><8> ), .B(n1257), .Y(n1541) );
  OAI21X1 U1239 ( .A(n1255), .B(n1336), .C(n1541), .Y(n2238) );
  NAND2X1 U1240 ( .A(\mem<21><9> ), .B(n1257), .Y(n1542) );
  OAI21X1 U1241 ( .A(n1255), .B(n1338), .C(n1542), .Y(n2237) );
  NAND2X1 U1242 ( .A(\mem<21><10> ), .B(n1257), .Y(n1543) );
  OAI21X1 U1243 ( .A(n1255), .B(n1340), .C(n1543), .Y(n2236) );
  NAND2X1 U1244 ( .A(\mem<21><11> ), .B(n1257), .Y(n1544) );
  OAI21X1 U1245 ( .A(n1255), .B(n1342), .C(n1544), .Y(n2235) );
  NAND2X1 U1246 ( .A(\mem<21><12> ), .B(n1257), .Y(n1545) );
  OAI21X1 U1247 ( .A(n1255), .B(n1344), .C(n1545), .Y(n2234) );
  NAND2X1 U1248 ( .A(\mem<21><13> ), .B(n1257), .Y(n1546) );
  OAI21X1 U1249 ( .A(n1255), .B(n1346), .C(n1546), .Y(n2233) );
  NAND2X1 U1250 ( .A(\mem<21><14> ), .B(n1257), .Y(n1547) );
  OAI21X1 U1251 ( .A(n1255), .B(n1348), .C(n1547), .Y(n2232) );
  NAND2X1 U1252 ( .A(\mem<21><15> ), .B(n1257), .Y(n1548) );
  OAI21X1 U1253 ( .A(n1255), .B(n1350), .C(n1548), .Y(n2231) );
  NAND2X1 U1254 ( .A(\mem<20><0> ), .B(n1260), .Y(n1549) );
  OAI21X1 U1255 ( .A(n1258), .B(n1319), .C(n1549), .Y(n2230) );
  NAND2X1 U1256 ( .A(\mem<20><1> ), .B(n1260), .Y(n1550) );
  OAI21X1 U1257 ( .A(n1258), .B(n1322), .C(n1550), .Y(n2229) );
  NAND2X1 U1258 ( .A(\mem<20><2> ), .B(n1260), .Y(n1551) );
  OAI21X1 U1259 ( .A(n1258), .B(n1324), .C(n1551), .Y(n2228) );
  NAND2X1 U1260 ( .A(\mem<20><3> ), .B(n1260), .Y(n1552) );
  OAI21X1 U1261 ( .A(n1258), .B(n1326), .C(n1552), .Y(n2227) );
  NAND2X1 U1262 ( .A(\mem<20><4> ), .B(n1260), .Y(n1553) );
  OAI21X1 U1263 ( .A(n1258), .B(n1328), .C(n1553), .Y(n2226) );
  NAND2X1 U1264 ( .A(\mem<20><5> ), .B(n1260), .Y(n1554) );
  OAI21X1 U1265 ( .A(n1258), .B(n1330), .C(n1554), .Y(n2225) );
  NAND2X1 U1266 ( .A(\mem<20><6> ), .B(n1260), .Y(n1555) );
  OAI21X1 U1267 ( .A(n1258), .B(n1332), .C(n1555), .Y(n2224) );
  NAND2X1 U1268 ( .A(\mem<20><7> ), .B(n1260), .Y(n1556) );
  OAI21X1 U1269 ( .A(n1258), .B(n1334), .C(n1556), .Y(n2223) );
  NAND2X1 U1270 ( .A(\mem<20><8> ), .B(n1261), .Y(n1557) );
  OAI21X1 U1271 ( .A(n1259), .B(n1336), .C(n1557), .Y(n2222) );
  NAND2X1 U1272 ( .A(\mem<20><9> ), .B(n1261), .Y(n1558) );
  OAI21X1 U1273 ( .A(n1259), .B(n1338), .C(n1558), .Y(n2221) );
  NAND2X1 U1274 ( .A(\mem<20><10> ), .B(n1261), .Y(n1559) );
  OAI21X1 U1275 ( .A(n1259), .B(n1340), .C(n1559), .Y(n2220) );
  NAND2X1 U1276 ( .A(\mem<20><11> ), .B(n1261), .Y(n1560) );
  OAI21X1 U1277 ( .A(n1259), .B(n1342), .C(n1560), .Y(n2219) );
  NAND2X1 U1278 ( .A(\mem<20><12> ), .B(n1261), .Y(n1561) );
  OAI21X1 U1279 ( .A(n1259), .B(n1344), .C(n1561), .Y(n2218) );
  NAND2X1 U1280 ( .A(\mem<20><13> ), .B(n1261), .Y(n1562) );
  OAI21X1 U1281 ( .A(n1259), .B(n1346), .C(n1562), .Y(n2217) );
  NAND2X1 U1282 ( .A(\mem<20><14> ), .B(n1261), .Y(n1563) );
  OAI21X1 U1283 ( .A(n1259), .B(n1348), .C(n1563), .Y(n2216) );
  NAND2X1 U1284 ( .A(\mem<20><15> ), .B(n1261), .Y(n1564) );
  OAI21X1 U1285 ( .A(n1259), .B(n1350), .C(n1564), .Y(n2215) );
  NAND2X1 U1286 ( .A(\mem<19><0> ), .B(n125), .Y(n1565) );
  OAI21X1 U1287 ( .A(n1262), .B(n1319), .C(n1565), .Y(n2214) );
  NAND2X1 U1288 ( .A(\mem<19><1> ), .B(n125), .Y(n1566) );
  OAI21X1 U1289 ( .A(n1262), .B(n1321), .C(n1566), .Y(n2213) );
  NAND2X1 U1290 ( .A(\mem<19><2> ), .B(n125), .Y(n1567) );
  OAI21X1 U1291 ( .A(n1262), .B(n1323), .C(n1567), .Y(n2212) );
  NAND2X1 U1292 ( .A(\mem<19><3> ), .B(n125), .Y(n1568) );
  OAI21X1 U1293 ( .A(n1262), .B(n1325), .C(n1568), .Y(n2211) );
  NAND2X1 U1294 ( .A(\mem<19><4> ), .B(n125), .Y(n1569) );
  OAI21X1 U1295 ( .A(n1262), .B(n1327), .C(n1569), .Y(n2210) );
  NAND2X1 U1296 ( .A(\mem<19><5> ), .B(n125), .Y(n1570) );
  OAI21X1 U1297 ( .A(n1262), .B(n1329), .C(n1570), .Y(n2209) );
  NAND2X1 U1298 ( .A(\mem<19><6> ), .B(n125), .Y(n1571) );
  OAI21X1 U1299 ( .A(n1262), .B(n1331), .C(n1571), .Y(n2208) );
  NAND2X1 U1300 ( .A(\mem<19><7> ), .B(n125), .Y(n1572) );
  OAI21X1 U1301 ( .A(n1262), .B(n1333), .C(n1572), .Y(n2207) );
  NAND2X1 U1302 ( .A(\mem<19><8> ), .B(n125), .Y(n1573) );
  OAI21X1 U1303 ( .A(n1263), .B(n1336), .C(n1573), .Y(n2206) );
  NAND2X1 U1304 ( .A(\mem<19><9> ), .B(n125), .Y(n1574) );
  OAI21X1 U1305 ( .A(n1263), .B(n1338), .C(n1574), .Y(n2205) );
  NAND2X1 U1306 ( .A(\mem<19><10> ), .B(n125), .Y(n1575) );
  OAI21X1 U1307 ( .A(n1263), .B(n1340), .C(n1575), .Y(n2204) );
  NAND2X1 U1308 ( .A(\mem<19><11> ), .B(n125), .Y(n1576) );
  OAI21X1 U1309 ( .A(n1263), .B(n1342), .C(n1576), .Y(n2203) );
  NAND2X1 U1310 ( .A(\mem<19><12> ), .B(n125), .Y(n1577) );
  OAI21X1 U1311 ( .A(n1263), .B(n1344), .C(n1577), .Y(n2202) );
  NAND2X1 U1312 ( .A(\mem<19><13> ), .B(n125), .Y(n1578) );
  OAI21X1 U1313 ( .A(n1263), .B(n1346), .C(n1578), .Y(n2201) );
  NAND2X1 U1314 ( .A(\mem<19><14> ), .B(n125), .Y(n1579) );
  OAI21X1 U1315 ( .A(n1263), .B(n1348), .C(n1579), .Y(n2200) );
  NAND2X1 U1316 ( .A(\mem<19><15> ), .B(n125), .Y(n1580) );
  OAI21X1 U1317 ( .A(n1263), .B(n1350), .C(n1580), .Y(n2199) );
  NAND2X1 U1318 ( .A(\mem<18><0> ), .B(n128), .Y(n1581) );
  OAI21X1 U1319 ( .A(n1264), .B(n1320), .C(n1581), .Y(n2198) );
  NAND2X1 U1320 ( .A(\mem<18><1> ), .B(n128), .Y(n1582) );
  OAI21X1 U1321 ( .A(n1264), .B(n1322), .C(n1582), .Y(n2197) );
  NAND2X1 U1322 ( .A(\mem<18><2> ), .B(n128), .Y(n1583) );
  OAI21X1 U1323 ( .A(n1264), .B(n1324), .C(n1583), .Y(n2196) );
  NAND2X1 U1324 ( .A(\mem<18><3> ), .B(n128), .Y(n1584) );
  OAI21X1 U1325 ( .A(n1264), .B(n1326), .C(n1584), .Y(n2195) );
  NAND2X1 U1326 ( .A(\mem<18><4> ), .B(n128), .Y(n1585) );
  OAI21X1 U1327 ( .A(n1264), .B(n1328), .C(n1585), .Y(n2194) );
  NAND2X1 U1328 ( .A(\mem<18><5> ), .B(n128), .Y(n1586) );
  OAI21X1 U1329 ( .A(n1264), .B(n1330), .C(n1586), .Y(n2193) );
  NAND2X1 U1330 ( .A(\mem<18><6> ), .B(n128), .Y(n1587) );
  OAI21X1 U1331 ( .A(n1264), .B(n1332), .C(n1587), .Y(n2192) );
  NAND2X1 U1332 ( .A(\mem<18><7> ), .B(n128), .Y(n1588) );
  OAI21X1 U1333 ( .A(n1264), .B(n1334), .C(n1588), .Y(n2191) );
  NAND2X1 U1334 ( .A(\mem<18><8> ), .B(n128), .Y(n1589) );
  OAI21X1 U1335 ( .A(n1265), .B(n1335), .C(n1589), .Y(n2190) );
  NAND2X1 U1336 ( .A(\mem<18><9> ), .B(n128), .Y(n1590) );
  OAI21X1 U1337 ( .A(n1265), .B(n1337), .C(n1590), .Y(n2189) );
  NAND2X1 U1338 ( .A(\mem<18><10> ), .B(n128), .Y(n1591) );
  OAI21X1 U1339 ( .A(n1265), .B(n1339), .C(n1591), .Y(n2188) );
  NAND2X1 U1340 ( .A(\mem<18><11> ), .B(n128), .Y(n1592) );
  OAI21X1 U1341 ( .A(n1265), .B(n1341), .C(n1592), .Y(n2187) );
  NAND2X1 U1342 ( .A(\mem<18><12> ), .B(n128), .Y(n1593) );
  OAI21X1 U1343 ( .A(n1265), .B(n1343), .C(n1593), .Y(n2186) );
  NAND2X1 U1344 ( .A(\mem<18><13> ), .B(n128), .Y(n1594) );
  OAI21X1 U1345 ( .A(n1265), .B(n1345), .C(n1594), .Y(n2185) );
  NAND2X1 U1346 ( .A(\mem<18><14> ), .B(n128), .Y(n1595) );
  OAI21X1 U1347 ( .A(n1265), .B(n1347), .C(n1595), .Y(n2184) );
  NAND2X1 U1348 ( .A(\mem<18><15> ), .B(n128), .Y(n1596) );
  OAI21X1 U1349 ( .A(n1265), .B(n1349), .C(n1596), .Y(n2183) );
  NAND2X1 U1350 ( .A(\mem<17><0> ), .B(n1268), .Y(n1597) );
  OAI21X1 U1351 ( .A(n1266), .B(n1319), .C(n1597), .Y(n2182) );
  NAND2X1 U1352 ( .A(\mem<17><1> ), .B(n1268), .Y(n1598) );
  OAI21X1 U1353 ( .A(n1266), .B(n1321), .C(n1598), .Y(n2181) );
  NAND2X1 U1354 ( .A(\mem<17><2> ), .B(n1268), .Y(n1599) );
  OAI21X1 U1355 ( .A(n1266), .B(n1323), .C(n1599), .Y(n2180) );
  NAND2X1 U1356 ( .A(\mem<17><3> ), .B(n1268), .Y(n1600) );
  OAI21X1 U1357 ( .A(n1266), .B(n1325), .C(n1600), .Y(n2179) );
  NAND2X1 U1358 ( .A(\mem<17><4> ), .B(n1268), .Y(n1601) );
  OAI21X1 U1359 ( .A(n1266), .B(n1327), .C(n1601), .Y(n2178) );
  NAND2X1 U1360 ( .A(\mem<17><5> ), .B(n1268), .Y(n1602) );
  OAI21X1 U1361 ( .A(n1266), .B(n1329), .C(n1602), .Y(n2177) );
  NAND2X1 U1362 ( .A(\mem<17><6> ), .B(n1268), .Y(n1603) );
  OAI21X1 U1363 ( .A(n1266), .B(n1331), .C(n1603), .Y(n2176) );
  NAND2X1 U1364 ( .A(\mem<17><7> ), .B(n1268), .Y(n1604) );
  OAI21X1 U1365 ( .A(n1266), .B(n1333), .C(n1604), .Y(n2175) );
  NAND2X1 U1366 ( .A(\mem<17><8> ), .B(n1269), .Y(n1605) );
  OAI21X1 U1367 ( .A(n1267), .B(n1336), .C(n1605), .Y(n2174) );
  NAND2X1 U1368 ( .A(\mem<17><9> ), .B(n1269), .Y(n1606) );
  OAI21X1 U1369 ( .A(n1267), .B(n1338), .C(n1606), .Y(n2173) );
  NAND2X1 U1370 ( .A(\mem<17><10> ), .B(n1269), .Y(n1607) );
  OAI21X1 U1371 ( .A(n1267), .B(n1340), .C(n1607), .Y(n2172) );
  NAND2X1 U1372 ( .A(\mem<17><11> ), .B(n1269), .Y(n1608) );
  OAI21X1 U1373 ( .A(n1267), .B(n1342), .C(n1608), .Y(n2171) );
  NAND2X1 U1374 ( .A(\mem<17><12> ), .B(n1269), .Y(n1609) );
  OAI21X1 U1375 ( .A(n1267), .B(n1344), .C(n1609), .Y(n2170) );
  NAND2X1 U1376 ( .A(\mem<17><13> ), .B(n1269), .Y(n1610) );
  OAI21X1 U1377 ( .A(n1267), .B(n1346), .C(n1610), .Y(n2169) );
  NAND2X1 U1378 ( .A(\mem<17><14> ), .B(n1269), .Y(n1611) );
  OAI21X1 U1379 ( .A(n1267), .B(n1348), .C(n1611), .Y(n2168) );
  NAND2X1 U1380 ( .A(\mem<17><15> ), .B(n1269), .Y(n1612) );
  OAI21X1 U1381 ( .A(n1267), .B(n1350), .C(n1612), .Y(n2167) );
  NAND2X1 U1382 ( .A(\mem<16><0> ), .B(n131), .Y(n1613) );
  OAI21X1 U1383 ( .A(n1270), .B(n1320), .C(n1613), .Y(n2166) );
  NAND2X1 U1384 ( .A(\mem<16><1> ), .B(n131), .Y(n1614) );
  OAI21X1 U1385 ( .A(n1270), .B(n1322), .C(n1614), .Y(n2165) );
  NAND2X1 U1386 ( .A(\mem<16><2> ), .B(n131), .Y(n1615) );
  OAI21X1 U1387 ( .A(n1270), .B(n1324), .C(n1615), .Y(n2164) );
  NAND2X1 U1388 ( .A(\mem<16><3> ), .B(n131), .Y(n1616) );
  OAI21X1 U1389 ( .A(n1270), .B(n1326), .C(n1616), .Y(n2163) );
  NAND2X1 U1390 ( .A(\mem<16><4> ), .B(n131), .Y(n1617) );
  OAI21X1 U1391 ( .A(n1270), .B(n1328), .C(n1617), .Y(n2162) );
  NAND2X1 U1392 ( .A(\mem<16><5> ), .B(n131), .Y(n1618) );
  OAI21X1 U1393 ( .A(n1270), .B(n1330), .C(n1618), .Y(n2161) );
  NAND2X1 U1394 ( .A(\mem<16><6> ), .B(n131), .Y(n1619) );
  OAI21X1 U1395 ( .A(n1270), .B(n1332), .C(n1619), .Y(n2160) );
  NAND2X1 U1396 ( .A(\mem<16><7> ), .B(n131), .Y(n1620) );
  OAI21X1 U1397 ( .A(n1270), .B(n1334), .C(n1620), .Y(n2159) );
  NAND2X1 U1398 ( .A(\mem<16><8> ), .B(n131), .Y(n1621) );
  OAI21X1 U1399 ( .A(n1270), .B(n1335), .C(n1621), .Y(n2158) );
  NAND2X1 U1400 ( .A(\mem<16><9> ), .B(n131), .Y(n1622) );
  OAI21X1 U1401 ( .A(n1270), .B(n1337), .C(n1622), .Y(n2157) );
  NAND2X1 U1402 ( .A(\mem<16><10> ), .B(n131), .Y(n1623) );
  OAI21X1 U1403 ( .A(n1270), .B(n1339), .C(n1623), .Y(n2156) );
  NAND2X1 U1404 ( .A(\mem<16><11> ), .B(n131), .Y(n1624) );
  OAI21X1 U1405 ( .A(n1270), .B(n1341), .C(n1624), .Y(n2155) );
  NAND2X1 U1406 ( .A(\mem<16><12> ), .B(n131), .Y(n1625) );
  OAI21X1 U1407 ( .A(n1270), .B(n1343), .C(n1625), .Y(n2154) );
  NAND2X1 U1408 ( .A(\mem<16><13> ), .B(n131), .Y(n1626) );
  OAI21X1 U1409 ( .A(n1270), .B(n1345), .C(n1626), .Y(n2153) );
  NAND2X1 U1410 ( .A(\mem<16><14> ), .B(n131), .Y(n1627) );
  OAI21X1 U1411 ( .A(n1270), .B(n1347), .C(n1627), .Y(n2152) );
  NAND2X1 U1412 ( .A(\mem<16><15> ), .B(n131), .Y(n1628) );
  OAI21X1 U1413 ( .A(n1270), .B(n1349), .C(n1628), .Y(n2151) );
  NAND3X1 U1414 ( .A(n1357), .B(n2407), .C(n1359), .Y(n1629) );
  NAND2X1 U1415 ( .A(\mem<15><0> ), .B(n1273), .Y(n1630) );
  OAI21X1 U1416 ( .A(n1271), .B(n1320), .C(n1630), .Y(n2150) );
  NAND2X1 U1417 ( .A(\mem<15><1> ), .B(n1273), .Y(n1631) );
  OAI21X1 U1418 ( .A(n1271), .B(n1322), .C(n1631), .Y(n2149) );
  NAND2X1 U1419 ( .A(\mem<15><2> ), .B(n1273), .Y(n1632) );
  OAI21X1 U1420 ( .A(n1271), .B(n1324), .C(n1632), .Y(n2148) );
  NAND2X1 U1421 ( .A(\mem<15><3> ), .B(n1273), .Y(n1633) );
  OAI21X1 U1422 ( .A(n1271), .B(n1326), .C(n1633), .Y(n2147) );
  NAND2X1 U1423 ( .A(\mem<15><4> ), .B(n1273), .Y(n1634) );
  OAI21X1 U1424 ( .A(n1271), .B(n1328), .C(n1634), .Y(n2146) );
  NAND2X1 U1425 ( .A(\mem<15><5> ), .B(n1273), .Y(n1635) );
  OAI21X1 U1426 ( .A(n1271), .B(n1330), .C(n1635), .Y(n2145) );
  NAND2X1 U1427 ( .A(\mem<15><6> ), .B(n1273), .Y(n1636) );
  OAI21X1 U1428 ( .A(n1271), .B(n1332), .C(n1636), .Y(n2144) );
  NAND2X1 U1429 ( .A(\mem<15><7> ), .B(n1273), .Y(n1637) );
  OAI21X1 U1430 ( .A(n1271), .B(n1334), .C(n1637), .Y(n2143) );
  NAND2X1 U1431 ( .A(\mem<15><8> ), .B(n1274), .Y(n1638) );
  OAI21X1 U1432 ( .A(n1272), .B(n1335), .C(n1638), .Y(n2142) );
  NAND2X1 U1433 ( .A(\mem<15><9> ), .B(n1274), .Y(n1639) );
  OAI21X1 U1434 ( .A(n1272), .B(n1337), .C(n1639), .Y(n2141) );
  NAND2X1 U1435 ( .A(\mem<15><10> ), .B(n1274), .Y(n1640) );
  OAI21X1 U1436 ( .A(n1272), .B(n1339), .C(n1640), .Y(n2140) );
  NAND2X1 U1437 ( .A(\mem<15><11> ), .B(n1274), .Y(n1641) );
  OAI21X1 U1438 ( .A(n1272), .B(n1341), .C(n1641), .Y(n2139) );
  NAND2X1 U1439 ( .A(\mem<15><12> ), .B(n1274), .Y(n1642) );
  OAI21X1 U1440 ( .A(n1272), .B(n1343), .C(n1642), .Y(n2138) );
  NAND2X1 U1441 ( .A(\mem<15><13> ), .B(n1274), .Y(n1643) );
  OAI21X1 U1442 ( .A(n1272), .B(n1345), .C(n1643), .Y(n2137) );
  NAND2X1 U1443 ( .A(\mem<15><14> ), .B(n1274), .Y(n1644) );
  OAI21X1 U1444 ( .A(n1272), .B(n1347), .C(n1644), .Y(n2136) );
  NAND2X1 U1445 ( .A(\mem<15><15> ), .B(n1274), .Y(n1645) );
  OAI21X1 U1446 ( .A(n1272), .B(n1349), .C(n1645), .Y(n2135) );
  NAND2X1 U1447 ( .A(\mem<14><0> ), .B(n1277), .Y(n1646) );
  OAI21X1 U1448 ( .A(n1275), .B(n1319), .C(n1646), .Y(n2134) );
  NAND2X1 U1449 ( .A(\mem<14><1> ), .B(n1277), .Y(n1647) );
  OAI21X1 U1450 ( .A(n1275), .B(n1321), .C(n1647), .Y(n2133) );
  NAND2X1 U1451 ( .A(\mem<14><2> ), .B(n1277), .Y(n1648) );
  OAI21X1 U1452 ( .A(n1275), .B(n1323), .C(n1648), .Y(n2132) );
  NAND2X1 U1453 ( .A(\mem<14><3> ), .B(n1277), .Y(n1649) );
  OAI21X1 U1454 ( .A(n1275), .B(n1325), .C(n1649), .Y(n2131) );
  NAND2X1 U1455 ( .A(\mem<14><4> ), .B(n1277), .Y(n1650) );
  OAI21X1 U1456 ( .A(n1275), .B(n1327), .C(n1650), .Y(n2130) );
  NAND2X1 U1457 ( .A(\mem<14><5> ), .B(n1277), .Y(n1651) );
  OAI21X1 U1458 ( .A(n1275), .B(n1329), .C(n1651), .Y(n2129) );
  NAND2X1 U1459 ( .A(\mem<14><6> ), .B(n1277), .Y(n1652) );
  OAI21X1 U1460 ( .A(n1275), .B(n1331), .C(n1652), .Y(n2128) );
  NAND2X1 U1461 ( .A(\mem<14><7> ), .B(n1277), .Y(n1653) );
  OAI21X1 U1462 ( .A(n1275), .B(n1333), .C(n1653), .Y(n2127) );
  NAND2X1 U1463 ( .A(\mem<14><8> ), .B(n1278), .Y(n1654) );
  OAI21X1 U1464 ( .A(n1276), .B(n1336), .C(n1654), .Y(n2126) );
  NAND2X1 U1465 ( .A(\mem<14><9> ), .B(n1278), .Y(n1655) );
  OAI21X1 U1466 ( .A(n1276), .B(n1338), .C(n1655), .Y(n2125) );
  NAND2X1 U1467 ( .A(\mem<14><10> ), .B(n1278), .Y(n1656) );
  OAI21X1 U1468 ( .A(n1276), .B(n1340), .C(n1656), .Y(n2124) );
  NAND2X1 U1469 ( .A(\mem<14><11> ), .B(n1278), .Y(n1657) );
  OAI21X1 U1470 ( .A(n1276), .B(n1342), .C(n1657), .Y(n2123) );
  NAND2X1 U1471 ( .A(\mem<14><12> ), .B(n1278), .Y(n1658) );
  OAI21X1 U1472 ( .A(n1276), .B(n1344), .C(n1658), .Y(n2122) );
  NAND2X1 U1473 ( .A(\mem<14><13> ), .B(n1278), .Y(n1659) );
  OAI21X1 U1474 ( .A(n1276), .B(n1346), .C(n1659), .Y(n2121) );
  NAND2X1 U1475 ( .A(\mem<14><14> ), .B(n1278), .Y(n1660) );
  OAI21X1 U1476 ( .A(n1276), .B(n1348), .C(n1660), .Y(n2120) );
  NAND2X1 U1477 ( .A(\mem<14><15> ), .B(n1278), .Y(n1661) );
  OAI21X1 U1478 ( .A(n1276), .B(n1350), .C(n1661), .Y(n2119) );
  NAND2X1 U1479 ( .A(\mem<13><0> ), .B(n1281), .Y(n1662) );
  OAI21X1 U1480 ( .A(n1279), .B(n1320), .C(n1662), .Y(n2118) );
  NAND2X1 U1481 ( .A(\mem<13><1> ), .B(n1281), .Y(n1663) );
  OAI21X1 U1482 ( .A(n1279), .B(n1322), .C(n1663), .Y(n2117) );
  NAND2X1 U1483 ( .A(\mem<13><2> ), .B(n1281), .Y(n1664) );
  OAI21X1 U1484 ( .A(n1279), .B(n1324), .C(n1664), .Y(n2116) );
  NAND2X1 U1485 ( .A(\mem<13><3> ), .B(n1281), .Y(n1665) );
  OAI21X1 U1486 ( .A(n1279), .B(n1326), .C(n1665), .Y(n2115) );
  NAND2X1 U1487 ( .A(\mem<13><4> ), .B(n1281), .Y(n1666) );
  OAI21X1 U1488 ( .A(n1279), .B(n1328), .C(n1666), .Y(n2114) );
  NAND2X1 U1489 ( .A(\mem<13><5> ), .B(n1281), .Y(n1667) );
  OAI21X1 U1490 ( .A(n1279), .B(n1330), .C(n1667), .Y(n2113) );
  NAND2X1 U1491 ( .A(\mem<13><6> ), .B(n1281), .Y(n1668) );
  OAI21X1 U1492 ( .A(n1279), .B(n1332), .C(n1668), .Y(n2112) );
  NAND2X1 U1493 ( .A(\mem<13><7> ), .B(n1281), .Y(n1669) );
  OAI21X1 U1494 ( .A(n1279), .B(n1334), .C(n1669), .Y(n2111) );
  NAND2X1 U1495 ( .A(\mem<13><8> ), .B(n1282), .Y(n1670) );
  OAI21X1 U1496 ( .A(n1280), .B(n1335), .C(n1670), .Y(n2110) );
  NAND2X1 U1497 ( .A(\mem<13><9> ), .B(n1282), .Y(n1671) );
  OAI21X1 U1498 ( .A(n1280), .B(n1337), .C(n1671), .Y(n2109) );
  NAND2X1 U1499 ( .A(\mem<13><10> ), .B(n1282), .Y(n1672) );
  OAI21X1 U1500 ( .A(n1280), .B(n1339), .C(n1672), .Y(n2108) );
  NAND2X1 U1501 ( .A(\mem<13><11> ), .B(n1282), .Y(n1673) );
  OAI21X1 U1502 ( .A(n1280), .B(n1341), .C(n1673), .Y(n2107) );
  NAND2X1 U1503 ( .A(\mem<13><12> ), .B(n1282), .Y(n1674) );
  OAI21X1 U1504 ( .A(n1280), .B(n1343), .C(n1674), .Y(n2106) );
  NAND2X1 U1505 ( .A(\mem<13><13> ), .B(n1282), .Y(n1675) );
  OAI21X1 U1506 ( .A(n1280), .B(n1345), .C(n1675), .Y(n2105) );
  NAND2X1 U1507 ( .A(\mem<13><14> ), .B(n1282), .Y(n1676) );
  OAI21X1 U1508 ( .A(n1280), .B(n1347), .C(n1676), .Y(n2104) );
  NAND2X1 U1509 ( .A(\mem<13><15> ), .B(n1282), .Y(n1677) );
  OAI21X1 U1510 ( .A(n1280), .B(n1349), .C(n1677), .Y(n2103) );
  NAND2X1 U1511 ( .A(\mem<12><0> ), .B(n1285), .Y(n1678) );
  OAI21X1 U1512 ( .A(n1283), .B(n1319), .C(n1678), .Y(n2102) );
  NAND2X1 U1513 ( .A(\mem<12><1> ), .B(n1285), .Y(n1679) );
  OAI21X1 U1514 ( .A(n1283), .B(n1321), .C(n1679), .Y(n2101) );
  NAND2X1 U1515 ( .A(\mem<12><2> ), .B(n1285), .Y(n1680) );
  OAI21X1 U1516 ( .A(n1283), .B(n1323), .C(n1680), .Y(n2100) );
  NAND2X1 U1517 ( .A(\mem<12><3> ), .B(n1285), .Y(n1681) );
  OAI21X1 U1518 ( .A(n1283), .B(n1325), .C(n1681), .Y(n2099) );
  NAND2X1 U1519 ( .A(\mem<12><4> ), .B(n1285), .Y(n1682) );
  OAI21X1 U1520 ( .A(n1283), .B(n1327), .C(n1682), .Y(n2098) );
  NAND2X1 U1521 ( .A(\mem<12><5> ), .B(n1285), .Y(n1683) );
  OAI21X1 U1522 ( .A(n1283), .B(n1329), .C(n1683), .Y(n2097) );
  NAND2X1 U1523 ( .A(\mem<12><6> ), .B(n1285), .Y(n1684) );
  OAI21X1 U1524 ( .A(n1283), .B(n1331), .C(n1684), .Y(n2096) );
  NAND2X1 U1525 ( .A(\mem<12><7> ), .B(n1285), .Y(n1685) );
  OAI21X1 U1526 ( .A(n1283), .B(n1333), .C(n1685), .Y(n2095) );
  NAND2X1 U1527 ( .A(\mem<12><8> ), .B(n1286), .Y(n1686) );
  OAI21X1 U1528 ( .A(n1284), .B(n1336), .C(n1686), .Y(n2094) );
  NAND2X1 U1529 ( .A(\mem<12><9> ), .B(n1286), .Y(n1687) );
  OAI21X1 U1530 ( .A(n1284), .B(n1338), .C(n1687), .Y(n2093) );
  NAND2X1 U1531 ( .A(\mem<12><10> ), .B(n1286), .Y(n1688) );
  OAI21X1 U1532 ( .A(n1284), .B(n1340), .C(n1688), .Y(n2092) );
  NAND2X1 U1533 ( .A(\mem<12><11> ), .B(n1286), .Y(n1689) );
  OAI21X1 U1534 ( .A(n1284), .B(n1342), .C(n1689), .Y(n2091) );
  NAND2X1 U1535 ( .A(\mem<12><12> ), .B(n1286), .Y(n1690) );
  OAI21X1 U1536 ( .A(n1284), .B(n1344), .C(n1690), .Y(n2090) );
  NAND2X1 U1537 ( .A(\mem<12><13> ), .B(n1286), .Y(n1691) );
  OAI21X1 U1538 ( .A(n1284), .B(n1346), .C(n1691), .Y(n2089) );
  NAND2X1 U1539 ( .A(\mem<12><14> ), .B(n1286), .Y(n1692) );
  OAI21X1 U1540 ( .A(n1284), .B(n1348), .C(n1692), .Y(n2088) );
  NAND2X1 U1541 ( .A(\mem<12><15> ), .B(n1286), .Y(n1693) );
  OAI21X1 U1542 ( .A(n1284), .B(n1350), .C(n1693), .Y(n2087) );
  NAND2X1 U1543 ( .A(\mem<11><0> ), .B(n1289), .Y(n1694) );
  OAI21X1 U1544 ( .A(n1287), .B(n1320), .C(n1694), .Y(n2086) );
  NAND2X1 U1545 ( .A(\mem<11><1> ), .B(n1289), .Y(n1695) );
  OAI21X1 U1546 ( .A(n1287), .B(n1321), .C(n1695), .Y(n2085) );
  NAND2X1 U1547 ( .A(\mem<11><2> ), .B(n1289), .Y(n1696) );
  OAI21X1 U1548 ( .A(n1287), .B(n1323), .C(n1696), .Y(n2084) );
  NAND2X1 U1549 ( .A(\mem<11><3> ), .B(n1289), .Y(n1697) );
  OAI21X1 U1550 ( .A(n1287), .B(n1325), .C(n1697), .Y(n2083) );
  NAND2X1 U1551 ( .A(\mem<11><4> ), .B(n1289), .Y(n1698) );
  OAI21X1 U1552 ( .A(n1287), .B(n1327), .C(n1698), .Y(n2082) );
  NAND2X1 U1553 ( .A(\mem<11><5> ), .B(n1289), .Y(n1699) );
  OAI21X1 U1554 ( .A(n1287), .B(n1329), .C(n1699), .Y(n2081) );
  NAND2X1 U1555 ( .A(\mem<11><6> ), .B(n1289), .Y(n1700) );
  OAI21X1 U1556 ( .A(n1287), .B(n1331), .C(n1700), .Y(n2080) );
  NAND2X1 U1557 ( .A(\mem<11><7> ), .B(n1289), .Y(n1701) );
  OAI21X1 U1558 ( .A(n1287), .B(n1333), .C(n1701), .Y(n2079) );
  NAND2X1 U1559 ( .A(\mem<11><8> ), .B(n1290), .Y(n1702) );
  OAI21X1 U1560 ( .A(n1288), .B(n1335), .C(n1702), .Y(n2078) );
  NAND2X1 U1561 ( .A(\mem<11><9> ), .B(n1290), .Y(n1703) );
  OAI21X1 U1562 ( .A(n1288), .B(n1337), .C(n1703), .Y(n2077) );
  NAND2X1 U1563 ( .A(\mem<11><10> ), .B(n1290), .Y(n1704) );
  OAI21X1 U1564 ( .A(n1288), .B(n1339), .C(n1704), .Y(n2076) );
  NAND2X1 U1565 ( .A(\mem<11><11> ), .B(n1290), .Y(n1705) );
  OAI21X1 U1566 ( .A(n1288), .B(n1341), .C(n1705), .Y(n2075) );
  NAND2X1 U1567 ( .A(\mem<11><12> ), .B(n1290), .Y(n1706) );
  OAI21X1 U1568 ( .A(n1288), .B(n1343), .C(n1706), .Y(n2074) );
  NAND2X1 U1569 ( .A(\mem<11><13> ), .B(n1290), .Y(n1707) );
  OAI21X1 U1570 ( .A(n1288), .B(n1345), .C(n1707), .Y(n2073) );
  NAND2X1 U1571 ( .A(\mem<11><14> ), .B(n1290), .Y(n1708) );
  OAI21X1 U1572 ( .A(n1288), .B(n1347), .C(n1708), .Y(n2072) );
  NAND2X1 U1573 ( .A(\mem<11><15> ), .B(n1290), .Y(n1709) );
  OAI21X1 U1574 ( .A(n1288), .B(n1349), .C(n1709), .Y(n2071) );
  NAND2X1 U1575 ( .A(\mem<10><0> ), .B(n1293), .Y(n1710) );
  OAI21X1 U1576 ( .A(n1291), .B(n1320), .C(n1710), .Y(n2070) );
  NAND2X1 U1577 ( .A(\mem<10><1> ), .B(n1293), .Y(n1711) );
  OAI21X1 U1578 ( .A(n1291), .B(n1321), .C(n1711), .Y(n2069) );
  NAND2X1 U1579 ( .A(\mem<10><2> ), .B(n1293), .Y(n1712) );
  OAI21X1 U1580 ( .A(n1291), .B(n1323), .C(n1712), .Y(n2068) );
  NAND2X1 U1581 ( .A(\mem<10><3> ), .B(n1293), .Y(n1713) );
  OAI21X1 U1582 ( .A(n1291), .B(n1325), .C(n1713), .Y(n2067) );
  NAND2X1 U1583 ( .A(\mem<10><4> ), .B(n1293), .Y(n1714) );
  OAI21X1 U1584 ( .A(n1291), .B(n1327), .C(n1714), .Y(n2066) );
  NAND2X1 U1585 ( .A(\mem<10><5> ), .B(n1293), .Y(n1715) );
  OAI21X1 U1586 ( .A(n1291), .B(n1329), .C(n1715), .Y(n2065) );
  NAND2X1 U1587 ( .A(\mem<10><6> ), .B(n1293), .Y(n1716) );
  OAI21X1 U1588 ( .A(n1291), .B(n1331), .C(n1716), .Y(n2064) );
  NAND2X1 U1589 ( .A(\mem<10><7> ), .B(n1293), .Y(n1717) );
  OAI21X1 U1590 ( .A(n1291), .B(n1333), .C(n1717), .Y(n2063) );
  NAND2X1 U1591 ( .A(\mem<10><8> ), .B(n1294), .Y(n1718) );
  OAI21X1 U1592 ( .A(n1292), .B(n1335), .C(n1718), .Y(n2062) );
  NAND2X1 U1593 ( .A(\mem<10><9> ), .B(n1294), .Y(n1719) );
  OAI21X1 U1594 ( .A(n1292), .B(n1337), .C(n1719), .Y(n2061) );
  NAND2X1 U1595 ( .A(\mem<10><10> ), .B(n1294), .Y(n1720) );
  OAI21X1 U1596 ( .A(n1292), .B(n1339), .C(n1720), .Y(n2060) );
  NAND2X1 U1597 ( .A(\mem<10><11> ), .B(n1294), .Y(n1721) );
  OAI21X1 U1598 ( .A(n1292), .B(n1341), .C(n1721), .Y(n2059) );
  NAND2X1 U1599 ( .A(\mem<10><12> ), .B(n1294), .Y(n1722) );
  OAI21X1 U1600 ( .A(n1292), .B(n1343), .C(n1722), .Y(n2058) );
  NAND2X1 U1601 ( .A(\mem<10><13> ), .B(n1294), .Y(n1723) );
  OAI21X1 U1602 ( .A(n1292), .B(n1345), .C(n1723), .Y(n2057) );
  NAND2X1 U1603 ( .A(\mem<10><14> ), .B(n1294), .Y(n1724) );
  OAI21X1 U1604 ( .A(n1292), .B(n1347), .C(n1724), .Y(n2056) );
  NAND2X1 U1605 ( .A(\mem<10><15> ), .B(n1294), .Y(n1725) );
  OAI21X1 U1606 ( .A(n1292), .B(n1349), .C(n1725), .Y(n2055) );
  NAND2X1 U1607 ( .A(\mem<9><0> ), .B(n1297), .Y(n1726) );
  OAI21X1 U1608 ( .A(n1295), .B(n1320), .C(n1726), .Y(n2054) );
  NAND2X1 U1609 ( .A(\mem<9><1> ), .B(n1297), .Y(n1727) );
  OAI21X1 U1610 ( .A(n1295), .B(n1321), .C(n1727), .Y(n2053) );
  NAND2X1 U1611 ( .A(\mem<9><2> ), .B(n1297), .Y(n1728) );
  OAI21X1 U1612 ( .A(n1295), .B(n1323), .C(n1728), .Y(n2052) );
  NAND2X1 U1613 ( .A(\mem<9><3> ), .B(n1297), .Y(n1729) );
  OAI21X1 U1614 ( .A(n1295), .B(n1325), .C(n1729), .Y(n2051) );
  NAND2X1 U1615 ( .A(\mem<9><4> ), .B(n1297), .Y(n1730) );
  OAI21X1 U1616 ( .A(n1295), .B(n1327), .C(n1730), .Y(n2050) );
  NAND2X1 U1617 ( .A(\mem<9><5> ), .B(n1297), .Y(n1731) );
  OAI21X1 U1618 ( .A(n1295), .B(n1329), .C(n1731), .Y(n2049) );
  NAND2X1 U1619 ( .A(\mem<9><6> ), .B(n1297), .Y(n1732) );
  OAI21X1 U1620 ( .A(n1295), .B(n1331), .C(n1732), .Y(n2048) );
  NAND2X1 U1621 ( .A(\mem<9><7> ), .B(n1297), .Y(n1733) );
  OAI21X1 U1622 ( .A(n1295), .B(n1333), .C(n1733), .Y(n2047) );
  NAND2X1 U1623 ( .A(\mem<9><8> ), .B(n1298), .Y(n1734) );
  OAI21X1 U1624 ( .A(n1296), .B(n1335), .C(n1734), .Y(n2046) );
  NAND2X1 U1625 ( .A(\mem<9><9> ), .B(n1298), .Y(n1735) );
  OAI21X1 U1626 ( .A(n1296), .B(n1337), .C(n1735), .Y(n2045) );
  NAND2X1 U1627 ( .A(\mem<9><10> ), .B(n1298), .Y(n1736) );
  OAI21X1 U1628 ( .A(n1296), .B(n1339), .C(n1736), .Y(n2044) );
  NAND2X1 U1629 ( .A(\mem<9><11> ), .B(n1298), .Y(n1737) );
  OAI21X1 U1630 ( .A(n1296), .B(n1341), .C(n1737), .Y(n2043) );
  NAND2X1 U1631 ( .A(\mem<9><12> ), .B(n1298), .Y(n1738) );
  OAI21X1 U1632 ( .A(n1296), .B(n1343), .C(n1738), .Y(n2042) );
  NAND2X1 U1633 ( .A(\mem<9><13> ), .B(n1298), .Y(n1739) );
  OAI21X1 U1634 ( .A(n1296), .B(n1345), .C(n1739), .Y(n2041) );
  NAND2X1 U1635 ( .A(\mem<9><14> ), .B(n1298), .Y(n1740) );
  OAI21X1 U1636 ( .A(n1296), .B(n1347), .C(n1740), .Y(n2040) );
  NAND2X1 U1637 ( .A(\mem<9><15> ), .B(n1298), .Y(n1741) );
  OAI21X1 U1638 ( .A(n1296), .B(n1349), .C(n1741), .Y(n2039) );
  NAND2X1 U1639 ( .A(\mem<8><0> ), .B(n1300), .Y(n1743) );
  OAI21X1 U1640 ( .A(n1299), .B(n1320), .C(n1743), .Y(n2038) );
  NAND2X1 U1641 ( .A(\mem<8><1> ), .B(n1300), .Y(n1744) );
  OAI21X1 U1642 ( .A(n1299), .B(n1321), .C(n1744), .Y(n2037) );
  NAND2X1 U1643 ( .A(\mem<8><2> ), .B(n1300), .Y(n1745) );
  OAI21X1 U1644 ( .A(n1299), .B(n1323), .C(n1745), .Y(n2036) );
  NAND2X1 U1645 ( .A(\mem<8><3> ), .B(n1300), .Y(n1746) );
  OAI21X1 U1646 ( .A(n1299), .B(n1325), .C(n1746), .Y(n2035) );
  NAND2X1 U1647 ( .A(\mem<8><4> ), .B(n1300), .Y(n1747) );
  OAI21X1 U1648 ( .A(n1299), .B(n1327), .C(n1747), .Y(n2034) );
  NAND2X1 U1649 ( .A(\mem<8><5> ), .B(n1300), .Y(n1748) );
  OAI21X1 U1650 ( .A(n1299), .B(n1329), .C(n1748), .Y(n2033) );
  NAND2X1 U1651 ( .A(\mem<8><6> ), .B(n1300), .Y(n1749) );
  OAI21X1 U1652 ( .A(n1299), .B(n1331), .C(n1749), .Y(n2032) );
  NAND2X1 U1653 ( .A(\mem<8><7> ), .B(n1300), .Y(n1750) );
  OAI21X1 U1654 ( .A(n1299), .B(n1333), .C(n1750), .Y(n2031) );
  NAND2X1 U1655 ( .A(\mem<8><8> ), .B(n1301), .Y(n1751) );
  OAI21X1 U1656 ( .A(n1299), .B(n1335), .C(n1751), .Y(n2030) );
  NAND2X1 U1657 ( .A(\mem<8><9> ), .B(n1301), .Y(n1752) );
  OAI21X1 U1658 ( .A(n1299), .B(n1337), .C(n1752), .Y(n2029) );
  NAND2X1 U1659 ( .A(\mem<8><10> ), .B(n1301), .Y(n1753) );
  OAI21X1 U1660 ( .A(n1299), .B(n1339), .C(n1753), .Y(n2028) );
  NAND2X1 U1661 ( .A(\mem<8><11> ), .B(n1301), .Y(n1754) );
  OAI21X1 U1662 ( .A(n1299), .B(n1341), .C(n1754), .Y(n2027) );
  NAND2X1 U1663 ( .A(\mem<8><12> ), .B(n1301), .Y(n1755) );
  OAI21X1 U1664 ( .A(n1299), .B(n1343), .C(n1755), .Y(n2026) );
  NAND2X1 U1665 ( .A(\mem<8><13> ), .B(n1301), .Y(n1756) );
  OAI21X1 U1666 ( .A(n1299), .B(n1345), .C(n1756), .Y(n2025) );
  NAND2X1 U1667 ( .A(\mem<8><14> ), .B(n1301), .Y(n1757) );
  OAI21X1 U1668 ( .A(n1299), .B(n1347), .C(n1757), .Y(n2024) );
  NAND2X1 U1669 ( .A(\mem<8><15> ), .B(n1301), .Y(n1758) );
  OAI21X1 U1670 ( .A(n1299), .B(n1349), .C(n1758), .Y(n2023) );
  NAND3X1 U1671 ( .A(n1358), .B(n2407), .C(n1359), .Y(n1759) );
  NAND2X1 U1672 ( .A(\mem<7><0> ), .B(n1304), .Y(n1760) );
  OAI21X1 U1673 ( .A(n1302), .B(n1320), .C(n1760), .Y(n2022) );
  NAND2X1 U1674 ( .A(\mem<7><1> ), .B(n1304), .Y(n1761) );
  OAI21X1 U1675 ( .A(n1302), .B(n1321), .C(n1761), .Y(n2021) );
  NAND2X1 U1676 ( .A(\mem<7><2> ), .B(n1304), .Y(n1762) );
  OAI21X1 U1677 ( .A(n1302), .B(n1323), .C(n1762), .Y(n2020) );
  NAND2X1 U1678 ( .A(\mem<7><3> ), .B(n1304), .Y(n1763) );
  OAI21X1 U1679 ( .A(n1302), .B(n1325), .C(n1763), .Y(n2019) );
  NAND2X1 U1680 ( .A(\mem<7><4> ), .B(n1304), .Y(n1764) );
  OAI21X1 U1681 ( .A(n1302), .B(n1327), .C(n1764), .Y(n2018) );
  NAND2X1 U1682 ( .A(\mem<7><5> ), .B(n1304), .Y(n1765) );
  OAI21X1 U1683 ( .A(n1302), .B(n1329), .C(n1765), .Y(n2017) );
  NAND2X1 U1684 ( .A(\mem<7><6> ), .B(n1304), .Y(n1766) );
  OAI21X1 U1685 ( .A(n1302), .B(n1331), .C(n1766), .Y(n2016) );
  NAND2X1 U1686 ( .A(\mem<7><7> ), .B(n1304), .Y(n1767) );
  OAI21X1 U1687 ( .A(n1302), .B(n1333), .C(n1767), .Y(n2015) );
  NAND2X1 U1688 ( .A(\mem<7><8> ), .B(n1305), .Y(n1768) );
  OAI21X1 U1689 ( .A(n1303), .B(n1335), .C(n1768), .Y(n2014) );
  NAND2X1 U1690 ( .A(\mem<7><9> ), .B(n1305), .Y(n1769) );
  OAI21X1 U1691 ( .A(n1303), .B(n1337), .C(n1769), .Y(n2013) );
  NAND2X1 U1692 ( .A(\mem<7><10> ), .B(n1305), .Y(n1770) );
  OAI21X1 U1693 ( .A(n1303), .B(n1339), .C(n1770), .Y(n2012) );
  NAND2X1 U1694 ( .A(\mem<7><11> ), .B(n1305), .Y(n1771) );
  OAI21X1 U1695 ( .A(n1303), .B(n1341), .C(n1771), .Y(n2011) );
  NAND2X1 U1696 ( .A(\mem<7><12> ), .B(n1305), .Y(n1772) );
  OAI21X1 U1697 ( .A(n1303), .B(n1343), .C(n1772), .Y(n2010) );
  NAND2X1 U1698 ( .A(\mem<7><13> ), .B(n1305), .Y(n1773) );
  OAI21X1 U1699 ( .A(n1303), .B(n1345), .C(n1773), .Y(n2009) );
  NAND2X1 U1700 ( .A(\mem<7><14> ), .B(n1305), .Y(n1774) );
  OAI21X1 U1701 ( .A(n1303), .B(n1347), .C(n1774), .Y(n2008) );
  NAND2X1 U1702 ( .A(\mem<7><15> ), .B(n1305), .Y(n1775) );
  OAI21X1 U1703 ( .A(n1303), .B(n1349), .C(n1775), .Y(n2007) );
  NAND2X1 U1704 ( .A(\mem<6><0> ), .B(n150), .Y(n1776) );
  OAI21X1 U1705 ( .A(n1306), .B(n1320), .C(n1776), .Y(n2006) );
  NAND2X1 U1706 ( .A(\mem<6><1> ), .B(n150), .Y(n1777) );
  OAI21X1 U1707 ( .A(n1306), .B(n1321), .C(n1777), .Y(n2005) );
  NAND2X1 U1708 ( .A(\mem<6><2> ), .B(n150), .Y(n1778) );
  OAI21X1 U1709 ( .A(n1306), .B(n1323), .C(n1778), .Y(n2004) );
  NAND2X1 U1710 ( .A(\mem<6><3> ), .B(n150), .Y(n1779) );
  OAI21X1 U1711 ( .A(n1306), .B(n1325), .C(n1779), .Y(n2003) );
  NAND2X1 U1712 ( .A(\mem<6><4> ), .B(n150), .Y(n1780) );
  OAI21X1 U1713 ( .A(n1306), .B(n1327), .C(n1780), .Y(n2002) );
  NAND2X1 U1714 ( .A(\mem<6><5> ), .B(n150), .Y(n1781) );
  OAI21X1 U1715 ( .A(n1306), .B(n1329), .C(n1781), .Y(n2001) );
  NAND2X1 U1716 ( .A(\mem<6><6> ), .B(n150), .Y(n1782) );
  OAI21X1 U1717 ( .A(n1306), .B(n1331), .C(n1782), .Y(n2000) );
  NAND2X1 U1718 ( .A(\mem<6><7> ), .B(n150), .Y(n1783) );
  OAI21X1 U1719 ( .A(n1306), .B(n1333), .C(n1783), .Y(n1999) );
  NAND2X1 U1720 ( .A(\mem<6><8> ), .B(n150), .Y(n1784) );
  OAI21X1 U1721 ( .A(n1307), .B(n1335), .C(n1784), .Y(n1998) );
  NAND2X1 U1722 ( .A(\mem<6><9> ), .B(n150), .Y(n1785) );
  OAI21X1 U1723 ( .A(n1307), .B(n1337), .C(n1785), .Y(n1997) );
  NAND2X1 U1724 ( .A(\mem<6><10> ), .B(n150), .Y(n1786) );
  OAI21X1 U1725 ( .A(n1307), .B(n1339), .C(n1786), .Y(n1996) );
  NAND2X1 U1726 ( .A(\mem<6><11> ), .B(n150), .Y(n1787) );
  OAI21X1 U1727 ( .A(n1307), .B(n1341), .C(n1787), .Y(n1995) );
  NAND2X1 U1728 ( .A(\mem<6><12> ), .B(n150), .Y(n1788) );
  OAI21X1 U1729 ( .A(n1307), .B(n1343), .C(n1788), .Y(n1994) );
  NAND2X1 U1730 ( .A(\mem<6><13> ), .B(n150), .Y(n1789) );
  OAI21X1 U1731 ( .A(n1307), .B(n1345), .C(n1789), .Y(n1993) );
  NAND2X1 U1732 ( .A(\mem<6><14> ), .B(n150), .Y(n1790) );
  OAI21X1 U1733 ( .A(n1307), .B(n1347), .C(n1790), .Y(n1992) );
  NAND2X1 U1734 ( .A(\mem<6><15> ), .B(n150), .Y(n1791) );
  OAI21X1 U1735 ( .A(n1307), .B(n1349), .C(n1791), .Y(n1991) );
  NAND2X1 U1736 ( .A(\mem<5><0> ), .B(n153), .Y(n1793) );
  OAI21X1 U1737 ( .A(n1308), .B(n1320), .C(n1793), .Y(n1990) );
  NAND2X1 U1738 ( .A(\mem<5><1> ), .B(n153), .Y(n1794) );
  OAI21X1 U1739 ( .A(n1308), .B(n1321), .C(n1794), .Y(n1989) );
  NAND2X1 U1740 ( .A(\mem<5><2> ), .B(n153), .Y(n1795) );
  OAI21X1 U1741 ( .A(n1308), .B(n1323), .C(n1795), .Y(n1988) );
  NAND2X1 U1742 ( .A(\mem<5><3> ), .B(n153), .Y(n1796) );
  OAI21X1 U1743 ( .A(n1308), .B(n1325), .C(n1796), .Y(n1987) );
  NAND2X1 U1744 ( .A(\mem<5><4> ), .B(n153), .Y(n1797) );
  OAI21X1 U1745 ( .A(n1308), .B(n1327), .C(n1797), .Y(n1986) );
  NAND2X1 U1746 ( .A(\mem<5><5> ), .B(n153), .Y(n1798) );
  OAI21X1 U1747 ( .A(n1308), .B(n1329), .C(n1798), .Y(n1985) );
  NAND2X1 U1748 ( .A(\mem<5><6> ), .B(n153), .Y(n1799) );
  OAI21X1 U1749 ( .A(n1308), .B(n1331), .C(n1799), .Y(n1984) );
  NAND2X1 U1750 ( .A(\mem<5><7> ), .B(n153), .Y(n1800) );
  OAI21X1 U1751 ( .A(n1308), .B(n1333), .C(n1800), .Y(n1983) );
  NAND2X1 U1752 ( .A(\mem<5><8> ), .B(n153), .Y(n1801) );
  OAI21X1 U1753 ( .A(n1309), .B(n1335), .C(n1801), .Y(n1982) );
  NAND2X1 U1754 ( .A(\mem<5><9> ), .B(n153), .Y(n1802) );
  OAI21X1 U1755 ( .A(n1309), .B(n1337), .C(n1802), .Y(n1981) );
  NAND2X1 U1756 ( .A(\mem<5><10> ), .B(n153), .Y(n1803) );
  OAI21X1 U1757 ( .A(n1309), .B(n1339), .C(n1803), .Y(n1980) );
  NAND2X1 U1758 ( .A(\mem<5><11> ), .B(n153), .Y(n1804) );
  OAI21X1 U1759 ( .A(n1309), .B(n1341), .C(n1804), .Y(n1979) );
  NAND2X1 U1760 ( .A(\mem<5><12> ), .B(n153), .Y(n1805) );
  OAI21X1 U1761 ( .A(n1309), .B(n1343), .C(n1805), .Y(n1978) );
  NAND2X1 U1762 ( .A(\mem<5><13> ), .B(n153), .Y(n1806) );
  OAI21X1 U1763 ( .A(n1309), .B(n1345), .C(n1806), .Y(n1977) );
  NAND2X1 U1764 ( .A(\mem<5><14> ), .B(n153), .Y(n1807) );
  OAI21X1 U1765 ( .A(n1309), .B(n1347), .C(n1807), .Y(n1976) );
  NAND2X1 U1766 ( .A(\mem<5><15> ), .B(n153), .Y(n1808) );
  OAI21X1 U1767 ( .A(n1309), .B(n1349), .C(n1808), .Y(n1975) );
  NAND2X1 U1768 ( .A(\mem<4><0> ), .B(n156), .Y(n1810) );
  OAI21X1 U1769 ( .A(n1310), .B(n1320), .C(n1810), .Y(n1974) );
  NAND2X1 U1770 ( .A(\mem<4><1> ), .B(n156), .Y(n1811) );
  OAI21X1 U1771 ( .A(n1310), .B(n1321), .C(n1811), .Y(n1973) );
  NAND2X1 U1772 ( .A(\mem<4><2> ), .B(n156), .Y(n1812) );
  OAI21X1 U1773 ( .A(n1310), .B(n1323), .C(n1812), .Y(n1972) );
  NAND2X1 U1774 ( .A(\mem<4><3> ), .B(n156), .Y(n1813) );
  OAI21X1 U1775 ( .A(n1310), .B(n1325), .C(n1813), .Y(n1971) );
  NAND2X1 U1776 ( .A(\mem<4><4> ), .B(n156), .Y(n1814) );
  OAI21X1 U1777 ( .A(n1310), .B(n1327), .C(n1814), .Y(n1970) );
  NAND2X1 U1778 ( .A(\mem<4><5> ), .B(n156), .Y(n1815) );
  OAI21X1 U1779 ( .A(n1310), .B(n1329), .C(n1815), .Y(n1969) );
  NAND2X1 U1780 ( .A(\mem<4><6> ), .B(n156), .Y(n1816) );
  OAI21X1 U1781 ( .A(n1310), .B(n1331), .C(n1816), .Y(n1968) );
  NAND2X1 U1782 ( .A(\mem<4><7> ), .B(n156), .Y(n1817) );
  OAI21X1 U1783 ( .A(n1310), .B(n1333), .C(n1817), .Y(n1967) );
  NAND2X1 U1784 ( .A(\mem<4><8> ), .B(n156), .Y(n1818) );
  OAI21X1 U1785 ( .A(n1311), .B(n1335), .C(n1818), .Y(n1966) );
  NAND2X1 U1786 ( .A(\mem<4><9> ), .B(n156), .Y(n1819) );
  OAI21X1 U1787 ( .A(n1311), .B(n1337), .C(n1819), .Y(n1965) );
  NAND2X1 U1788 ( .A(\mem<4><10> ), .B(n156), .Y(n1820) );
  OAI21X1 U1789 ( .A(n1311), .B(n1339), .C(n1820), .Y(n1964) );
  NAND2X1 U1790 ( .A(\mem<4><11> ), .B(n156), .Y(n1821) );
  OAI21X1 U1791 ( .A(n1311), .B(n1341), .C(n1821), .Y(n1963) );
  NAND2X1 U1792 ( .A(\mem<4><12> ), .B(n156), .Y(n1822) );
  OAI21X1 U1793 ( .A(n1311), .B(n1343), .C(n1822), .Y(n1962) );
  NAND2X1 U1794 ( .A(\mem<4><13> ), .B(n156), .Y(n1823) );
  OAI21X1 U1795 ( .A(n1311), .B(n1345), .C(n1823), .Y(n1961) );
  NAND2X1 U1796 ( .A(\mem<4><14> ), .B(n156), .Y(n1824) );
  OAI21X1 U1797 ( .A(n1311), .B(n1347), .C(n1824), .Y(n1960) );
  NAND2X1 U1798 ( .A(\mem<4><15> ), .B(n156), .Y(n1825) );
  OAI21X1 U1799 ( .A(n1311), .B(n1349), .C(n1825), .Y(n1959) );
  NAND2X1 U1800 ( .A(\mem<3><0> ), .B(n159), .Y(n1827) );
  OAI21X1 U1801 ( .A(n1312), .B(n1320), .C(n1827), .Y(n1958) );
  NAND2X1 U1802 ( .A(\mem<3><1> ), .B(n159), .Y(n1828) );
  OAI21X1 U1803 ( .A(n1312), .B(n1321), .C(n1828), .Y(n1957) );
  NAND2X1 U1804 ( .A(\mem<3><2> ), .B(n159), .Y(n1829) );
  OAI21X1 U1805 ( .A(n1312), .B(n1323), .C(n1829), .Y(n1956) );
  NAND2X1 U1806 ( .A(\mem<3><3> ), .B(n159), .Y(n1830) );
  OAI21X1 U1807 ( .A(n1312), .B(n1325), .C(n1830), .Y(n1955) );
  NAND2X1 U1808 ( .A(\mem<3><4> ), .B(n159), .Y(n1831) );
  OAI21X1 U1809 ( .A(n1312), .B(n1327), .C(n1831), .Y(n1954) );
  NAND2X1 U1810 ( .A(\mem<3><5> ), .B(n159), .Y(n1832) );
  OAI21X1 U1811 ( .A(n1312), .B(n1329), .C(n1832), .Y(n1953) );
  NAND2X1 U1812 ( .A(\mem<3><6> ), .B(n159), .Y(n1833) );
  OAI21X1 U1813 ( .A(n1312), .B(n1331), .C(n1833), .Y(n1952) );
  NAND2X1 U1814 ( .A(\mem<3><7> ), .B(n159), .Y(n1834) );
  OAI21X1 U1815 ( .A(n1312), .B(n1333), .C(n1834), .Y(n1951) );
  NAND2X1 U1816 ( .A(\mem<3><8> ), .B(n159), .Y(n1835) );
  OAI21X1 U1817 ( .A(n1313), .B(n1335), .C(n1835), .Y(n1950) );
  NAND2X1 U1818 ( .A(\mem<3><9> ), .B(n159), .Y(n1836) );
  OAI21X1 U1819 ( .A(n1313), .B(n1337), .C(n1836), .Y(n1949) );
  NAND2X1 U1820 ( .A(\mem<3><10> ), .B(n159), .Y(n1837) );
  OAI21X1 U1821 ( .A(n1313), .B(n1339), .C(n1837), .Y(n1948) );
  NAND2X1 U1822 ( .A(\mem<3><11> ), .B(n159), .Y(n1838) );
  OAI21X1 U1823 ( .A(n1313), .B(n1341), .C(n1838), .Y(n1947) );
  NAND2X1 U1824 ( .A(\mem<3><12> ), .B(n159), .Y(n1839) );
  OAI21X1 U1825 ( .A(n1313), .B(n1343), .C(n1839), .Y(n1946) );
  NAND2X1 U1826 ( .A(\mem<3><13> ), .B(n159), .Y(n1840) );
  OAI21X1 U1827 ( .A(n1313), .B(n1345), .C(n1840), .Y(n1945) );
  NAND2X1 U1828 ( .A(\mem<3><14> ), .B(n159), .Y(n1841) );
  OAI21X1 U1829 ( .A(n1313), .B(n1347), .C(n1841), .Y(n1944) );
  NAND2X1 U1830 ( .A(\mem<3><15> ), .B(n159), .Y(n1842) );
  OAI21X1 U1831 ( .A(n1313), .B(n1349), .C(n1842), .Y(n1943) );
  NAND2X1 U1832 ( .A(\mem<2><0> ), .B(n162), .Y(n1844) );
  OAI21X1 U1833 ( .A(n1314), .B(n1320), .C(n1844), .Y(n1942) );
  NAND2X1 U1834 ( .A(\mem<2><1> ), .B(n162), .Y(n1845) );
  OAI21X1 U1835 ( .A(n1314), .B(n1321), .C(n1845), .Y(n1941) );
  NAND2X1 U1836 ( .A(\mem<2><2> ), .B(n162), .Y(n1846) );
  OAI21X1 U1837 ( .A(n1314), .B(n1323), .C(n1846), .Y(n1940) );
  NAND2X1 U1838 ( .A(\mem<2><3> ), .B(n162), .Y(n1847) );
  OAI21X1 U1839 ( .A(n1314), .B(n1325), .C(n1847), .Y(n1939) );
  NAND2X1 U1840 ( .A(\mem<2><4> ), .B(n162), .Y(n1848) );
  OAI21X1 U1841 ( .A(n1314), .B(n1327), .C(n1848), .Y(n1938) );
  NAND2X1 U1842 ( .A(\mem<2><5> ), .B(n162), .Y(n1849) );
  OAI21X1 U1843 ( .A(n1314), .B(n1329), .C(n1849), .Y(n1937) );
  NAND2X1 U1844 ( .A(\mem<2><6> ), .B(n162), .Y(n1850) );
  OAI21X1 U1845 ( .A(n1314), .B(n1331), .C(n1850), .Y(n1936) );
  NAND2X1 U1846 ( .A(\mem<2><7> ), .B(n162), .Y(n1851) );
  OAI21X1 U1847 ( .A(n1314), .B(n1333), .C(n1851), .Y(n1935) );
  NAND2X1 U1848 ( .A(\mem<2><8> ), .B(n162), .Y(n1852) );
  OAI21X1 U1849 ( .A(n1315), .B(n1335), .C(n1852), .Y(n1934) );
  NAND2X1 U1850 ( .A(\mem<2><9> ), .B(n162), .Y(n1853) );
  OAI21X1 U1851 ( .A(n1315), .B(n1337), .C(n1853), .Y(n1933) );
  NAND2X1 U1852 ( .A(\mem<2><10> ), .B(n162), .Y(n1854) );
  OAI21X1 U1853 ( .A(n1315), .B(n1339), .C(n1854), .Y(n1932) );
  NAND2X1 U1854 ( .A(\mem<2><11> ), .B(n162), .Y(n1855) );
  OAI21X1 U1855 ( .A(n1315), .B(n1341), .C(n1855), .Y(n1931) );
  NAND2X1 U1856 ( .A(\mem<2><12> ), .B(n162), .Y(n1856) );
  OAI21X1 U1857 ( .A(n1315), .B(n1343), .C(n1856), .Y(n1930) );
  NAND2X1 U1858 ( .A(\mem<2><13> ), .B(n162), .Y(n1857) );
  OAI21X1 U1859 ( .A(n1315), .B(n1345), .C(n1857), .Y(n1929) );
  NAND2X1 U1860 ( .A(\mem<2><14> ), .B(n162), .Y(n1858) );
  OAI21X1 U1861 ( .A(n1315), .B(n1347), .C(n1858), .Y(n1928) );
  NAND2X1 U1862 ( .A(\mem<2><15> ), .B(n162), .Y(n1859) );
  OAI21X1 U1863 ( .A(n1315), .B(n1349), .C(n1859), .Y(n1927) );
  NAND2X1 U1864 ( .A(\mem<1><0> ), .B(n165), .Y(n1861) );
  OAI21X1 U1865 ( .A(n1316), .B(n1320), .C(n1861), .Y(n1926) );
  NAND2X1 U1866 ( .A(\mem<1><1> ), .B(n165), .Y(n1862) );
  OAI21X1 U1867 ( .A(n1316), .B(n1321), .C(n1862), .Y(n1925) );
  NAND2X1 U1868 ( .A(\mem<1><2> ), .B(n165), .Y(n1863) );
  OAI21X1 U1869 ( .A(n1316), .B(n1323), .C(n1863), .Y(n1924) );
  NAND2X1 U1870 ( .A(\mem<1><3> ), .B(n165), .Y(n1864) );
  OAI21X1 U1871 ( .A(n1316), .B(n1325), .C(n1864), .Y(n1923) );
  NAND2X1 U1872 ( .A(\mem<1><4> ), .B(n165), .Y(n1865) );
  OAI21X1 U1873 ( .A(n1316), .B(n1327), .C(n1865), .Y(n1922) );
  NAND2X1 U1874 ( .A(\mem<1><5> ), .B(n165), .Y(n1866) );
  OAI21X1 U1875 ( .A(n1316), .B(n1329), .C(n1866), .Y(n1921) );
  NAND2X1 U1876 ( .A(\mem<1><6> ), .B(n165), .Y(n1867) );
  OAI21X1 U1877 ( .A(n1316), .B(n1331), .C(n1867), .Y(n1920) );
  NAND2X1 U1878 ( .A(\mem<1><7> ), .B(n165), .Y(n1868) );
  OAI21X1 U1879 ( .A(n1316), .B(n1333), .C(n1868), .Y(n1919) );
  NAND2X1 U1880 ( .A(\mem<1><8> ), .B(n165), .Y(n1869) );
  OAI21X1 U1881 ( .A(n1317), .B(n1335), .C(n1869), .Y(n1918) );
  NAND2X1 U1882 ( .A(\mem<1><9> ), .B(n165), .Y(n1870) );
  OAI21X1 U1883 ( .A(n1317), .B(n1337), .C(n1870), .Y(n1917) );
  NAND2X1 U1884 ( .A(\mem<1><10> ), .B(n165), .Y(n1871) );
  OAI21X1 U1885 ( .A(n1317), .B(n1339), .C(n1871), .Y(n1916) );
  NAND2X1 U1886 ( .A(\mem<1><11> ), .B(n165), .Y(n1872) );
  OAI21X1 U1887 ( .A(n1317), .B(n1341), .C(n1872), .Y(n1915) );
  NAND2X1 U1888 ( .A(\mem<1><12> ), .B(n165), .Y(n1873) );
  OAI21X1 U1889 ( .A(n1317), .B(n1343), .C(n1873), .Y(n1914) );
  NAND2X1 U1890 ( .A(\mem<1><13> ), .B(n165), .Y(n1874) );
  OAI21X1 U1891 ( .A(n1317), .B(n1345), .C(n1874), .Y(n1913) );
  NAND2X1 U1892 ( .A(\mem<1><14> ), .B(n165), .Y(n1875) );
  OAI21X1 U1893 ( .A(n1317), .B(n1347), .C(n1875), .Y(n1912) );
  NAND2X1 U1894 ( .A(\mem<1><15> ), .B(n165), .Y(n1876) );
  OAI21X1 U1895 ( .A(n1317), .B(n1349), .C(n1876), .Y(n1911) );
  NAND2X1 U1896 ( .A(\mem<0><0> ), .B(n166), .Y(n1879) );
  OAI21X1 U1897 ( .A(n1318), .B(n1320), .C(n1879), .Y(n1910) );
  NAND2X1 U1898 ( .A(\mem<0><1> ), .B(n166), .Y(n1880) );
  OAI21X1 U1899 ( .A(n1318), .B(n1321), .C(n1880), .Y(n1909) );
  NAND2X1 U1900 ( .A(\mem<0><2> ), .B(n166), .Y(n1881) );
  OAI21X1 U1901 ( .A(n1318), .B(n1323), .C(n1881), .Y(n1908) );
  NAND2X1 U1902 ( .A(\mem<0><3> ), .B(n166), .Y(n1882) );
  OAI21X1 U1903 ( .A(n1318), .B(n1325), .C(n1882), .Y(n1907) );
  NAND2X1 U1904 ( .A(\mem<0><4> ), .B(n166), .Y(n1883) );
  OAI21X1 U1905 ( .A(n1318), .B(n1327), .C(n1883), .Y(n1906) );
  NAND2X1 U1906 ( .A(\mem<0><5> ), .B(n166), .Y(n1884) );
  OAI21X1 U1907 ( .A(n1318), .B(n1329), .C(n1884), .Y(n1905) );
  NAND2X1 U1908 ( .A(\mem<0><6> ), .B(n166), .Y(n1885) );
  OAI21X1 U1909 ( .A(n1318), .B(n1331), .C(n1885), .Y(n1904) );
  NAND2X1 U1910 ( .A(\mem<0><7> ), .B(n166), .Y(n1886) );
  OAI21X1 U1911 ( .A(n1318), .B(n1333), .C(n1886), .Y(n1903) );
  NAND2X1 U1912 ( .A(\mem<0><8> ), .B(n166), .Y(n1887) );
  OAI21X1 U1913 ( .A(n1318), .B(n1335), .C(n1887), .Y(n1902) );
  NAND2X1 U1914 ( .A(\mem<0><9> ), .B(n166), .Y(n1888) );
  OAI21X1 U1915 ( .A(n1318), .B(n1337), .C(n1888), .Y(n1901) );
  NAND2X1 U1916 ( .A(\mem<0><10> ), .B(n166), .Y(n1889) );
  OAI21X1 U1917 ( .A(n1318), .B(n1339), .C(n1889), .Y(n1900) );
  NAND2X1 U1918 ( .A(\mem<0><11> ), .B(n166), .Y(n1890) );
  OAI21X1 U1919 ( .A(n1318), .B(n1341), .C(n1890), .Y(n1899) );
  NAND2X1 U1920 ( .A(\mem<0><12> ), .B(n166), .Y(n1891) );
  OAI21X1 U1921 ( .A(n1318), .B(n1343), .C(n1891), .Y(n1898) );
  NAND2X1 U1922 ( .A(\mem<0><13> ), .B(n166), .Y(n1892) );
  OAI21X1 U1923 ( .A(n1318), .B(n1345), .C(n1892), .Y(n1897) );
  NAND2X1 U1924 ( .A(\mem<0><14> ), .B(n166), .Y(n1893) );
  OAI21X1 U1925 ( .A(n1318), .B(n1347), .C(n1893), .Y(n1896) );
  NAND2X1 U1926 ( .A(\mem<0><15> ), .B(n166), .Y(n1894) );
  OAI21X1 U1927 ( .A(n1318), .B(n1349), .C(n1894), .Y(n1895) );
endmodule


module memc_Size5_0 ( .data_out({\data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        write, clk, rst, createdump, .file_id({\file_id<4> , \file_id<3> , 
        \file_id<2> , \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<4> , \data_in<3> , \data_in<2> ,
         \data_in<1> , \data_in<0> , write, clk, rst, createdump, \file_id<4> ,
         \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> ,
         \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><4> , \mem<0><3> , \mem<0><2> ,
         \mem<0><1> , \mem<0><0> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><4> , \mem<3><3> , \mem<3><2> ,
         \mem<3><1> , \mem<3><0> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><4> , \mem<5><3> , \mem<5><2> ,
         \mem<5><1> , \mem<5><0> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><4> , \mem<8><3> , \mem<8><2> ,
         \mem<8><1> , \mem<8><0> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><4> , \mem<10><3> , \mem<10><2> ,
         \mem<10><1> , \mem<10><0> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><4> , \mem<13><3> , \mem<13><2> ,
         \mem<13><1> , \mem<13><0> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><4> , \mem<15><3> , \mem<15><2> ,
         \mem<15><1> , \mem<15><0> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><4> , \mem<18><3> , \mem<18><2> ,
         \mem<18><1> , \mem<18><0> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><4> , \mem<20><3> , \mem<20><2> ,
         \mem<20><1> , \mem<20><0> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><4> , \mem<23><3> , \mem<23><2> ,
         \mem<23><1> , \mem<23><0> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><4> , \mem<25><3> , \mem<25><2> ,
         \mem<25><1> , \mem<25><0> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><4> , \mem<28><3> , \mem<28><2> ,
         \mem<28><1> , \mem<28><0> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><4> , \mem<30><3> , \mem<30><2> ,
         \mem<30><1> , \mem<30><0> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , N17, N18, N19, N20, N21, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n58, n59, n60, n61, n62, n63,
         n64, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79,
         n80, n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n106, n107, n108, n109,
         n110, n111, n112, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n287, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><4>  ( .D(n831), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n832), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n833), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n834), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n835), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n836), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n837), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n838), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n839), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n840), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n841), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n842), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n843), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n844), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n845), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n846), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n847), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n848), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n849), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n850), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n851), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n852), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n853), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n854), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n855), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n856), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n857), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n858), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n859), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n860), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n861), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n862), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n863), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n864), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n865), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n866), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n867), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n868), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n869), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n870), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n871), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n872), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n873), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n874), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n875), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n876), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n877), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n878), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n879), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n880), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n881), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n882), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n883), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n884), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n885), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n886), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n887), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n888), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n889), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n890), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n891), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n892), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n893), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n894), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n895), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n896), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n897), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n898), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n899), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n900), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n901), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n902), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n903), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n904), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n905), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n906), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n907), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n908), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n909), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n910), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n911), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n912), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n913), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n914), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n915), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n916), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n917), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n918), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n919), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n920), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n921), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n922), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n923), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n924), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n925), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n926), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n927), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n928), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n929), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n930), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n931), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n932), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n933), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n934), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n935), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n936), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n937), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n938), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n939), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n940), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n941), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n942), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n943), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n944), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n945), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n946), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n947), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n948), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n949), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n950), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n951), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n952), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n953), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n954), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n955), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n956), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n957), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n958), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n959), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n960), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n961), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n962), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n963), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n964), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n965), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n966), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n967), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n968), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n969), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n970), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n971), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n972), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n973), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n974), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n975), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n976), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n977), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n978), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n979), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n980), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n981), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n982), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n983), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n984), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n985), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n986), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n987), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n988), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n989), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n990), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(n647), .B(n820), .Y(n1004) );
  OAI21X1 U50 ( .A(n578), .B(n819), .C(n212), .Y(n990) );
  OAI21X1 U52 ( .A(n578), .B(n818), .C(n210), .Y(n989) );
  OAI21X1 U54 ( .A(n578), .B(n817), .C(n208), .Y(n988) );
  OAI21X1 U56 ( .A(n578), .B(n816), .C(n206), .Y(n987) );
  OAI21X1 U58 ( .A(n578), .B(n815), .C(n204), .Y(n986) );
  OAI21X1 U62 ( .A(n819), .B(n641), .C(n202), .Y(n985) );
  OAI21X1 U64 ( .A(n818), .B(n641), .C(n200), .Y(n984) );
  OAI21X1 U66 ( .A(n817), .B(n641), .C(n198), .Y(n983) );
  OAI21X1 U68 ( .A(n816), .B(n641), .C(n196), .Y(n982) );
  OAI21X1 U70 ( .A(n815), .B(n641), .C(n194), .Y(n981) );
  OAI21X1 U74 ( .A(n819), .B(n639), .C(n192), .Y(n980) );
  OAI21X1 U76 ( .A(n818), .B(n639), .C(n190), .Y(n979) );
  OAI21X1 U78 ( .A(n817), .B(n639), .C(n188), .Y(n978) );
  OAI21X1 U80 ( .A(n816), .B(n639), .C(n186), .Y(n977) );
  OAI21X1 U82 ( .A(n815), .B(n639), .C(n184), .Y(n976) );
  OAI21X1 U86 ( .A(n819), .B(n637), .C(n182), .Y(n975) );
  OAI21X1 U88 ( .A(n818), .B(n637), .C(n180), .Y(n974) );
  OAI21X1 U90 ( .A(n817), .B(n637), .C(n178), .Y(n973) );
  OAI21X1 U92 ( .A(n816), .B(n637), .C(n176), .Y(n972) );
  OAI21X1 U94 ( .A(n815), .B(n637), .C(n174), .Y(n971) );
  OAI21X1 U98 ( .A(n819), .B(n635), .C(n171), .Y(n970) );
  OAI21X1 U100 ( .A(n818), .B(n635), .C(n169), .Y(n969) );
  OAI21X1 U102 ( .A(n817), .B(n635), .C(n167), .Y(n968) );
  OAI21X1 U104 ( .A(n816), .B(n635), .C(n165), .Y(n967) );
  OAI21X1 U106 ( .A(n815), .B(n635), .C(n163), .Y(n966) );
  OAI21X1 U110 ( .A(n819), .B(n633), .C(n497), .Y(n965) );
  OAI21X1 U112 ( .A(n818), .B(n633), .C(n495), .Y(n964) );
  OAI21X1 U114 ( .A(n817), .B(n633), .C(n493), .Y(n963) );
  OAI21X1 U116 ( .A(n816), .B(n633), .C(n491), .Y(n962) );
  OAI21X1 U118 ( .A(n815), .B(n633), .C(n161), .Y(n961) );
  OAI21X1 U122 ( .A(n819), .B(n631), .C(n159), .Y(n960) );
  OAI21X1 U124 ( .A(n818), .B(n631), .C(n157), .Y(n959) );
  OAI21X1 U126 ( .A(n817), .B(n631), .C(n155), .Y(n958) );
  OAI21X1 U128 ( .A(n816), .B(n631), .C(n153), .Y(n957) );
  OAI21X1 U130 ( .A(n815), .B(n631), .C(n151), .Y(n956) );
  OAI21X1 U134 ( .A(n819), .B(n629), .C(n489), .Y(n955) );
  OAI21X1 U136 ( .A(n818), .B(n629), .C(n487), .Y(n954) );
  OAI21X1 U138 ( .A(n817), .B(n629), .C(n485), .Y(n953) );
  OAI21X1 U140 ( .A(n816), .B(n629), .C(n483), .Y(n952) );
  OAI21X1 U142 ( .A(n815), .B(n629), .C(n149), .Y(n951) );
  NAND3X1 U146 ( .A(N13), .B(n994), .C(N14), .Y(n995) );
  OAI21X1 U147 ( .A(n819), .B(n626), .C(n147), .Y(n950) );
  OAI21X1 U149 ( .A(n818), .B(n626), .C(n145), .Y(n949) );
  OAI21X1 U151 ( .A(n817), .B(n626), .C(n143), .Y(n948) );
  OAI21X1 U153 ( .A(n816), .B(n626), .C(n141), .Y(n947) );
  OAI21X1 U155 ( .A(n815), .B(n626), .C(n139), .Y(n946) );
  OAI21X1 U159 ( .A(n819), .B(n624), .C(n137), .Y(n945) );
  OAI21X1 U161 ( .A(n818), .B(n624), .C(n135), .Y(n944) );
  OAI21X1 U163 ( .A(n817), .B(n624), .C(n133), .Y(n943) );
  OAI21X1 U165 ( .A(n816), .B(n624), .C(n131), .Y(n942) );
  OAI21X1 U167 ( .A(n815), .B(n624), .C(n129), .Y(n941) );
  OAI21X1 U171 ( .A(n819), .B(n622), .C(n127), .Y(n940) );
  OAI21X1 U173 ( .A(n818), .B(n622), .C(n125), .Y(n939) );
  OAI21X1 U175 ( .A(n817), .B(n622), .C(n123), .Y(n938) );
  OAI21X1 U177 ( .A(n816), .B(n622), .C(n121), .Y(n937) );
  OAI21X1 U179 ( .A(n815), .B(n622), .C(n119), .Y(n936) );
  OAI21X1 U183 ( .A(n819), .B(n621), .C(n117), .Y(n935) );
  OAI21X1 U185 ( .A(n818), .B(n621), .C(n112), .Y(n934) );
  OAI21X1 U187 ( .A(n817), .B(n621), .C(n110), .Y(n933) );
  OAI21X1 U189 ( .A(n816), .B(n621), .C(n108), .Y(n932) );
  OAI21X1 U191 ( .A(n815), .B(n621), .C(n106), .Y(n931) );
  OAI21X1 U195 ( .A(n819), .B(n618), .C(n103), .Y(n930) );
  OAI21X1 U197 ( .A(n818), .B(n618), .C(n101), .Y(n929) );
  OAI21X1 U199 ( .A(n817), .B(n618), .C(n99), .Y(n928) );
  OAI21X1 U201 ( .A(n816), .B(n618), .C(n96), .Y(n927) );
  OAI21X1 U203 ( .A(n815), .B(n618), .C(n94), .Y(n926) );
  OAI21X1 U207 ( .A(n819), .B(n617), .C(n481), .Y(n925) );
  OAI21X1 U209 ( .A(n818), .B(n617), .C(n479), .Y(n924) );
  OAI21X1 U211 ( .A(n817), .B(n617), .C(n477), .Y(n923) );
  OAI21X1 U213 ( .A(n816), .B(n617), .C(n475), .Y(n922) );
  OAI21X1 U215 ( .A(n815), .B(n617), .C(n92), .Y(n921) );
  OAI21X1 U219 ( .A(n819), .B(n615), .C(n90), .Y(n920) );
  OAI21X1 U221 ( .A(n818), .B(n615), .C(n87), .Y(n919) );
  OAI21X1 U223 ( .A(n817), .B(n615), .C(n85), .Y(n918) );
  OAI21X1 U225 ( .A(n816), .B(n615), .C(n83), .Y(n917) );
  OAI21X1 U227 ( .A(n815), .B(n615), .C(n80), .Y(n916) );
  OAI21X1 U231 ( .A(n819), .B(n613), .C(n473), .Y(n915) );
  OAI21X1 U233 ( .A(n818), .B(n613), .C(n471), .Y(n914) );
  OAI21X1 U235 ( .A(n817), .B(n613), .C(n469), .Y(n913) );
  OAI21X1 U237 ( .A(n816), .B(n613), .C(n467), .Y(n912) );
  OAI21X1 U239 ( .A(n815), .B(n613), .C(n78), .Y(n911) );
  NAND3X1 U243 ( .A(n994), .B(n646), .C(N14), .Y(n993) );
  OAI21X1 U244 ( .A(n819), .B(n610), .C(n76), .Y(n910) );
  OAI21X1 U246 ( .A(n818), .B(n610), .C(n74), .Y(n909) );
  OAI21X1 U248 ( .A(n817), .B(n610), .C(n465), .Y(n908) );
  OAI21X1 U250 ( .A(n816), .B(n610), .C(n463), .Y(n907) );
  OAI21X1 U252 ( .A(n815), .B(n610), .C(n71), .Y(n906) );
  OAI21X1 U256 ( .A(n819), .B(n608), .C(n461), .Y(n905) );
  OAI21X1 U258 ( .A(n818), .B(n608), .C(n459), .Y(n904) );
  OAI21X1 U260 ( .A(n817), .B(n608), .C(n69), .Y(n903) );
  OAI21X1 U262 ( .A(n816), .B(n608), .C(n67), .Y(n902) );
  OAI21X1 U264 ( .A(n815), .B(n608), .C(n64), .Y(n901) );
  OAI21X1 U268 ( .A(n819), .B(n606), .C(n62), .Y(n900) );
  OAI21X1 U270 ( .A(n818), .B(n606), .C(n60), .Y(n899) );
  OAI21X1 U272 ( .A(n817), .B(n606), .C(n58), .Y(n898) );
  OAI21X1 U274 ( .A(n816), .B(n606), .C(n54), .Y(n897) );
  OAI21X1 U276 ( .A(n815), .B(n606), .C(n52), .Y(n896) );
  OAI21X1 U280 ( .A(n819), .B(n605), .C(n457), .Y(n895) );
  OAI21X1 U282 ( .A(n818), .B(n605), .C(n455), .Y(n894) );
  OAI21X1 U284 ( .A(n817), .B(n605), .C(n453), .Y(n893) );
  OAI21X1 U286 ( .A(n816), .B(n605), .C(n451), .Y(n892) );
  OAI21X1 U288 ( .A(n815), .B(n605), .C(n50), .Y(n891) );
  OAI21X1 U292 ( .A(n819), .B(n602), .C(n449), .Y(n890) );
  OAI21X1 U294 ( .A(n818), .B(n602), .C(n287), .Y(n889) );
  OAI21X1 U296 ( .A(n817), .B(n602), .C(n284), .Y(n888) );
  OAI21X1 U298 ( .A(n816), .B(n602), .C(n48), .Y(n887) );
  OAI21X1 U300 ( .A(n815), .B(n602), .C(n46), .Y(n886) );
  OAI21X1 U304 ( .A(n819), .B(n601), .C(n282), .Y(n885) );
  OAI21X1 U306 ( .A(n818), .B(n601), .C(n280), .Y(n884) );
  OAI21X1 U308 ( .A(n817), .B(n601), .C(n278), .Y(n883) );
  OAI21X1 U310 ( .A(n816), .B(n601), .C(n276), .Y(n882) );
  OAI21X1 U312 ( .A(n815), .B(n601), .C(n44), .Y(n881) );
  OAI21X1 U316 ( .A(n819), .B(n599), .C(n274), .Y(n880) );
  OAI21X1 U318 ( .A(n818), .B(n599), .C(n272), .Y(n879) );
  OAI21X1 U320 ( .A(n817), .B(n599), .C(n270), .Y(n878) );
  OAI21X1 U322 ( .A(n816), .B(n599), .C(n42), .Y(n877) );
  OAI21X1 U324 ( .A(n815), .B(n599), .C(n40), .Y(n876) );
  OAI21X1 U328 ( .A(n819), .B(n597), .C(n268), .Y(n875) );
  OAI21X1 U330 ( .A(n818), .B(n597), .C(n266), .Y(n874) );
  OAI21X1 U332 ( .A(n817), .B(n597), .C(n264), .Y(n873) );
  OAI21X1 U334 ( .A(n816), .B(n597), .C(n38), .Y(n872) );
  OAI21X1 U336 ( .A(n815), .B(n597), .C(n36), .Y(n871) );
  NAND3X1 U340 ( .A(n994), .B(n826), .C(N13), .Y(n992) );
  OAI21X1 U341 ( .A(n819), .B(n594), .C(n34), .Y(n870) );
  OAI21X1 U343 ( .A(n818), .B(n594), .C(n32), .Y(n869) );
  OAI21X1 U345 ( .A(n817), .B(n594), .C(n30), .Y(n868) );
  OAI21X1 U347 ( .A(n816), .B(n594), .C(n28), .Y(n867) );
  OAI21X1 U349 ( .A(n815), .B(n594), .C(n26), .Y(n866) );
  NOR3X1 U353 ( .A(n823), .B(n644), .C(n825), .Y(n1003) );
  OAI21X1 U354 ( .A(n819), .B(n592), .C(n262), .Y(n865) );
  OAI21X1 U356 ( .A(n818), .B(n592), .C(n260), .Y(n864) );
  OAI21X1 U358 ( .A(n817), .B(n592), .C(n258), .Y(n863) );
  OAI21X1 U360 ( .A(n816), .B(n592), .C(n256), .Y(n862) );
  OAI21X1 U362 ( .A(n815), .B(n592), .C(n24), .Y(n861) );
  NOR3X1 U366 ( .A(n823), .B(n814), .C(n825), .Y(n1002) );
  OAI21X1 U367 ( .A(n819), .B(n591), .C(n22), .Y(n860) );
  OAI21X1 U369 ( .A(n818), .B(n591), .C(n20), .Y(n859) );
  OAI21X1 U371 ( .A(n817), .B(n591), .C(n18), .Y(n858) );
  OAI21X1 U373 ( .A(n816), .B(n591), .C(n16), .Y(n857) );
  OAI21X1 U375 ( .A(n815), .B(n591), .C(n14), .Y(n856) );
  NOR3X1 U379 ( .A(n644), .B(n805), .C(n825), .Y(n1001) );
  OAI21X1 U380 ( .A(n819), .B(n589), .C(n254), .Y(n855) );
  OAI21X1 U382 ( .A(n818), .B(n589), .C(n252), .Y(n854) );
  OAI21X1 U384 ( .A(n817), .B(n589), .C(n250), .Y(n853) );
  OAI21X1 U386 ( .A(n816), .B(n589), .C(n248), .Y(n852) );
  OAI21X1 U388 ( .A(n815), .B(n589), .C(n12), .Y(n851) );
  NOR3X1 U392 ( .A(n643), .B(n805), .C(n825), .Y(n1000) );
  OAI21X1 U393 ( .A(n819), .B(n587), .C(n246), .Y(n850) );
  OAI21X1 U395 ( .A(n818), .B(n587), .C(n244), .Y(n849) );
  OAI21X1 U397 ( .A(n817), .B(n587), .C(n242), .Y(n848) );
  OAI21X1 U399 ( .A(n816), .B(n587), .C(n240), .Y(n847) );
  OAI21X1 U401 ( .A(n815), .B(n587), .C(n10), .Y(n846) );
  NOR3X1 U405 ( .A(n644), .B(n824), .C(n823), .Y(n999) );
  OAI21X1 U406 ( .A(n819), .B(n585), .C(n238), .Y(n845) );
  OAI21X1 U408 ( .A(n818), .B(n585), .C(n236), .Y(n844) );
  OAI21X1 U410 ( .A(n817), .B(n585), .C(n234), .Y(n843) );
  OAI21X1 U412 ( .A(n816), .B(n585), .C(n232), .Y(n842) );
  OAI21X1 U414 ( .A(n815), .B(n585), .C(n8), .Y(n841) );
  NOR3X1 U418 ( .A(n812), .B(n824), .C(n823), .Y(n998) );
  OAI21X1 U419 ( .A(n819), .B(n583), .C(n230), .Y(n840) );
  OAI21X1 U421 ( .A(n818), .B(n583), .C(n227), .Y(n839) );
  OAI21X1 U423 ( .A(n817), .B(n583), .C(n225), .Y(n838) );
  OAI21X1 U425 ( .A(n816), .B(n583), .C(n223), .Y(n837) );
  OAI21X1 U427 ( .A(n815), .B(n583), .C(n6), .Y(n836) );
  NOR3X1 U431 ( .A(n805), .B(n824), .C(n644), .Y(n997) );
  OAI21X1 U432 ( .A(n819), .B(n581), .C(n221), .Y(n835) );
  OAI21X1 U435 ( .A(n818), .B(n581), .C(n219), .Y(n834) );
  OAI21X1 U438 ( .A(n817), .B(n581), .C(n217), .Y(n833) );
  OAI21X1 U441 ( .A(n816), .B(n581), .C(n215), .Y(n832) );
  OAI21X1 U444 ( .A(n815), .B(n581), .C(n4), .Y(n831) );
  NOR3X1 U448 ( .A(n805), .B(n824), .C(n645), .Y(n996) );
  NAND3X1 U449 ( .A(n646), .B(n826), .C(n994), .Y(n991) );
  NOR3X1 U450 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n994) );
  INVX2 U3 ( .A(n513), .Y(n819) );
  INVX2 U4 ( .A(n512), .Y(n818) );
  INVX2 U5 ( .A(n511), .Y(n817) );
  INVX2 U6 ( .A(n510), .Y(n816) );
  INVX2 U7 ( .A(n509), .Y(n815) );
  AND2X1 U8 ( .A(\mem<31><0> ), .B(n577), .Y(n211) );
  AND2X1 U9 ( .A(\mem<31><1> ), .B(n577), .Y(n209) );
  AND2X1 U10 ( .A(\mem<31><2> ), .B(n577), .Y(n207) );
  AND2X1 U11 ( .A(\mem<31><4> ), .B(n577), .Y(n203) );
  AND2X1 U12 ( .A(\mem<30><1> ), .B(n575), .Y(n199) );
  AND2X1 U13 ( .A(\mem<30><4> ), .B(n575), .Y(n193) );
  AND2X1 U14 ( .A(\mem<29><0> ), .B(n573), .Y(n191) );
  AND2X1 U15 ( .A(\mem<29><1> ), .B(n573), .Y(n189) );
  AND2X1 U16 ( .A(\mem<29><2> ), .B(n573), .Y(n187) );
  AND2X1 U17 ( .A(\mem<29><4> ), .B(n573), .Y(n183) );
  AND2X1 U18 ( .A(\mem<28><1> ), .B(n571), .Y(n179) );
  AND2X1 U19 ( .A(\mem<28><4> ), .B(n571), .Y(n173) );
  AND2X1 U20 ( .A(\mem<27><1> ), .B(n569), .Y(n168) );
  AND2X1 U21 ( .A(\mem<27><4> ), .B(n569), .Y(n162) );
  AND2X1 U22 ( .A(\mem<26><4> ), .B(n567), .Y(n160) );
  AND2X1 U23 ( .A(\mem<25><1> ), .B(n565), .Y(n156) );
  AND2X1 U24 ( .A(\mem<25><4> ), .B(n565), .Y(n150) );
  AND2X1 U25 ( .A(\mem<24><4> ), .B(n563), .Y(n148) );
  AND2X1 U26 ( .A(\mem<23><0> ), .B(n561), .Y(n146) );
  AND2X1 U27 ( .A(\mem<23><1> ), .B(n561), .Y(n144) );
  AND2X1 U28 ( .A(\mem<23><2> ), .B(n561), .Y(n142) );
  AND2X1 U29 ( .A(\mem<23><4> ), .B(n561), .Y(n138) );
  AND2X1 U30 ( .A(\mem<22><1> ), .B(n559), .Y(n134) );
  AND2X1 U31 ( .A(\mem<22><4> ), .B(n559), .Y(n128) );
  AND2X1 U32 ( .A(\mem<21><0> ), .B(n557), .Y(n126) );
  AND2X1 U33 ( .A(\mem<21><1> ), .B(n557), .Y(n124) );
  AND2X1 U34 ( .A(\mem<21><2> ), .B(n557), .Y(n122) );
  AND2X1 U35 ( .A(\mem<21><4> ), .B(n557), .Y(n118) );
  AND2X1 U36 ( .A(\mem<20><1> ), .B(n555), .Y(n111) );
  AND2X1 U37 ( .A(\mem<20><4> ), .B(n555), .Y(n104) );
  AND2X1 U38 ( .A(\mem<19><1> ), .B(n553), .Y(n100) );
  AND2X1 U39 ( .A(\mem<19><4> ), .B(n553), .Y(n93) );
  AND2X1 U40 ( .A(\mem<18><4> ), .B(n551), .Y(n91) );
  AND2X1 U41 ( .A(\mem<17><1> ), .B(n549), .Y(n86) );
  AND2X1 U42 ( .A(\mem<17><4> ), .B(n549), .Y(n79) );
  AND2X1 U43 ( .A(\mem<16><4> ), .B(n547), .Y(n77) );
  AND2X1 U44 ( .A(\mem<15><1> ), .B(n545), .Y(n72) );
  AND2X1 U45 ( .A(\mem<15><4> ), .B(n545), .Y(n70) );
  AND2X1 U46 ( .A(\mem<14><4> ), .B(n543), .Y(n63) );
  AND2X1 U47 ( .A(\mem<13><1> ), .B(n541), .Y(n59) );
  AND2X1 U48 ( .A(\mem<13><4> ), .B(n541), .Y(n51) );
  AND2X1 U49 ( .A(\mem<12><4> ), .B(n539), .Y(n49) );
  AND2X1 U51 ( .A(\mem<11><4> ), .B(n537), .Y(n45) );
  AND2X1 U53 ( .A(\mem<10><4> ), .B(n535), .Y(n43) );
  AND2X1 U55 ( .A(\mem<9><4> ), .B(n533), .Y(n39) );
  AND2X1 U57 ( .A(\mem<8><4> ), .B(n531), .Y(n35) );
  AND2X1 U59 ( .A(\mem<7><1> ), .B(n529), .Y(n31) );
  AND2X1 U60 ( .A(\mem<7><4> ), .B(n529), .Y(n25) );
  AND2X1 U61 ( .A(\mem<6><4> ), .B(n527), .Y(n23) );
  AND2X1 U63 ( .A(\mem<5><1> ), .B(n525), .Y(n19) );
  AND2X1 U65 ( .A(\mem<5><4> ), .B(n525), .Y(n13) );
  AND2X1 U67 ( .A(\mem<4><4> ), .B(n523), .Y(n11) );
  AND2X1 U69 ( .A(\mem<3><4> ), .B(n521), .Y(n9) );
  AND2X1 U71 ( .A(\mem<2><4> ), .B(n519), .Y(n7) );
  AND2X1 U72 ( .A(\mem<1><4> ), .B(n517), .Y(n5) );
  AND2X1 U73 ( .A(\mem<0><4> ), .B(n515), .Y(n3) );
  INVX1 U75 ( .A(N14), .Y(n826) );
  INVX2 U77 ( .A(N13), .Y(n646) );
  INVX1 U79 ( .A(rst), .Y(n820) );
  INVX8 U81 ( .A(n825), .Y(n802) );
  INVX4 U83 ( .A(n821), .Y(n809) );
  INVX1 U84 ( .A(n825), .Y(n824) );
  OR2X2 U85 ( .A(write), .B(rst), .Y(n1) );
  INVX1 U87 ( .A(n1), .Y(n2) );
  INVX1 U89 ( .A(n3), .Y(n4) );
  INVX1 U91 ( .A(n5), .Y(n6) );
  INVX1 U93 ( .A(n7), .Y(n8) );
  INVX1 U95 ( .A(n9), .Y(n10) );
  INVX1 U96 ( .A(n11), .Y(n12) );
  INVX1 U97 ( .A(n13), .Y(n14) );
  AND2X2 U99 ( .A(\mem<5><3> ), .B(n525), .Y(n15) );
  INVX1 U101 ( .A(n15), .Y(n16) );
  AND2X2 U103 ( .A(\mem<5><2> ), .B(n525), .Y(n17) );
  INVX1 U105 ( .A(n17), .Y(n18) );
  INVX1 U107 ( .A(n19), .Y(n20) );
  AND2X2 U108 ( .A(\mem<5><0> ), .B(n525), .Y(n21) );
  INVX1 U109 ( .A(n21), .Y(n22) );
  INVX1 U111 ( .A(n23), .Y(n24) );
  INVX1 U113 ( .A(n25), .Y(n26) );
  AND2X2 U115 ( .A(\mem<7><3> ), .B(n529), .Y(n27) );
  INVX1 U117 ( .A(n27), .Y(n28) );
  AND2X2 U119 ( .A(\mem<7><2> ), .B(n529), .Y(n29) );
  INVX1 U120 ( .A(n29), .Y(n30) );
  INVX1 U121 ( .A(n31), .Y(n32) );
  AND2X2 U123 ( .A(\mem<7><0> ), .B(n529), .Y(n33) );
  INVX1 U125 ( .A(n33), .Y(n34) );
  INVX1 U127 ( .A(n35), .Y(n36) );
  AND2X2 U129 ( .A(\mem<8><3> ), .B(n531), .Y(n37) );
  INVX1 U131 ( .A(n37), .Y(n38) );
  INVX1 U132 ( .A(n39), .Y(n40) );
  AND2X2 U133 ( .A(\mem<9><3> ), .B(n533), .Y(n41) );
  INVX1 U135 ( .A(n41), .Y(n42) );
  INVX1 U137 ( .A(n43), .Y(n44) );
  INVX1 U139 ( .A(n45), .Y(n46) );
  AND2X2 U141 ( .A(\mem<11><3> ), .B(n537), .Y(n47) );
  INVX1 U143 ( .A(n47), .Y(n48) );
  INVX1 U144 ( .A(n49), .Y(n50) );
  INVX1 U145 ( .A(n51), .Y(n52) );
  AND2X2 U148 ( .A(\mem<13><3> ), .B(n541), .Y(n53) );
  INVX1 U150 ( .A(n53), .Y(n54) );
  AND2X2 U152 ( .A(\mem<13><2> ), .B(n541), .Y(n55) );
  INVX1 U154 ( .A(n55), .Y(n58) );
  INVX1 U156 ( .A(n59), .Y(n60) );
  AND2X2 U157 ( .A(\mem<13><0> ), .B(n541), .Y(n61) );
  INVX1 U158 ( .A(n61), .Y(n62) );
  INVX1 U160 ( .A(n63), .Y(n64) );
  AND2X2 U162 ( .A(\mem<14><3> ), .B(n543), .Y(n66) );
  INVX1 U164 ( .A(n66), .Y(n67) );
  AND2X2 U166 ( .A(\mem<14><2> ), .B(n543), .Y(n68) );
  INVX1 U168 ( .A(n68), .Y(n69) );
  INVX1 U169 ( .A(n70), .Y(n71) );
  INVX1 U170 ( .A(n72), .Y(n74) );
  AND2X2 U172 ( .A(\mem<15><0> ), .B(n545), .Y(n75) );
  INVX1 U174 ( .A(n75), .Y(n76) );
  INVX1 U176 ( .A(n77), .Y(n78) );
  INVX1 U178 ( .A(n79), .Y(n80) );
  AND2X2 U180 ( .A(\mem<17><3> ), .B(n549), .Y(n82) );
  INVX1 U181 ( .A(n82), .Y(n83) );
  AND2X2 U182 ( .A(\mem<17><2> ), .B(n549), .Y(n84) );
  INVX1 U184 ( .A(n84), .Y(n85) );
  INVX1 U186 ( .A(n86), .Y(n87) );
  AND2X2 U188 ( .A(\mem<17><0> ), .B(n549), .Y(n88) );
  INVX1 U190 ( .A(n88), .Y(n90) );
  INVX1 U192 ( .A(n91), .Y(n92) );
  INVX1 U193 ( .A(n93), .Y(n94) );
  AND2X2 U194 ( .A(\mem<19><3> ), .B(n553), .Y(n95) );
  INVX1 U196 ( .A(n95), .Y(n96) );
  AND2X2 U198 ( .A(\mem<19><2> ), .B(n553), .Y(n98) );
  INVX1 U200 ( .A(n98), .Y(n99) );
  INVX1 U202 ( .A(n100), .Y(n101) );
  AND2X2 U204 ( .A(\mem<19><0> ), .B(n553), .Y(n102) );
  INVX1 U205 ( .A(n102), .Y(n103) );
  INVX1 U206 ( .A(n104), .Y(n106) );
  AND2X2 U208 ( .A(\mem<20><3> ), .B(n555), .Y(n107) );
  INVX1 U210 ( .A(n107), .Y(n108) );
  AND2X2 U212 ( .A(\mem<20><2> ), .B(n555), .Y(n109) );
  INVX1 U214 ( .A(n109), .Y(n110) );
  INVX1 U216 ( .A(n111), .Y(n112) );
  AND2X2 U217 ( .A(\mem<20><0> ), .B(n555), .Y(n116) );
  INVX1 U218 ( .A(n116), .Y(n117) );
  INVX1 U220 ( .A(n118), .Y(n119) );
  AND2X2 U222 ( .A(\mem<21><3> ), .B(n557), .Y(n120) );
  INVX1 U224 ( .A(n120), .Y(n121) );
  INVX1 U226 ( .A(n122), .Y(n123) );
  INVX1 U228 ( .A(n124), .Y(n125) );
  INVX1 U229 ( .A(n126), .Y(n127) );
  INVX1 U230 ( .A(n128), .Y(n129) );
  AND2X2 U232 ( .A(\mem<22><3> ), .B(n559), .Y(n130) );
  INVX1 U234 ( .A(n130), .Y(n131) );
  AND2X2 U236 ( .A(\mem<22><2> ), .B(n559), .Y(n132) );
  INVX1 U238 ( .A(n132), .Y(n133) );
  INVX1 U240 ( .A(n134), .Y(n135) );
  AND2X2 U241 ( .A(\mem<22><0> ), .B(n559), .Y(n136) );
  INVX1 U242 ( .A(n136), .Y(n137) );
  INVX1 U245 ( .A(n138), .Y(n139) );
  AND2X2 U247 ( .A(\mem<23><3> ), .B(n561), .Y(n140) );
  INVX1 U249 ( .A(n140), .Y(n141) );
  INVX1 U251 ( .A(n142), .Y(n143) );
  INVX1 U253 ( .A(n144), .Y(n145) );
  INVX1 U254 ( .A(n146), .Y(n147) );
  INVX1 U255 ( .A(n148), .Y(n149) );
  INVX1 U257 ( .A(n150), .Y(n151) );
  AND2X2 U259 ( .A(\mem<25><3> ), .B(n565), .Y(n152) );
  INVX1 U261 ( .A(n152), .Y(n153) );
  AND2X2 U263 ( .A(\mem<25><2> ), .B(n565), .Y(n154) );
  INVX1 U265 ( .A(n154), .Y(n155) );
  INVX1 U266 ( .A(n156), .Y(n157) );
  AND2X2 U267 ( .A(\mem<25><0> ), .B(n565), .Y(n158) );
  INVX1 U269 ( .A(n158), .Y(n159) );
  INVX1 U271 ( .A(n160), .Y(n161) );
  INVX1 U273 ( .A(n162), .Y(n163) );
  AND2X2 U275 ( .A(\mem<27><3> ), .B(n569), .Y(n164) );
  INVX1 U277 ( .A(n164), .Y(n165) );
  AND2X2 U278 ( .A(\mem<27><2> ), .B(n569), .Y(n166) );
  INVX1 U279 ( .A(n166), .Y(n167) );
  INVX1 U281 ( .A(n168), .Y(n169) );
  AND2X2 U283 ( .A(\mem<27><0> ), .B(n569), .Y(n170) );
  INVX1 U285 ( .A(n170), .Y(n171) );
  INVX1 U287 ( .A(n173), .Y(n174) );
  AND2X2 U289 ( .A(\mem<28><3> ), .B(n571), .Y(n175) );
  INVX1 U290 ( .A(n175), .Y(n176) );
  AND2X2 U291 ( .A(\mem<28><2> ), .B(n571), .Y(n177) );
  INVX1 U293 ( .A(n177), .Y(n178) );
  INVX1 U295 ( .A(n179), .Y(n180) );
  AND2X2 U297 ( .A(\mem<28><0> ), .B(n571), .Y(n181) );
  INVX1 U299 ( .A(n181), .Y(n182) );
  INVX1 U301 ( .A(n183), .Y(n184) );
  AND2X2 U302 ( .A(\mem<29><3> ), .B(n573), .Y(n185) );
  INVX1 U303 ( .A(n185), .Y(n186) );
  INVX1 U305 ( .A(n187), .Y(n188) );
  INVX1 U307 ( .A(n189), .Y(n190) );
  INVX1 U309 ( .A(n191), .Y(n192) );
  INVX1 U311 ( .A(n193), .Y(n194) );
  AND2X2 U313 ( .A(\mem<30><3> ), .B(n575), .Y(n195) );
  INVX1 U314 ( .A(n195), .Y(n196) );
  AND2X2 U315 ( .A(\mem<30><2> ), .B(n575), .Y(n197) );
  INVX1 U317 ( .A(n197), .Y(n198) );
  INVX1 U319 ( .A(n199), .Y(n200) );
  AND2X2 U321 ( .A(\mem<30><0> ), .B(n575), .Y(n201) );
  INVX1 U323 ( .A(n201), .Y(n202) );
  INVX1 U325 ( .A(n203), .Y(n204) );
  AND2X2 U326 ( .A(\mem<31><3> ), .B(n577), .Y(n205) );
  INVX1 U327 ( .A(n205), .Y(n206) );
  INVX1 U329 ( .A(n207), .Y(n208) );
  INVX1 U331 ( .A(n209), .Y(n210) );
  INVX1 U333 ( .A(n211), .Y(n212) );
  AND2X2 U335 ( .A(n501), .B(n499), .Y(n213) );
  AND2X2 U337 ( .A(\mem<0><3> ), .B(n515), .Y(n214) );
  INVX1 U338 ( .A(n214), .Y(n215) );
  AND2X2 U339 ( .A(\mem<0><2> ), .B(n515), .Y(n216) );
  INVX1 U342 ( .A(n216), .Y(n217) );
  AND2X2 U344 ( .A(\mem<0><1> ), .B(n515), .Y(n218) );
  INVX1 U346 ( .A(n218), .Y(n219) );
  AND2X2 U348 ( .A(\mem<0><0> ), .B(n515), .Y(n220) );
  INVX1 U350 ( .A(n220), .Y(n221) );
  AND2X2 U351 ( .A(\mem<1><3> ), .B(n517), .Y(n222) );
  INVX1 U352 ( .A(n222), .Y(n223) );
  AND2X2 U355 ( .A(\mem<1><2> ), .B(n517), .Y(n224) );
  INVX1 U357 ( .A(n224), .Y(n225) );
  AND2X2 U359 ( .A(\mem<1><1> ), .B(n517), .Y(n226) );
  INVX1 U361 ( .A(n226), .Y(n227) );
  AND2X2 U363 ( .A(\mem<1><0> ), .B(n517), .Y(n228) );
  INVX1 U364 ( .A(n228), .Y(n230) );
  AND2X2 U365 ( .A(\mem<2><3> ), .B(n519), .Y(n231) );
  INVX1 U368 ( .A(n231), .Y(n232) );
  AND2X2 U370 ( .A(\mem<2><2> ), .B(n519), .Y(n233) );
  INVX1 U372 ( .A(n233), .Y(n234) );
  AND2X2 U374 ( .A(\mem<2><1> ), .B(n519), .Y(n235) );
  INVX1 U376 ( .A(n235), .Y(n236) );
  AND2X2 U377 ( .A(\mem<2><0> ), .B(n519), .Y(n237) );
  INVX1 U378 ( .A(n237), .Y(n238) );
  AND2X2 U381 ( .A(\mem<3><3> ), .B(n521), .Y(n239) );
  INVX1 U383 ( .A(n239), .Y(n240) );
  AND2X2 U385 ( .A(\mem<3><2> ), .B(n521), .Y(n241) );
  INVX1 U387 ( .A(n241), .Y(n242) );
  AND2X2 U389 ( .A(\mem<3><1> ), .B(n521), .Y(n243) );
  INVX1 U390 ( .A(n243), .Y(n244) );
  AND2X2 U391 ( .A(\mem<3><0> ), .B(n521), .Y(n245) );
  INVX1 U394 ( .A(n245), .Y(n246) );
  AND2X2 U396 ( .A(\mem<4><3> ), .B(n523), .Y(n247) );
  INVX1 U398 ( .A(n247), .Y(n248) );
  AND2X2 U400 ( .A(\mem<4><2> ), .B(n523), .Y(n249) );
  INVX1 U402 ( .A(n249), .Y(n250) );
  AND2X2 U403 ( .A(\mem<4><1> ), .B(n523), .Y(n251) );
  INVX1 U404 ( .A(n251), .Y(n252) );
  AND2X2 U407 ( .A(\mem<4><0> ), .B(n523), .Y(n253) );
  INVX1 U409 ( .A(n253), .Y(n254) );
  AND2X2 U411 ( .A(\mem<6><3> ), .B(n527), .Y(n255) );
  INVX1 U413 ( .A(n255), .Y(n256) );
  AND2X2 U415 ( .A(\mem<6><2> ), .B(n527), .Y(n257) );
  INVX1 U416 ( .A(n257), .Y(n258) );
  AND2X2 U417 ( .A(\mem<6><1> ), .B(n527), .Y(n259) );
  INVX1 U420 ( .A(n259), .Y(n260) );
  AND2X2 U422 ( .A(\mem<6><0> ), .B(n527), .Y(n261) );
  INVX1 U424 ( .A(n261), .Y(n262) );
  AND2X2 U426 ( .A(\mem<8><2> ), .B(n531), .Y(n263) );
  INVX1 U428 ( .A(n263), .Y(n264) );
  AND2X2 U429 ( .A(\mem<8><1> ), .B(n531), .Y(n265) );
  INVX1 U430 ( .A(n265), .Y(n266) );
  AND2X2 U433 ( .A(\mem<8><0> ), .B(n531), .Y(n267) );
  INVX1 U434 ( .A(n267), .Y(n268) );
  AND2X2 U436 ( .A(\mem<9><2> ), .B(n533), .Y(n269) );
  INVX1 U437 ( .A(n269), .Y(n270) );
  AND2X2 U439 ( .A(\mem<9><1> ), .B(n533), .Y(n271) );
  INVX1 U440 ( .A(n271), .Y(n272) );
  AND2X2 U442 ( .A(\mem<9><0> ), .B(n533), .Y(n273) );
  INVX1 U443 ( .A(n273), .Y(n274) );
  AND2X2 U445 ( .A(\mem<10><3> ), .B(n535), .Y(n275) );
  INVX1 U446 ( .A(n275), .Y(n276) );
  AND2X2 U447 ( .A(\mem<10><2> ), .B(n535), .Y(n277) );
  INVX1 U451 ( .A(n277), .Y(n278) );
  AND2X2 U452 ( .A(\mem<10><1> ), .B(n535), .Y(n279) );
  INVX1 U453 ( .A(n279), .Y(n280) );
  AND2X2 U454 ( .A(\mem<10><0> ), .B(n535), .Y(n281) );
  INVX1 U455 ( .A(n281), .Y(n282) );
  AND2X2 U456 ( .A(\mem<11><2> ), .B(n537), .Y(n283) );
  INVX1 U457 ( .A(n283), .Y(n284) );
  AND2X2 U458 ( .A(\mem<11><1> ), .B(n537), .Y(n285) );
  INVX1 U459 ( .A(n285), .Y(n287) );
  AND2X2 U460 ( .A(\mem<11><0> ), .B(n537), .Y(n448) );
  INVX1 U461 ( .A(n448), .Y(n449) );
  AND2X2 U462 ( .A(\mem<12><3> ), .B(n539), .Y(n450) );
  INVX1 U463 ( .A(n450), .Y(n451) );
  AND2X2 U464 ( .A(\mem<12><2> ), .B(n539), .Y(n452) );
  INVX1 U465 ( .A(n452), .Y(n453) );
  AND2X2 U466 ( .A(\mem<12><1> ), .B(n539), .Y(n454) );
  INVX1 U467 ( .A(n454), .Y(n455) );
  AND2X2 U468 ( .A(\mem<12><0> ), .B(n539), .Y(n456) );
  INVX1 U469 ( .A(n456), .Y(n457) );
  AND2X2 U470 ( .A(\mem<14><1> ), .B(n543), .Y(n458) );
  INVX1 U471 ( .A(n458), .Y(n459) );
  AND2X2 U472 ( .A(\mem<14><0> ), .B(n543), .Y(n460) );
  INVX1 U473 ( .A(n460), .Y(n461) );
  AND2X2 U474 ( .A(\mem<15><3> ), .B(n545), .Y(n462) );
  INVX1 U475 ( .A(n462), .Y(n463) );
  AND2X2 U476 ( .A(\mem<15><2> ), .B(n545), .Y(n464) );
  INVX1 U477 ( .A(n464), .Y(n465) );
  AND2X2 U478 ( .A(\mem<16><3> ), .B(n547), .Y(n466) );
  INVX1 U479 ( .A(n466), .Y(n467) );
  AND2X2 U480 ( .A(\mem<16><2> ), .B(n547), .Y(n468) );
  INVX1 U481 ( .A(n468), .Y(n469) );
  AND2X2 U482 ( .A(\mem<16><1> ), .B(n547), .Y(n470) );
  INVX1 U483 ( .A(n470), .Y(n471) );
  AND2X2 U484 ( .A(\mem<16><0> ), .B(n547), .Y(n472) );
  INVX1 U485 ( .A(n472), .Y(n473) );
  AND2X2 U486 ( .A(\mem<18><3> ), .B(n551), .Y(n474) );
  INVX1 U487 ( .A(n474), .Y(n475) );
  AND2X2 U488 ( .A(\mem<18><2> ), .B(n551), .Y(n476) );
  INVX1 U489 ( .A(n476), .Y(n477) );
  AND2X2 U490 ( .A(\mem<18><1> ), .B(n551), .Y(n478) );
  INVX1 U491 ( .A(n478), .Y(n479) );
  AND2X2 U492 ( .A(\mem<18><0> ), .B(n551), .Y(n480) );
  INVX1 U493 ( .A(n480), .Y(n481) );
  AND2X2 U494 ( .A(\mem<24><3> ), .B(n563), .Y(n482) );
  INVX1 U495 ( .A(n482), .Y(n483) );
  AND2X2 U496 ( .A(\mem<24><2> ), .B(n563), .Y(n484) );
  INVX1 U497 ( .A(n484), .Y(n485) );
  AND2X2 U498 ( .A(\mem<24><1> ), .B(n563), .Y(n486) );
  INVX1 U499 ( .A(n486), .Y(n487) );
  AND2X2 U500 ( .A(\mem<24><0> ), .B(n563), .Y(n488) );
  INVX1 U501 ( .A(n488), .Y(n489) );
  AND2X2 U502 ( .A(\mem<26><3> ), .B(n567), .Y(n490) );
  INVX1 U503 ( .A(n490), .Y(n491) );
  AND2X2 U504 ( .A(\mem<26><2> ), .B(n567), .Y(n492) );
  INVX1 U505 ( .A(n492), .Y(n493) );
  AND2X2 U506 ( .A(\mem<26><1> ), .B(n567), .Y(n494) );
  INVX1 U507 ( .A(n494), .Y(n495) );
  AND2X2 U508 ( .A(\mem<26><0> ), .B(n567), .Y(n496) );
  INVX1 U509 ( .A(n496), .Y(n497) );
  AND2X2 U510 ( .A(n753), .B(n802), .Y(n498) );
  INVX1 U511 ( .A(n498), .Y(n499) );
  AND2X2 U512 ( .A(n756), .B(n825), .Y(n500) );
  INVX1 U513 ( .A(n500), .Y(n501) );
  OR2X2 U514 ( .A(write), .B(rst), .Y(n502) );
  INVX1 U515 ( .A(n1), .Y(n503) );
  INVX1 U516 ( .A(n502), .Y(n504) );
  BUFX2 U517 ( .A(n991), .Y(n505) );
  INVX1 U518 ( .A(n505), .Y(n827) );
  BUFX2 U519 ( .A(n992), .Y(n506) );
  INVX1 U520 ( .A(n506), .Y(n828) );
  BUFX2 U521 ( .A(n993), .Y(n507) );
  INVX1 U522 ( .A(n507), .Y(n829) );
  BUFX2 U523 ( .A(n995), .Y(n508) );
  INVX1 U524 ( .A(n508), .Y(n830) );
  AND2X1 U525 ( .A(\data_in<4> ), .B(n1004), .Y(n509) );
  AND2X1 U526 ( .A(\data_in<3> ), .B(n1004), .Y(n510) );
  AND2X1 U527 ( .A(\data_in<2> ), .B(n1004), .Y(n511) );
  AND2X1 U528 ( .A(\data_in<1> ), .B(n1004), .Y(n512) );
  AND2X1 U529 ( .A(\data_in<0> ), .B(n1004), .Y(n513) );
  AND2X1 U530 ( .A(n580), .B(n1004), .Y(n514) );
  INVX1 U531 ( .A(n514), .Y(n515) );
  AND2X1 U532 ( .A(n582), .B(n1004), .Y(n516) );
  INVX1 U533 ( .A(n516), .Y(n517) );
  AND2X1 U534 ( .A(n584), .B(n1004), .Y(n518) );
  INVX1 U535 ( .A(n518), .Y(n519) );
  AND2X1 U536 ( .A(n586), .B(n1004), .Y(n520) );
  INVX1 U537 ( .A(n520), .Y(n521) );
  AND2X1 U538 ( .A(n588), .B(n1004), .Y(n522) );
  INVX1 U539 ( .A(n522), .Y(n523) );
  AND2X1 U540 ( .A(n590), .B(n1004), .Y(n524) );
  INVX1 U541 ( .A(n524), .Y(n525) );
  AND2X1 U542 ( .A(n593), .B(n1004), .Y(n526) );
  INVX1 U543 ( .A(n526), .Y(n527) );
  AND2X1 U544 ( .A(n595), .B(n1004), .Y(n528) );
  INVX1 U545 ( .A(n528), .Y(n529) );
  AND2X1 U546 ( .A(n596), .B(n1004), .Y(n530) );
  INVX1 U547 ( .A(n530), .Y(n531) );
  AND2X1 U548 ( .A(n598), .B(n1004), .Y(n532) );
  INVX1 U549 ( .A(n532), .Y(n533) );
  AND2X1 U550 ( .A(n600), .B(n1004), .Y(n534) );
  INVX1 U551 ( .A(n534), .Y(n535) );
  AND2X1 U552 ( .A(n603), .B(n1004), .Y(n536) );
  INVX1 U553 ( .A(n536), .Y(n537) );
  AND2X1 U554 ( .A(n604), .B(n1004), .Y(n538) );
  INVX1 U555 ( .A(n538), .Y(n539) );
  AND2X1 U556 ( .A(n607), .B(n1004), .Y(n540) );
  INVX1 U557 ( .A(n540), .Y(n541) );
  AND2X1 U558 ( .A(n609), .B(n1004), .Y(n542) );
  INVX1 U559 ( .A(n542), .Y(n543) );
  AND2X1 U560 ( .A(n611), .B(n1004), .Y(n544) );
  INVX1 U561 ( .A(n544), .Y(n545) );
  AND2X1 U562 ( .A(n612), .B(n1004), .Y(n546) );
  INVX1 U563 ( .A(n546), .Y(n547) );
  AND2X1 U564 ( .A(n614), .B(n1004), .Y(n548) );
  INVX1 U565 ( .A(n548), .Y(n549) );
  AND2X1 U566 ( .A(n616), .B(n1004), .Y(n550) );
  INVX1 U567 ( .A(n550), .Y(n551) );
  AND2X1 U568 ( .A(n619), .B(n1004), .Y(n552) );
  INVX1 U569 ( .A(n552), .Y(n553) );
  AND2X1 U570 ( .A(n620), .B(n1004), .Y(n554) );
  INVX1 U571 ( .A(n554), .Y(n555) );
  AND2X1 U572 ( .A(n623), .B(n1004), .Y(n556) );
  INVX1 U573 ( .A(n556), .Y(n557) );
  AND2X1 U574 ( .A(n625), .B(n1004), .Y(n558) );
  INVX1 U575 ( .A(n558), .Y(n559) );
  AND2X1 U576 ( .A(n627), .B(n1004), .Y(n560) );
  INVX1 U577 ( .A(n560), .Y(n561) );
  AND2X1 U578 ( .A(n628), .B(n1004), .Y(n562) );
  INVX1 U579 ( .A(n562), .Y(n563) );
  AND2X1 U580 ( .A(n630), .B(n1004), .Y(n564) );
  INVX1 U581 ( .A(n564), .Y(n565) );
  AND2X1 U582 ( .A(n632), .B(n1004), .Y(n566) );
  INVX1 U583 ( .A(n566), .Y(n567) );
  AND2X1 U584 ( .A(n634), .B(n1004), .Y(n568) );
  INVX1 U585 ( .A(n568), .Y(n569) );
  AND2X1 U586 ( .A(n636), .B(n1004), .Y(n570) );
  INVX1 U587 ( .A(n570), .Y(n571) );
  AND2X1 U588 ( .A(n638), .B(n1004), .Y(n572) );
  INVX1 U589 ( .A(n572), .Y(n573) );
  AND2X1 U590 ( .A(n640), .B(n1004), .Y(n574) );
  INVX1 U591 ( .A(n574), .Y(n575) );
  AND2X1 U592 ( .A(n579), .B(n1004), .Y(n576) );
  INVX1 U593 ( .A(n576), .Y(n577) );
  INVX1 U594 ( .A(n579), .Y(n578) );
  AND2X1 U595 ( .A(n1003), .B(n830), .Y(n579) );
  AND2X1 U596 ( .A(n827), .B(n996), .Y(n580) );
  INVX1 U597 ( .A(n580), .Y(n581) );
  AND2X1 U598 ( .A(n827), .B(n997), .Y(n582) );
  INVX1 U599 ( .A(n582), .Y(n583) );
  AND2X1 U600 ( .A(n827), .B(n998), .Y(n584) );
  INVX1 U601 ( .A(n584), .Y(n585) );
  AND2X1 U602 ( .A(n827), .B(n999), .Y(n586) );
  INVX1 U603 ( .A(n586), .Y(n587) );
  AND2X1 U604 ( .A(n827), .B(n1000), .Y(n588) );
  INVX1 U605 ( .A(n588), .Y(n589) );
  AND2X1 U606 ( .A(n827), .B(n1001), .Y(n590) );
  INVX1 U607 ( .A(n590), .Y(n591) );
  INVX1 U608 ( .A(n593), .Y(n592) );
  AND2X1 U609 ( .A(n827), .B(n1002), .Y(n593) );
  INVX1 U610 ( .A(n595), .Y(n594) );
  AND2X1 U611 ( .A(n827), .B(n1003), .Y(n595) );
  AND2X1 U612 ( .A(n828), .B(n996), .Y(n596) );
  INVX1 U613 ( .A(n596), .Y(n597) );
  AND2X1 U614 ( .A(n828), .B(n997), .Y(n598) );
  INVX1 U615 ( .A(n598), .Y(n599) );
  AND2X1 U616 ( .A(n828), .B(n998), .Y(n600) );
  INVX1 U617 ( .A(n600), .Y(n601) );
  INVX1 U618 ( .A(n603), .Y(n602) );
  AND2X1 U619 ( .A(n828), .B(n999), .Y(n603) );
  AND2X1 U620 ( .A(n828), .B(n1000), .Y(n604) );
  INVX1 U621 ( .A(n604), .Y(n605) );
  INVX1 U622 ( .A(n607), .Y(n606) );
  AND2X1 U623 ( .A(n828), .B(n1001), .Y(n607) );
  INVX1 U624 ( .A(n609), .Y(n608) );
  AND2X1 U625 ( .A(n828), .B(n1002), .Y(n609) );
  INVX1 U626 ( .A(n611), .Y(n610) );
  AND2X1 U627 ( .A(n828), .B(n1003), .Y(n611) );
  AND2X1 U628 ( .A(n829), .B(n996), .Y(n612) );
  INVX1 U629 ( .A(n612), .Y(n613) );
  AND2X1 U630 ( .A(n829), .B(n997), .Y(n614) );
  INVX1 U631 ( .A(n614), .Y(n615) );
  AND2X1 U632 ( .A(n829), .B(n998), .Y(n616) );
  INVX1 U633 ( .A(n616), .Y(n617) );
  INVX1 U634 ( .A(n619), .Y(n618) );
  AND2X1 U635 ( .A(n829), .B(n999), .Y(n619) );
  AND2X1 U636 ( .A(n829), .B(n1000), .Y(n620) );
  INVX1 U637 ( .A(n620), .Y(n621) );
  INVX1 U638 ( .A(n623), .Y(n622) );
  AND2X1 U639 ( .A(n829), .B(n1001), .Y(n623) );
  INVX1 U640 ( .A(n625), .Y(n624) );
  AND2X1 U641 ( .A(n829), .B(n1002), .Y(n625) );
  INVX1 U642 ( .A(n627), .Y(n626) );
  AND2X1 U643 ( .A(n829), .B(n1003), .Y(n627) );
  AND2X1 U644 ( .A(n996), .B(n830), .Y(n628) );
  INVX1 U645 ( .A(n628), .Y(n629) );
  AND2X1 U646 ( .A(n997), .B(n830), .Y(n630) );
  INVX1 U647 ( .A(n630), .Y(n631) );
  AND2X1 U648 ( .A(n998), .B(n830), .Y(n632) );
  INVX1 U649 ( .A(n632), .Y(n633) );
  AND2X1 U650 ( .A(n999), .B(n830), .Y(n634) );
  INVX1 U651 ( .A(n634), .Y(n635) );
  AND2X1 U652 ( .A(n1000), .B(n830), .Y(n636) );
  INVX1 U653 ( .A(n636), .Y(n637) );
  AND2X1 U654 ( .A(n1001), .B(n830), .Y(n638) );
  INVX1 U655 ( .A(n638), .Y(n639) );
  AND2X1 U656 ( .A(n1002), .B(n830), .Y(n640) );
  INVX1 U657 ( .A(n640), .Y(n641) );
  BUFX4 U658 ( .A(n822), .Y(n642) );
  INVX1 U659 ( .A(N10), .Y(n822) );
  INVX1 U660 ( .A(n822), .Y(n821) );
  MUX2X1 U661 ( .B(n674), .A(n673), .S(n804), .Y(n672) );
  MUX2X1 U662 ( .B(\mem<15><3> ), .A(\mem<14><3> ), .S(n809), .Y(n755) );
  INVX1 U663 ( .A(n801), .Y(N17) );
  MUX2X1 U664 ( .B(n787), .A(n786), .S(n823), .Y(n785) );
  INVX1 U665 ( .A(n823), .Y(n805) );
  MUX2X1 U666 ( .B(\mem<15><2> ), .A(\mem<14><2> ), .S(n809), .Y(n725) );
  INVX8 U667 ( .A(n642), .Y(n643) );
  BUFX2 U668 ( .A(n822), .Y(n644) );
  INVX1 U669 ( .A(n642), .Y(n645) );
  MUX2X1 U670 ( .B(n692), .A(n691), .S(n646), .Y(n690) );
  MUX2X1 U671 ( .B(\mem<11><0> ), .A(\mem<10><0> ), .S(n644), .Y(n668) );
  BUFX2 U672 ( .A(write), .Y(n647) );
  MUX2X1 U673 ( .B(n649), .A(n650), .S(n808), .Y(n648) );
  MUX2X1 U674 ( .B(n652), .A(n653), .S(n808), .Y(n651) );
  MUX2X1 U675 ( .B(n655), .A(n656), .S(n808), .Y(n654) );
  MUX2X1 U676 ( .B(n658), .A(n659), .S(n808), .Y(n657) );
  MUX2X1 U677 ( .B(n661), .A(n662), .S(N13), .Y(n660) );
  MUX2X1 U678 ( .B(n664), .A(n665), .S(n808), .Y(n663) );
  MUX2X1 U679 ( .B(n667), .A(n668), .S(n808), .Y(n666) );
  MUX2X1 U680 ( .B(n670), .A(n671), .S(n808), .Y(n669) );
  MUX2X1 U681 ( .B(n676), .A(n677), .S(N13), .Y(n675) );
  MUX2X1 U682 ( .B(n679), .A(n680), .S(n808), .Y(n678) );
  MUX2X1 U683 ( .B(n682), .A(n683), .S(n808), .Y(n681) );
  MUX2X1 U684 ( .B(n685), .A(n686), .S(n808), .Y(n684) );
  MUX2X1 U685 ( .B(n688), .A(n689), .S(n808), .Y(n687) );
  MUX2X1 U686 ( .B(n694), .A(n695), .S(n807), .Y(n693) );
  MUX2X1 U687 ( .B(n697), .A(n698), .S(n807), .Y(n696) );
  MUX2X1 U688 ( .B(n700), .A(n701), .S(n807), .Y(n699) );
  MUX2X1 U689 ( .B(n703), .A(n704), .S(n807), .Y(n702) );
  MUX2X1 U690 ( .B(n706), .A(n707), .S(N13), .Y(n705) );
  MUX2X1 U691 ( .B(n709), .A(n710), .S(n807), .Y(n708) );
  MUX2X1 U692 ( .B(n712), .A(n713), .S(n807), .Y(n711) );
  MUX2X1 U693 ( .B(n715), .A(n716), .S(n807), .Y(n714) );
  MUX2X1 U694 ( .B(n718), .A(n719), .S(n807), .Y(n717) );
  MUX2X1 U695 ( .B(n721), .A(n722), .S(N13), .Y(n720) );
  MUX2X1 U696 ( .B(n724), .A(n725), .S(n807), .Y(n723) );
  MUX2X1 U697 ( .B(n727), .A(n728), .S(n807), .Y(n726) );
  MUX2X1 U698 ( .B(n730), .A(n731), .S(n807), .Y(n729) );
  MUX2X1 U699 ( .B(n733), .A(n734), .S(n807), .Y(n732) );
  MUX2X1 U700 ( .B(n736), .A(n737), .S(N13), .Y(n735) );
  MUX2X1 U701 ( .B(n739), .A(n740), .S(n806), .Y(n738) );
  MUX2X1 U702 ( .B(n742), .A(n743), .S(n806), .Y(n741) );
  MUX2X1 U703 ( .B(n745), .A(n746), .S(n806), .Y(n744) );
  MUX2X1 U704 ( .B(n748), .A(n749), .S(n806), .Y(n747) );
  MUX2X1 U705 ( .B(n751), .A(n752), .S(N13), .Y(n750) );
  MUX2X1 U706 ( .B(n754), .A(n755), .S(n806), .Y(n753) );
  MUX2X1 U707 ( .B(n757), .A(n758), .S(n806), .Y(n756) );
  MUX2X1 U708 ( .B(n760), .A(n761), .S(n806), .Y(n759) );
  MUX2X1 U709 ( .B(n763), .A(n764), .S(n806), .Y(n762) );
  MUX2X1 U710 ( .B(n766), .A(n213), .S(N13), .Y(n765) );
  MUX2X1 U711 ( .B(n768), .A(n769), .S(n806), .Y(n767) );
  MUX2X1 U712 ( .B(n771), .A(n772), .S(n806), .Y(n770) );
  MUX2X1 U713 ( .B(n774), .A(n775), .S(n806), .Y(n773) );
  MUX2X1 U714 ( .B(n777), .A(n778), .S(n806), .Y(n776) );
  MUX2X1 U715 ( .B(n780), .A(n781), .S(N13), .Y(n779) );
  MUX2X1 U716 ( .B(n783), .A(n784), .S(n805), .Y(n782) );
  MUX2X1 U717 ( .B(n789), .A(n790), .S(n805), .Y(n788) );
  MUX2X1 U718 ( .B(n792), .A(n793), .S(n805), .Y(n791) );
  MUX2X1 U719 ( .B(n795), .A(n796), .S(N13), .Y(n794) );
  MUX2X1 U720 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n643), .Y(n650) );
  MUX2X1 U721 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n643), .Y(n649) );
  MUX2X1 U722 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n643), .Y(n653) );
  MUX2X1 U723 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n643), .Y(n652) );
  MUX2X1 U724 ( .B(n651), .A(n648), .S(n803), .Y(n662) );
  MUX2X1 U725 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n814), .Y(n656) );
  MUX2X1 U726 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n812), .Y(n655) );
  MUX2X1 U727 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n814), .Y(n659) );
  MUX2X1 U728 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n814), .Y(n658) );
  MUX2X1 U729 ( .B(n657), .A(n654), .S(n803), .Y(n661) );
  MUX2X1 U730 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n812), .Y(n665) );
  MUX2X1 U731 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n645), .Y(n664) );
  MUX2X1 U732 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n812), .Y(n667) );
  MUX2X1 U733 ( .B(n666), .A(n663), .S(n803), .Y(n677) );
  MUX2X1 U734 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n813), .Y(n671) );
  MUX2X1 U735 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n812), .Y(n670) );
  MUX2X1 U736 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n814), .Y(n674) );
  MUX2X1 U737 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n643), .Y(n673) );
  MUX2X1 U738 ( .B(n672), .A(n669), .S(n803), .Y(n676) );
  MUX2X1 U739 ( .B(n675), .A(n660), .S(N14), .Y(n797) );
  MUX2X1 U740 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n643), .Y(n680) );
  MUX2X1 U741 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n812), .Y(n679) );
  MUX2X1 U742 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n812), .Y(n683) );
  MUX2X1 U743 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n812), .Y(n682) );
  MUX2X1 U744 ( .B(n681), .A(n678), .S(n803), .Y(n692) );
  MUX2X1 U745 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n813), .Y(n686) );
  MUX2X1 U746 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n812), .Y(n685) );
  MUX2X1 U747 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n813), .Y(n689) );
  MUX2X1 U748 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n813), .Y(n688) );
  MUX2X1 U749 ( .B(n687), .A(n684), .S(n803), .Y(n691) );
  MUX2X1 U750 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n813), .Y(n695) );
  MUX2X1 U751 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n814), .Y(n694) );
  MUX2X1 U752 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n813), .Y(n698) );
  MUX2X1 U753 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n813), .Y(n697) );
  MUX2X1 U754 ( .B(n696), .A(n693), .S(n803), .Y(n707) );
  MUX2X1 U755 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n813), .Y(n701) );
  MUX2X1 U756 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n814), .Y(n700) );
  MUX2X1 U757 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n645), .Y(n704) );
  MUX2X1 U758 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n814), .Y(n703) );
  MUX2X1 U759 ( .B(n702), .A(n699), .S(n803), .Y(n706) );
  MUX2X1 U760 ( .B(n705), .A(n690), .S(N14), .Y(n798) );
  MUX2X1 U761 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n813), .Y(n710) );
  MUX2X1 U762 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n814), .Y(n709) );
  MUX2X1 U763 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n812), .Y(n713) );
  MUX2X1 U764 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n814), .Y(n712) );
  MUX2X1 U765 ( .B(n711), .A(n708), .S(n803), .Y(n722) );
  MUX2X1 U766 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n813), .Y(n716) );
  MUX2X1 U767 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n813), .Y(n715) );
  MUX2X1 U768 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n813), .Y(n719) );
  MUX2X1 U769 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n813), .Y(n718) );
  MUX2X1 U770 ( .B(n717), .A(n714), .S(n803), .Y(n721) );
  MUX2X1 U771 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n643), .Y(n724) );
  MUX2X1 U772 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n814), .Y(n728) );
  MUX2X1 U773 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n814), .Y(n727) );
  MUX2X1 U774 ( .B(n726), .A(n723), .S(n803), .Y(n737) );
  MUX2X1 U775 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n813), .Y(n731) );
  MUX2X1 U776 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n643), .Y(n730) );
  MUX2X1 U777 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n814), .Y(n734) );
  MUX2X1 U778 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n643), .Y(n733) );
  MUX2X1 U779 ( .B(n732), .A(n729), .S(n803), .Y(n736) );
  MUX2X1 U780 ( .B(n735), .A(n720), .S(N14), .Y(n799) );
  MUX2X1 U781 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n810), .Y(n740) );
  MUX2X1 U782 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n811), .Y(n739) );
  MUX2X1 U783 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n811), .Y(n743) );
  MUX2X1 U784 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n811), .Y(n742) );
  MUX2X1 U785 ( .B(n741), .A(n738), .S(n802), .Y(n752) );
  MUX2X1 U786 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n810), .Y(n746) );
  MUX2X1 U787 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n810), .Y(n745) );
  MUX2X1 U788 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n811), .Y(n749) );
  MUX2X1 U789 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n810), .Y(n748) );
  MUX2X1 U790 ( .B(n747), .A(n744), .S(n802), .Y(n751) );
  MUX2X1 U791 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n810), .Y(n754) );
  MUX2X1 U792 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n811), .Y(n758) );
  MUX2X1 U793 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n814), .Y(n757) );
  MUX2X1 U794 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n811), .Y(n761) );
  MUX2X1 U795 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n810), .Y(n760) );
  MUX2X1 U796 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n643), .Y(n764) );
  MUX2X1 U797 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n812), .Y(n763) );
  MUX2X1 U798 ( .B(n762), .A(n759), .S(n802), .Y(n766) );
  MUX2X1 U799 ( .B(n765), .A(n750), .S(N14), .Y(n800) );
  MUX2X1 U800 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n811), .Y(n769) );
  MUX2X1 U801 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n810), .Y(n768) );
  MUX2X1 U802 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n810), .Y(n772) );
  MUX2X1 U803 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n810), .Y(n771) );
  MUX2X1 U804 ( .B(n770), .A(n767), .S(n802), .Y(n781) );
  MUX2X1 U805 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n811), .Y(n775) );
  MUX2X1 U806 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n811), .Y(n774) );
  MUX2X1 U807 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n811), .Y(n778) );
  MUX2X1 U808 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n811), .Y(n777) );
  MUX2X1 U809 ( .B(n776), .A(n773), .S(n802), .Y(n780) );
  MUX2X1 U810 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n810), .Y(n784) );
  MUX2X1 U811 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n810), .Y(n783) );
  MUX2X1 U812 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n813), .Y(n787) );
  MUX2X1 U813 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n813), .Y(n786) );
  MUX2X1 U814 ( .B(n785), .A(n782), .S(n802), .Y(n796) );
  MUX2X1 U815 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n810), .Y(n790) );
  MUX2X1 U816 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n811), .Y(n789) );
  MUX2X1 U817 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n813), .Y(n793) );
  MUX2X1 U818 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n813), .Y(n792) );
  MUX2X1 U819 ( .B(n791), .A(n788), .S(n802), .Y(n795) );
  MUX2X1 U820 ( .B(n794), .A(n779), .S(N14), .Y(n801) );
  INVX8 U821 ( .A(n825), .Y(n803) );
  INVX8 U822 ( .A(N11), .Y(n804) );
  INVX8 U823 ( .A(n823), .Y(n806) );
  INVX8 U824 ( .A(n823), .Y(n807) );
  INVX8 U825 ( .A(n804), .Y(n808) );
  INVX8 U826 ( .A(n809), .Y(n810) );
  INVX8 U827 ( .A(n809), .Y(n811) );
  INVX8 U828 ( .A(n642), .Y(n812) );
  INVX8 U829 ( .A(n642), .Y(n813) );
  INVX8 U830 ( .A(n809), .Y(n814) );
  INVX1 U831 ( .A(n799), .Y(N19) );
  INVX1 U832 ( .A(n798), .Y(N20) );
  INVX1 U833 ( .A(n800), .Y(N18) );
  INVX1 U834 ( .A(n797), .Y(N21) );
  INVX8 U835 ( .A(N11), .Y(n823) );
  INVX8 U836 ( .A(N12), .Y(n825) );
  AND2X2 U837 ( .A(n2), .B(N21), .Y(\data_out<0> ) );
  AND2X2 U838 ( .A(n2), .B(N20), .Y(\data_out<1> ) );
  AND2X2 U839 ( .A(n503), .B(N19), .Y(\data_out<2> ) );
  AND2X2 U840 ( .A(n504), .B(N18), .Y(\data_out<3> ) );
  AND2X2 U841 ( .A(N17), .B(n503), .Y(\data_out<4> ) );
endmodule


module memc_Size1_0 ( .data_out(\data_out<0> ), .addr({\addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
    .data_in(\data_in<0> ), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<0> , write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><0> , \mem<1><0> , \mem<2><0> ,
         \mem<3><0> , \mem<4><0> , \mem<5><0> , \mem<6><0> , \mem<7><0> ,
         \mem<8><0> , \mem<9><0> , \mem<10><0> , \mem<11><0> , \mem<12><0> ,
         \mem<13><0> , \mem<14><0> , \mem<15><0> , \mem<16><0> , \mem<17><0> ,
         \mem<18><0> , \mem<19><0> , \mem<20><0> , \mem<21><0> , \mem<22><0> ,
         \mem<23><0> , \mem<24><0> , \mem<25><0> , \mem<26><0> , \mem<27><0> ,
         \mem<28><0> , \mem<29><0> , \mem<30><0> , \mem<31><0> , N17, n1, n2,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><0>  ( .D(n203), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n204), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n205), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n206), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n207), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n208), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n209), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n210), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n211), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n212), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n213), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n214), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n215), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n216), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n217), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n218), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n219), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n220), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n221), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n222), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n223), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n224), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n225), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n226), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n227), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n228), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n229), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n230), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n231), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n232), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n233), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n234), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(\data_in<0> ), .B(n143), .Y(n95) );
  AND2X2 U3 ( .A(\data_in<0> ), .B(n144), .Y(n94) );
  AND2X2 U4 ( .A(\data_in<0> ), .B(n146), .Y(n107) );
  INVX1 U5 ( .A(n140), .Y(N17) );
  INVX1 U6 ( .A(n150), .Y(n141) );
  INVX1 U7 ( .A(rst), .Y(n147) );
  OR2X1 U8 ( .A(write), .B(n58), .Y(n2) );
  INVX1 U9 ( .A(N12), .Y(n152) );
  INVX1 U10 ( .A(n96), .Y(n186) );
  INVX1 U11 ( .A(n97), .Y(n189) );
  INVX1 U12 ( .A(n98), .Y(n192) );
  INVX1 U13 ( .A(n99), .Y(n195) );
  INVX1 U14 ( .A(n100), .Y(n198) );
  INVX2 U15 ( .A(n148), .Y(n142) );
  AND2X1 U16 ( .A(n148), .B(n56), .Y(n103) );
  INVX2 U17 ( .A(n109), .Y(n1) );
  INVX1 U18 ( .A(n109), .Y(n145) );
  INVX1 U19 ( .A(n145), .Y(n166) );
  INVX1 U20 ( .A(n2), .Y(\data_out<0> ) );
  AND2X2 U21 ( .A(\data_in<0> ), .B(n166), .Y(n4) );
  AND2X2 U22 ( .A(n105), .B(n94), .Y(n5) );
  INVX1 U23 ( .A(n5), .Y(n6) );
  AND2X2 U24 ( .A(n101), .B(n94), .Y(n7) );
  INVX1 U25 ( .A(n7), .Y(n8) );
  AND2X2 U26 ( .A(n186), .B(n94), .Y(n9) );
  INVX1 U27 ( .A(n9), .Y(n10) );
  AND2X2 U28 ( .A(n189), .B(n94), .Y(n11) );
  INVX1 U29 ( .A(n11), .Y(n12) );
  AND2X2 U30 ( .A(n192), .B(n94), .Y(n13) );
  INVX1 U31 ( .A(n13), .Y(n14) );
  AND2X2 U32 ( .A(n195), .B(n94), .Y(n15) );
  INVX1 U33 ( .A(n15), .Y(n16) );
  AND2X2 U34 ( .A(n198), .B(n94), .Y(n17) );
  INVX1 U35 ( .A(n17), .Y(n18) );
  AND2X2 U36 ( .A(n103), .B(n94), .Y(n19) );
  INVX1 U37 ( .A(n19), .Y(n20) );
  AND2X2 U38 ( .A(n105), .B(n95), .Y(n21) );
  INVX1 U39 ( .A(n21), .Y(n22) );
  AND2X2 U40 ( .A(n101), .B(n95), .Y(n23) );
  INVX1 U41 ( .A(n23), .Y(n24) );
  AND2X2 U42 ( .A(n186), .B(n95), .Y(n25) );
  INVX1 U43 ( .A(n25), .Y(n26) );
  AND2X2 U44 ( .A(n189), .B(n95), .Y(n27) );
  INVX1 U45 ( .A(n27), .Y(n28) );
  AND2X2 U46 ( .A(n192), .B(n95), .Y(n29) );
  INVX1 U47 ( .A(n29), .Y(n30) );
  AND2X2 U48 ( .A(n195), .B(n95), .Y(n31) );
  INVX1 U49 ( .A(n31), .Y(n32) );
  AND2X2 U50 ( .A(n198), .B(n95), .Y(n33) );
  INVX1 U51 ( .A(n33), .Y(n34) );
  AND2X2 U52 ( .A(n103), .B(n95), .Y(n35) );
  INVX1 U53 ( .A(n35), .Y(n36) );
  AND2X2 U54 ( .A(n105), .B(n4), .Y(n37) );
  INVX1 U55 ( .A(n37), .Y(n38) );
  AND2X2 U56 ( .A(n101), .B(n4), .Y(n39) );
  INVX1 U57 ( .A(n39), .Y(n40) );
  AND2X2 U58 ( .A(n186), .B(n4), .Y(n41) );
  INVX1 U59 ( .A(n41), .Y(n42) );
  AND2X2 U60 ( .A(n189), .B(n4), .Y(n43) );
  INVX1 U61 ( .A(n43), .Y(n44) );
  AND2X2 U62 ( .A(n192), .B(n4), .Y(n45) );
  INVX1 U63 ( .A(n45), .Y(n46) );
  AND2X2 U64 ( .A(n195), .B(n4), .Y(n47) );
  INVX1 U65 ( .A(n47), .Y(n48) );
  AND2X2 U66 ( .A(n198), .B(n4), .Y(n49) );
  INVX1 U67 ( .A(n49), .Y(n50) );
  AND2X2 U68 ( .A(n103), .B(n4), .Y(n51) );
  INVX1 U69 ( .A(n51), .Y(n52) );
  BUFX2 U70 ( .A(n156), .Y(n53) );
  OR2X2 U71 ( .A(\addr<5> ), .B(n53), .Y(n54) );
  INVX1 U72 ( .A(n152), .Y(n151) );
  INVX1 U73 ( .A(n150), .Y(n149) );
  OR2X1 U74 ( .A(n149), .B(n151), .Y(n55) );
  INVX1 U75 ( .A(n55), .Y(n56) );
  AND2X1 U76 ( .A(N17), .B(n147), .Y(n57) );
  INVX1 U77 ( .A(n57), .Y(n58) );
  OR2X1 U78 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n59) );
  INVX1 U79 ( .A(n59), .Y(n60) );
  AND2X1 U80 ( .A(n151), .B(n149), .Y(n93) );
  BUFX2 U81 ( .A(n187), .Y(n96) );
  BUFX2 U82 ( .A(n190), .Y(n97) );
  BUFX2 U83 ( .A(n193), .Y(n98) );
  BUFX2 U84 ( .A(n196), .Y(n99) );
  BUFX2 U85 ( .A(n199), .Y(n100) );
  AND2X1 U86 ( .A(n148), .B(n93), .Y(n101) );
  INVX1 U87 ( .A(n101), .Y(n102) );
  INVX1 U88 ( .A(n103), .Y(n104) );
  AND2X1 U89 ( .A(n142), .B(n93), .Y(n105) );
  INVX1 U90 ( .A(n105), .Y(n106) );
  INVX1 U91 ( .A(n107), .Y(n108) );
  NOR3X1 U92 ( .A(n155), .B(n54), .C(N13), .Y(n109) );
  INVX1 U93 ( .A(N11), .Y(n150) );
  MUX2X1 U94 ( .B(n111), .A(n112), .S(n141), .Y(n110) );
  MUX2X1 U95 ( .B(n114), .A(n115), .S(n141), .Y(n113) );
  MUX2X1 U96 ( .B(n117), .A(n118), .S(n141), .Y(n116) );
  MUX2X1 U97 ( .B(n120), .A(n121), .S(n141), .Y(n119) );
  MUX2X1 U98 ( .B(n123), .A(n124), .S(n153), .Y(n122) );
  MUX2X1 U99 ( .B(n126), .A(n127), .S(n141), .Y(n125) );
  MUX2X1 U100 ( .B(n129), .A(n130), .S(n141), .Y(n128) );
  MUX2X1 U101 ( .B(n132), .A(n133), .S(n141), .Y(n131) );
  MUX2X1 U102 ( .B(n135), .A(n136), .S(n141), .Y(n134) );
  MUX2X1 U103 ( .B(n138), .A(n139), .S(n153), .Y(n137) );
  MUX2X1 U104 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n142), .Y(n112) );
  MUX2X1 U105 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n142), .Y(n111) );
  MUX2X1 U106 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n142), .Y(n115) );
  MUX2X1 U107 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n142), .Y(n114) );
  MUX2X1 U108 ( .B(n113), .A(n110), .S(n151), .Y(n124) );
  MUX2X1 U109 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n142), .Y(n118) );
  MUX2X1 U110 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n142), .Y(n117) );
  MUX2X1 U111 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n142), .Y(n121) );
  MUX2X1 U112 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n142), .Y(n120) );
  MUX2X1 U113 ( .B(n119), .A(n116), .S(n151), .Y(n123) );
  MUX2X1 U114 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n142), .Y(n127) );
  MUX2X1 U115 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n142), .Y(n126) );
  MUX2X1 U116 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n142), .Y(n130) );
  MUX2X1 U117 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n142), .Y(n129) );
  MUX2X1 U118 ( .B(n128), .A(n125), .S(n151), .Y(n139) );
  MUX2X1 U119 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n142), .Y(n133) );
  MUX2X1 U120 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n142), .Y(n132) );
  MUX2X1 U121 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n142), .Y(n136) );
  MUX2X1 U122 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n142), .Y(n135) );
  MUX2X1 U123 ( .B(n134), .A(n131), .S(n151), .Y(n138) );
  MUX2X1 U124 ( .B(n137), .A(n122), .S(N14), .Y(n140) );
  NOR3X1 U125 ( .A(N13), .B(n54), .C(N14), .Y(n143) );
  INVX4 U126 ( .A(n143), .Y(n201) );
  INVX1 U127 ( .A(N13), .Y(n154) );
  NOR3X1 U128 ( .A(n154), .B(n54), .C(N14), .Y(n144) );
  INVX4 U129 ( .A(n144), .Y(n182) );
  INVX1 U130 ( .A(N14), .Y(n155) );
  NOR3X1 U131 ( .A(n155), .B(n154), .C(n54), .Y(n146) );
  INVX2 U132 ( .A(n146), .Y(n164) );
  INVX1 U133 ( .A(n154), .Y(n153) );
  INVX1 U134 ( .A(N10), .Y(n148) );
  NAND3X1 U135 ( .A(n60), .B(n147), .C(write), .Y(n156) );
  OAI21X1 U136 ( .A(n164), .B(n106), .C(\mem<31><0> ), .Y(n157) );
  OAI21X1 U137 ( .A(n108), .B(n106), .C(n157), .Y(n234) );
  OAI21X1 U138 ( .A(n102), .B(n164), .C(\mem<30><0> ), .Y(n158) );
  OAI21X1 U139 ( .A(n102), .B(n108), .C(n158), .Y(n233) );
  NAND3X1 U140 ( .A(n142), .B(n151), .C(n150), .Y(n187) );
  OAI21X1 U141 ( .A(n96), .B(n164), .C(\mem<29><0> ), .Y(n159) );
  OAI21X1 U142 ( .A(n96), .B(n108), .C(n159), .Y(n232) );
  NAND3X1 U143 ( .A(n151), .B(n150), .C(n148), .Y(n190) );
  OAI21X1 U144 ( .A(n97), .B(n164), .C(\mem<28><0> ), .Y(n160) );
  OAI21X1 U145 ( .A(n97), .B(n108), .C(n160), .Y(n231) );
  NAND3X1 U146 ( .A(n142), .B(n149), .C(n152), .Y(n193) );
  OAI21X1 U147 ( .A(n98), .B(n164), .C(\mem<27><0> ), .Y(n161) );
  OAI21X1 U148 ( .A(n98), .B(n108), .C(n161), .Y(n230) );
  NAND3X1 U149 ( .A(n152), .B(n149), .C(n148), .Y(n196) );
  OAI21X1 U150 ( .A(n99), .B(n164), .C(\mem<26><0> ), .Y(n162) );
  OAI21X1 U151 ( .A(n99), .B(n108), .C(n162), .Y(n229) );
  NAND3X1 U152 ( .A(n142), .B(n152), .C(n150), .Y(n199) );
  OAI21X1 U153 ( .A(n100), .B(n164), .C(\mem<25><0> ), .Y(n163) );
  OAI21X1 U154 ( .A(n100), .B(n108), .C(n163), .Y(n228) );
  OAI21X1 U155 ( .A(n104), .B(n164), .C(\mem<24><0> ), .Y(n165) );
  OAI21X1 U156 ( .A(n104), .B(n108), .C(n165), .Y(n227) );
  OAI21X1 U157 ( .A(n1), .B(n106), .C(\mem<23><0> ), .Y(n167) );
  NAND2X1 U158 ( .A(n38), .B(n167), .Y(n226) );
  OAI21X1 U159 ( .A(n1), .B(n102), .C(\mem<22><0> ), .Y(n168) );
  NAND2X1 U160 ( .A(n40), .B(n168), .Y(n225) );
  OAI21X1 U161 ( .A(n1), .B(n96), .C(\mem<21><0> ), .Y(n169) );
  NAND2X1 U162 ( .A(n42), .B(n169), .Y(n224) );
  OAI21X1 U163 ( .A(n1), .B(n97), .C(\mem<20><0> ), .Y(n170) );
  NAND2X1 U164 ( .A(n44), .B(n170), .Y(n223) );
  OAI21X1 U165 ( .A(n1), .B(n98), .C(\mem<19><0> ), .Y(n171) );
  NAND2X1 U166 ( .A(n46), .B(n171), .Y(n222) );
  OAI21X1 U167 ( .A(n1), .B(n99), .C(\mem<18><0> ), .Y(n172) );
  NAND2X1 U168 ( .A(n48), .B(n172), .Y(n221) );
  OAI21X1 U169 ( .A(n1), .B(n100), .C(\mem<17><0> ), .Y(n173) );
  NAND2X1 U170 ( .A(n50), .B(n173), .Y(n220) );
  OAI21X1 U171 ( .A(n145), .B(n104), .C(\mem<16><0> ), .Y(n174) );
  NAND2X1 U172 ( .A(n52), .B(n174), .Y(n219) );
  OAI21X1 U173 ( .A(n182), .B(n106), .C(\mem<15><0> ), .Y(n175) );
  NAND2X1 U174 ( .A(n6), .B(n175), .Y(n218) );
  OAI21X1 U175 ( .A(n182), .B(n102), .C(\mem<14><0> ), .Y(n176) );
  NAND2X1 U176 ( .A(n8), .B(n176), .Y(n217) );
  OAI21X1 U177 ( .A(n182), .B(n96), .C(\mem<13><0> ), .Y(n177) );
  NAND2X1 U178 ( .A(n10), .B(n177), .Y(n216) );
  OAI21X1 U179 ( .A(n182), .B(n97), .C(\mem<12><0> ), .Y(n178) );
  NAND2X1 U180 ( .A(n12), .B(n178), .Y(n215) );
  OAI21X1 U181 ( .A(n182), .B(n98), .C(\mem<11><0> ), .Y(n179) );
  NAND2X1 U182 ( .A(n14), .B(n179), .Y(n214) );
  OAI21X1 U183 ( .A(n182), .B(n99), .C(\mem<10><0> ), .Y(n180) );
  NAND2X1 U184 ( .A(n16), .B(n180), .Y(n213) );
  OAI21X1 U185 ( .A(n182), .B(n100), .C(\mem<9><0> ), .Y(n181) );
  NAND2X1 U186 ( .A(n18), .B(n181), .Y(n212) );
  OAI21X1 U187 ( .A(n182), .B(n104), .C(\mem<8><0> ), .Y(n183) );
  NAND2X1 U188 ( .A(n20), .B(n183), .Y(n211) );
  OAI21X1 U189 ( .A(n201), .B(n106), .C(\mem<7><0> ), .Y(n184) );
  NAND2X1 U190 ( .A(n22), .B(n184), .Y(n210) );
  OAI21X1 U191 ( .A(n201), .B(n102), .C(\mem<6><0> ), .Y(n185) );
  NAND2X1 U192 ( .A(n24), .B(n185), .Y(n209) );
  OAI21X1 U193 ( .A(n201), .B(n96), .C(\mem<5><0> ), .Y(n188) );
  NAND2X1 U194 ( .A(n26), .B(n188), .Y(n208) );
  OAI21X1 U195 ( .A(n201), .B(n97), .C(\mem<4><0> ), .Y(n191) );
  NAND2X1 U196 ( .A(n28), .B(n191), .Y(n207) );
  OAI21X1 U197 ( .A(n201), .B(n98), .C(\mem<3><0> ), .Y(n194) );
  NAND2X1 U198 ( .A(n30), .B(n194), .Y(n206) );
  OAI21X1 U199 ( .A(n201), .B(n99), .C(\mem<2><0> ), .Y(n197) );
  NAND2X1 U200 ( .A(n32), .B(n197), .Y(n205) );
  OAI21X1 U201 ( .A(n201), .B(n100), .C(\mem<1><0> ), .Y(n200) );
  NAND2X1 U202 ( .A(n34), .B(n200), .Y(n204) );
  OAI21X1 U203 ( .A(n201), .B(n104), .C(\mem<0><0> ), .Y(n202) );
  NAND2X1 U204 ( .A(n36), .B(n202), .Y(n203) );
endmodule


module memv_0 ( data_out, .addr({\addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), data_in, write, clk, rst, 
        createdump, .file_id({\file_id<4> , \file_id<3> , \file_id<2> , 
        \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , data_in, write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output data_out;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \mem<0> , \mem<1> , \mem<2> ,
         \mem<3> , \mem<4> , \mem<5> , \mem<6> , \mem<7> , \mem<8> , \mem<9> ,
         \mem<10> , \mem<11> , \mem<12> , \mem<13> , \mem<14> , \mem<15> ,
         \mem<16> , \mem<17> , \mem<18> , \mem<19> , \mem<20> , \mem<21> ,
         \mem<22> , \mem<23> , \mem<24> , \mem<25> , \mem<26> , \mem<27> ,
         \mem<28> , \mem<29> , \mem<30> , \mem<31> , \mem<32> , \mem<33> ,
         \mem<34> , \mem<35> , \mem<36> , \mem<37> , \mem<38> , \mem<39> ,
         \mem<40> , \mem<41> , \mem<42> , \mem<43> , \mem<44> , \mem<45> ,
         \mem<46> , \mem<47> , \mem<48> , \mem<49> , \mem<50> , \mem<51> ,
         \mem<52> , \mem<53> , \mem<54> , \mem<55> , \mem<56> , \mem<57> ,
         \mem<58> , \mem<59> , \mem<60> , \mem<61> , \mem<62> , \mem<63> ,
         \mem<64> , \mem<65> , \mem<66> , \mem<67> , \mem<68> , \mem<69> ,
         \mem<70> , \mem<71> , \mem<72> , \mem<73> , \mem<74> , \mem<75> ,
         \mem<76> , \mem<77> , \mem<78> , \mem<79> , \mem<80> , \mem<81> ,
         \mem<82> , \mem<83> , \mem<84> , \mem<85> , \mem<86> , \mem<87> ,
         \mem<88> , \mem<89> , \mem<90> , \mem<91> , \mem<92> , \mem<93> ,
         \mem<94> , \mem<95> , \mem<96> , \mem<97> , \mem<98> , \mem<99> ,
         \mem<100> , \mem<101> , \mem<102> , \mem<103> , \mem<104> ,
         \mem<105> , \mem<106> , \mem<107> , \mem<108> , \mem<109> ,
         \mem<110> , \mem<111> , \mem<112> , \mem<113> , \mem<114> ,
         \mem<115> , \mem<116> , \mem<117> , \mem<118> , \mem<119> ,
         \mem<120> , \mem<121> , \mem<122> , \mem<123> , \mem<124> ,
         \mem<125> , \mem<126> , \mem<127> , \mem<128> , \mem<129> ,
         \mem<130> , \mem<131> , \mem<132> , \mem<133> , \mem<134> ,
         \mem<135> , \mem<136> , \mem<137> , \mem<138> , \mem<139> ,
         \mem<140> , \mem<141> , \mem<142> , \mem<143> , \mem<144> ,
         \mem<145> , \mem<146> , \mem<147> , \mem<148> , \mem<149> ,
         \mem<150> , \mem<151> , \mem<152> , \mem<153> , \mem<154> ,
         \mem<155> , \mem<156> , \mem<157> , \mem<158> , \mem<159> ,
         \mem<160> , \mem<161> , \mem<162> , \mem<163> , \mem<164> ,
         \mem<165> , \mem<166> , \mem<167> , \mem<168> , \mem<169> ,
         \mem<170> , \mem<171> , \mem<172> , \mem<173> , \mem<174> ,
         \mem<175> , \mem<176> , \mem<177> , \mem<178> , \mem<179> ,
         \mem<180> , \mem<181> , \mem<182> , \mem<183> , \mem<184> ,
         \mem<185> , \mem<186> , \mem<187> , \mem<188> , \mem<189> ,
         \mem<190> , \mem<191> , \mem<192> , \mem<193> , \mem<194> ,
         \mem<195> , \mem<196> , \mem<197> , \mem<198> , \mem<199> ,
         \mem<200> , \mem<201> , \mem<202> , \mem<203> , \mem<204> ,
         \mem<205> , \mem<206> , \mem<207> , \mem<208> , \mem<209> ,
         \mem<210> , \mem<211> , \mem<212> , \mem<213> , \mem<214> ,
         \mem<215> , \mem<216> , \mem<217> , \mem<218> , \mem<219> ,
         \mem<220> , \mem<221> , \mem<222> , \mem<223> , \mem<224> ,
         \mem<225> , \mem<226> , \mem<227> , \mem<228> , \mem<229> ,
         \mem<230> , \mem<231> , \mem<232> , \mem<233> , \mem<234> ,
         \mem<235> , \mem<236> , \mem<237> , \mem<238> , \mem<239> ,
         \mem<240> , \mem<241> , \mem<242> , \mem<243> , \mem<244> ,
         \mem<245> , \mem<246> , \mem<247> , \mem<248> , \mem<249> ,
         \mem<250> , \mem<251> , \mem<252> , \mem<253> , \mem<254> ,
         \mem<255> , N28, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n43, n44, n45, n47, n48, n50, n51, n53, n54, n56, n57, n59, n60,
         n62, n63, n65, n66, n68, n69, n71, n72, n74, n75, n77, n78, n80, n81,
         n83, n84, n86, n87, n89, n93, n95, n112, n114, n130, n131, n133, n149,
         n150, n152, n169, n171, n187, n189, n205, n207, n223, n225, n241,
         n242, n244, n260, n262, n278, n280, n296, n298, n314, n315, n317,
         n333, n335, n351, n353, n354, n360, n362, n369, n374, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511;
  assign N18 = \addr<0> ;
  assign N19 = \addr<1> ;
  assign N20 = \addr<2> ;
  assign N21 = \addr<3> ;
  assign N22 = \addr<4> ;
  assign N23 = \addr<5> ;
  assign N24 = \addr<6> ;
  assign N25 = \addr<7> ;

  DFFPOSX1 \mem_reg<0>  ( .D(n991), .CLK(clk), .Q(\mem<0> ) );
  DFFPOSX1 \mem_reg<1>  ( .D(n992), .CLK(clk), .Q(\mem<1> ) );
  DFFPOSX1 \mem_reg<2>  ( .D(n993), .CLK(clk), .Q(\mem<2> ) );
  DFFPOSX1 \mem_reg<3>  ( .D(n994), .CLK(clk), .Q(\mem<3> ) );
  DFFPOSX1 \mem_reg<4>  ( .D(n995), .CLK(clk), .Q(\mem<4> ) );
  DFFPOSX1 \mem_reg<5>  ( .D(n996), .CLK(clk), .Q(\mem<5> ) );
  DFFPOSX1 \mem_reg<6>  ( .D(n997), .CLK(clk), .Q(\mem<6> ) );
  DFFPOSX1 \mem_reg<7>  ( .D(n998), .CLK(clk), .Q(\mem<7> ) );
  DFFPOSX1 \mem_reg<8>  ( .D(n999), .CLK(clk), .Q(\mem<8> ) );
  DFFPOSX1 \mem_reg<9>  ( .D(n1000), .CLK(clk), .Q(\mem<9> ) );
  DFFPOSX1 \mem_reg<10>  ( .D(n1001), .CLK(clk), .Q(\mem<10> ) );
  DFFPOSX1 \mem_reg<11>  ( .D(n1002), .CLK(clk), .Q(\mem<11> ) );
  DFFPOSX1 \mem_reg<12>  ( .D(n1003), .CLK(clk), .Q(\mem<12> ) );
  DFFPOSX1 \mem_reg<13>  ( .D(n1004), .CLK(clk), .Q(\mem<13> ) );
  DFFPOSX1 \mem_reg<14>  ( .D(n1005), .CLK(clk), .Q(\mem<14> ) );
  DFFPOSX1 \mem_reg<15>  ( .D(n1006), .CLK(clk), .Q(\mem<15> ) );
  DFFPOSX1 \mem_reg<16>  ( .D(n1007), .CLK(clk), .Q(\mem<16> ) );
  DFFPOSX1 \mem_reg<17>  ( .D(n1008), .CLK(clk), .Q(\mem<17> ) );
  DFFPOSX1 \mem_reg<18>  ( .D(n1009), .CLK(clk), .Q(\mem<18> ) );
  DFFPOSX1 \mem_reg<19>  ( .D(n1010), .CLK(clk), .Q(\mem<19> ) );
  DFFPOSX1 \mem_reg<20>  ( .D(n1011), .CLK(clk), .Q(\mem<20> ) );
  DFFPOSX1 \mem_reg<21>  ( .D(n1012), .CLK(clk), .Q(\mem<21> ) );
  DFFPOSX1 \mem_reg<22>  ( .D(n1013), .CLK(clk), .Q(\mem<22> ) );
  DFFPOSX1 \mem_reg<23>  ( .D(n1014), .CLK(clk), .Q(\mem<23> ) );
  DFFPOSX1 \mem_reg<24>  ( .D(n1015), .CLK(clk), .Q(\mem<24> ) );
  DFFPOSX1 \mem_reg<25>  ( .D(n1016), .CLK(clk), .Q(\mem<25> ) );
  DFFPOSX1 \mem_reg<26>  ( .D(n1017), .CLK(clk), .Q(\mem<26> ) );
  DFFPOSX1 \mem_reg<27>  ( .D(n1018), .CLK(clk), .Q(\mem<27> ) );
  DFFPOSX1 \mem_reg<28>  ( .D(n1019), .CLK(clk), .Q(\mem<28> ) );
  DFFPOSX1 \mem_reg<29>  ( .D(n1020), .CLK(clk), .Q(\mem<29> ) );
  DFFPOSX1 \mem_reg<30>  ( .D(n1021), .CLK(clk), .Q(\mem<30> ) );
  DFFPOSX1 \mem_reg<31>  ( .D(n1022), .CLK(clk), .Q(\mem<31> ) );
  DFFPOSX1 \mem_reg<32>  ( .D(n1023), .CLK(clk), .Q(\mem<32> ) );
  DFFPOSX1 \mem_reg<33>  ( .D(n1024), .CLK(clk), .Q(\mem<33> ) );
  DFFPOSX1 \mem_reg<34>  ( .D(n1025), .CLK(clk), .Q(\mem<34> ) );
  DFFPOSX1 \mem_reg<35>  ( .D(n1026), .CLK(clk), .Q(\mem<35> ) );
  DFFPOSX1 \mem_reg<36>  ( .D(n1027), .CLK(clk), .Q(\mem<36> ) );
  DFFPOSX1 \mem_reg<37>  ( .D(n1028), .CLK(clk), .Q(\mem<37> ) );
  DFFPOSX1 \mem_reg<38>  ( .D(n1029), .CLK(clk), .Q(\mem<38> ) );
  DFFPOSX1 \mem_reg<39>  ( .D(n1030), .CLK(clk), .Q(\mem<39> ) );
  DFFPOSX1 \mem_reg<40>  ( .D(n1031), .CLK(clk), .Q(\mem<40> ) );
  DFFPOSX1 \mem_reg<41>  ( .D(n1032), .CLK(clk), .Q(\mem<41> ) );
  DFFPOSX1 \mem_reg<42>  ( .D(n1033), .CLK(clk), .Q(\mem<42> ) );
  DFFPOSX1 \mem_reg<43>  ( .D(n1034), .CLK(clk), .Q(\mem<43> ) );
  DFFPOSX1 \mem_reg<44>  ( .D(n1035), .CLK(clk), .Q(\mem<44> ) );
  DFFPOSX1 \mem_reg<45>  ( .D(n1036), .CLK(clk), .Q(\mem<45> ) );
  DFFPOSX1 \mem_reg<46>  ( .D(n1037), .CLK(clk), .Q(\mem<46> ) );
  DFFPOSX1 \mem_reg<47>  ( .D(n1038), .CLK(clk), .Q(\mem<47> ) );
  DFFPOSX1 \mem_reg<48>  ( .D(n1039), .CLK(clk), .Q(\mem<48> ) );
  DFFPOSX1 \mem_reg<49>  ( .D(n1040), .CLK(clk), .Q(\mem<49> ) );
  DFFPOSX1 \mem_reg<50>  ( .D(n1041), .CLK(clk), .Q(\mem<50> ) );
  DFFPOSX1 \mem_reg<51>  ( .D(n1042), .CLK(clk), .Q(\mem<51> ) );
  DFFPOSX1 \mem_reg<52>  ( .D(n1043), .CLK(clk), .Q(\mem<52> ) );
  DFFPOSX1 \mem_reg<53>  ( .D(n1044), .CLK(clk), .Q(\mem<53> ) );
  DFFPOSX1 \mem_reg<54>  ( .D(n1045), .CLK(clk), .Q(\mem<54> ) );
  DFFPOSX1 \mem_reg<55>  ( .D(n1046), .CLK(clk), .Q(\mem<55> ) );
  DFFPOSX1 \mem_reg<56>  ( .D(n1047), .CLK(clk), .Q(\mem<56> ) );
  DFFPOSX1 \mem_reg<57>  ( .D(n1048), .CLK(clk), .Q(\mem<57> ) );
  DFFPOSX1 \mem_reg<58>  ( .D(n1049), .CLK(clk), .Q(\mem<58> ) );
  DFFPOSX1 \mem_reg<59>  ( .D(n1050), .CLK(clk), .Q(\mem<59> ) );
  DFFPOSX1 \mem_reg<60>  ( .D(n1051), .CLK(clk), .Q(\mem<60> ) );
  DFFPOSX1 \mem_reg<61>  ( .D(n1052), .CLK(clk), .Q(\mem<61> ) );
  DFFPOSX1 \mem_reg<62>  ( .D(n1053), .CLK(clk), .Q(\mem<62> ) );
  DFFPOSX1 \mem_reg<63>  ( .D(n1054), .CLK(clk), .Q(\mem<63> ) );
  DFFPOSX1 \mem_reg<64>  ( .D(n1055), .CLK(clk), .Q(\mem<64> ) );
  DFFPOSX1 \mem_reg<65>  ( .D(n1056), .CLK(clk), .Q(\mem<65> ) );
  DFFPOSX1 \mem_reg<66>  ( .D(n1057), .CLK(clk), .Q(\mem<66> ) );
  DFFPOSX1 \mem_reg<67>  ( .D(n1058), .CLK(clk), .Q(\mem<67> ) );
  DFFPOSX1 \mem_reg<68>  ( .D(n1059), .CLK(clk), .Q(\mem<68> ) );
  DFFPOSX1 \mem_reg<69>  ( .D(n1060), .CLK(clk), .Q(\mem<69> ) );
  DFFPOSX1 \mem_reg<70>  ( .D(n1061), .CLK(clk), .Q(\mem<70> ) );
  DFFPOSX1 \mem_reg<71>  ( .D(n1062), .CLK(clk), .Q(\mem<71> ) );
  DFFPOSX1 \mem_reg<72>  ( .D(n1063), .CLK(clk), .Q(\mem<72> ) );
  DFFPOSX1 \mem_reg<73>  ( .D(n1064), .CLK(clk), .Q(\mem<73> ) );
  DFFPOSX1 \mem_reg<74>  ( .D(n1065), .CLK(clk), .Q(\mem<74> ) );
  DFFPOSX1 \mem_reg<75>  ( .D(n1066), .CLK(clk), .Q(\mem<75> ) );
  DFFPOSX1 \mem_reg<76>  ( .D(n1067), .CLK(clk), .Q(\mem<76> ) );
  DFFPOSX1 \mem_reg<77>  ( .D(n1068), .CLK(clk), .Q(\mem<77> ) );
  DFFPOSX1 \mem_reg<78>  ( .D(n1069), .CLK(clk), .Q(\mem<78> ) );
  DFFPOSX1 \mem_reg<79>  ( .D(n1070), .CLK(clk), .Q(\mem<79> ) );
  DFFPOSX1 \mem_reg<80>  ( .D(n1071), .CLK(clk), .Q(\mem<80> ) );
  DFFPOSX1 \mem_reg<81>  ( .D(n1072), .CLK(clk), .Q(\mem<81> ) );
  DFFPOSX1 \mem_reg<82>  ( .D(n1073), .CLK(clk), .Q(\mem<82> ) );
  DFFPOSX1 \mem_reg<83>  ( .D(n1074), .CLK(clk), .Q(\mem<83> ) );
  DFFPOSX1 \mem_reg<84>  ( .D(n1075), .CLK(clk), .Q(\mem<84> ) );
  DFFPOSX1 \mem_reg<85>  ( .D(n1076), .CLK(clk), .Q(\mem<85> ) );
  DFFPOSX1 \mem_reg<86>  ( .D(n1077), .CLK(clk), .Q(\mem<86> ) );
  DFFPOSX1 \mem_reg<87>  ( .D(n1078), .CLK(clk), .Q(\mem<87> ) );
  DFFPOSX1 \mem_reg<88>  ( .D(n1079), .CLK(clk), .Q(\mem<88> ) );
  DFFPOSX1 \mem_reg<89>  ( .D(n1080), .CLK(clk), .Q(\mem<89> ) );
  DFFPOSX1 \mem_reg<90>  ( .D(n1081), .CLK(clk), .Q(\mem<90> ) );
  DFFPOSX1 \mem_reg<91>  ( .D(n1082), .CLK(clk), .Q(\mem<91> ) );
  DFFPOSX1 \mem_reg<92>  ( .D(n1083), .CLK(clk), .Q(\mem<92> ) );
  DFFPOSX1 \mem_reg<93>  ( .D(n1084), .CLK(clk), .Q(\mem<93> ) );
  DFFPOSX1 \mem_reg<94>  ( .D(n1085), .CLK(clk), .Q(\mem<94> ) );
  DFFPOSX1 \mem_reg<95>  ( .D(n1086), .CLK(clk), .Q(\mem<95> ) );
  DFFPOSX1 \mem_reg<96>  ( .D(n1087), .CLK(clk), .Q(\mem<96> ) );
  DFFPOSX1 \mem_reg<97>  ( .D(n1088), .CLK(clk), .Q(\mem<97> ) );
  DFFPOSX1 \mem_reg<98>  ( .D(n1089), .CLK(clk), .Q(\mem<98> ) );
  DFFPOSX1 \mem_reg<99>  ( .D(n1090), .CLK(clk), .Q(\mem<99> ) );
  DFFPOSX1 \mem_reg<100>  ( .D(n1091), .CLK(clk), .Q(\mem<100> ) );
  DFFPOSX1 \mem_reg<101>  ( .D(n1092), .CLK(clk), .Q(\mem<101> ) );
  DFFPOSX1 \mem_reg<102>  ( .D(n1093), .CLK(clk), .Q(\mem<102> ) );
  DFFPOSX1 \mem_reg<103>  ( .D(n1094), .CLK(clk), .Q(\mem<103> ) );
  DFFPOSX1 \mem_reg<104>  ( .D(n1095), .CLK(clk), .Q(\mem<104> ) );
  DFFPOSX1 \mem_reg<105>  ( .D(n1096), .CLK(clk), .Q(\mem<105> ) );
  DFFPOSX1 \mem_reg<106>  ( .D(n1097), .CLK(clk), .Q(\mem<106> ) );
  DFFPOSX1 \mem_reg<107>  ( .D(n1098), .CLK(clk), .Q(\mem<107> ) );
  DFFPOSX1 \mem_reg<108>  ( .D(n1099), .CLK(clk), .Q(\mem<108> ) );
  DFFPOSX1 \mem_reg<109>  ( .D(n1100), .CLK(clk), .Q(\mem<109> ) );
  DFFPOSX1 \mem_reg<110>  ( .D(n1101), .CLK(clk), .Q(\mem<110> ) );
  DFFPOSX1 \mem_reg<111>  ( .D(n1102), .CLK(clk), .Q(\mem<111> ) );
  DFFPOSX1 \mem_reg<112>  ( .D(n1103), .CLK(clk), .Q(\mem<112> ) );
  DFFPOSX1 \mem_reg<113>  ( .D(n1104), .CLK(clk), .Q(\mem<113> ) );
  DFFPOSX1 \mem_reg<114>  ( .D(n1105), .CLK(clk), .Q(\mem<114> ) );
  DFFPOSX1 \mem_reg<115>  ( .D(n1106), .CLK(clk), .Q(\mem<115> ) );
  DFFPOSX1 \mem_reg<116>  ( .D(n1107), .CLK(clk), .Q(\mem<116> ) );
  DFFPOSX1 \mem_reg<117>  ( .D(n1108), .CLK(clk), .Q(\mem<117> ) );
  DFFPOSX1 \mem_reg<118>  ( .D(n1109), .CLK(clk), .Q(\mem<118> ) );
  DFFPOSX1 \mem_reg<119>  ( .D(n1110), .CLK(clk), .Q(\mem<119> ) );
  DFFPOSX1 \mem_reg<120>  ( .D(n1111), .CLK(clk), .Q(\mem<120> ) );
  DFFPOSX1 \mem_reg<121>  ( .D(n1112), .CLK(clk), .Q(\mem<121> ) );
  DFFPOSX1 \mem_reg<122>  ( .D(n1113), .CLK(clk), .Q(\mem<122> ) );
  DFFPOSX1 \mem_reg<123>  ( .D(n1114), .CLK(clk), .Q(\mem<123> ) );
  DFFPOSX1 \mem_reg<124>  ( .D(n1115), .CLK(clk), .Q(\mem<124> ) );
  DFFPOSX1 \mem_reg<125>  ( .D(n1116), .CLK(clk), .Q(\mem<125> ) );
  DFFPOSX1 \mem_reg<126>  ( .D(n1117), .CLK(clk), .Q(\mem<126> ) );
  DFFPOSX1 \mem_reg<127>  ( .D(n1118), .CLK(clk), .Q(\mem<127> ) );
  DFFPOSX1 \mem_reg<128>  ( .D(n1119), .CLK(clk), .Q(\mem<128> ) );
  DFFPOSX1 \mem_reg<129>  ( .D(n1120), .CLK(clk), .Q(\mem<129> ) );
  DFFPOSX1 \mem_reg<130>  ( .D(n1121), .CLK(clk), .Q(\mem<130> ) );
  DFFPOSX1 \mem_reg<131>  ( .D(n1122), .CLK(clk), .Q(\mem<131> ) );
  DFFPOSX1 \mem_reg<132>  ( .D(n1123), .CLK(clk), .Q(\mem<132> ) );
  DFFPOSX1 \mem_reg<133>  ( .D(n1124), .CLK(clk), .Q(\mem<133> ) );
  DFFPOSX1 \mem_reg<134>  ( .D(n1125), .CLK(clk), .Q(\mem<134> ) );
  DFFPOSX1 \mem_reg<135>  ( .D(n1126), .CLK(clk), .Q(\mem<135> ) );
  DFFPOSX1 \mem_reg<136>  ( .D(n1127), .CLK(clk), .Q(\mem<136> ) );
  DFFPOSX1 \mem_reg<137>  ( .D(n1128), .CLK(clk), .Q(\mem<137> ) );
  DFFPOSX1 \mem_reg<138>  ( .D(n1129), .CLK(clk), .Q(\mem<138> ) );
  DFFPOSX1 \mem_reg<139>  ( .D(n1130), .CLK(clk), .Q(\mem<139> ) );
  DFFPOSX1 \mem_reg<140>  ( .D(n1131), .CLK(clk), .Q(\mem<140> ) );
  DFFPOSX1 \mem_reg<141>  ( .D(n1132), .CLK(clk), .Q(\mem<141> ) );
  DFFPOSX1 \mem_reg<142>  ( .D(n1133), .CLK(clk), .Q(\mem<142> ) );
  DFFPOSX1 \mem_reg<143>  ( .D(n1134), .CLK(clk), .Q(\mem<143> ) );
  DFFPOSX1 \mem_reg<144>  ( .D(n1135), .CLK(clk), .Q(\mem<144> ) );
  DFFPOSX1 \mem_reg<145>  ( .D(n1136), .CLK(clk), .Q(\mem<145> ) );
  DFFPOSX1 \mem_reg<146>  ( .D(n1137), .CLK(clk), .Q(\mem<146> ) );
  DFFPOSX1 \mem_reg<147>  ( .D(n1138), .CLK(clk), .Q(\mem<147> ) );
  DFFPOSX1 \mem_reg<148>  ( .D(n1139), .CLK(clk), .Q(\mem<148> ) );
  DFFPOSX1 \mem_reg<149>  ( .D(n1140), .CLK(clk), .Q(\mem<149> ) );
  DFFPOSX1 \mem_reg<150>  ( .D(n1141), .CLK(clk), .Q(\mem<150> ) );
  DFFPOSX1 \mem_reg<151>  ( .D(n1142), .CLK(clk), .Q(\mem<151> ) );
  DFFPOSX1 \mem_reg<152>  ( .D(n1143), .CLK(clk), .Q(\mem<152> ) );
  DFFPOSX1 \mem_reg<153>  ( .D(n1144), .CLK(clk), .Q(\mem<153> ) );
  DFFPOSX1 \mem_reg<154>  ( .D(n1145), .CLK(clk), .Q(\mem<154> ) );
  DFFPOSX1 \mem_reg<155>  ( .D(n1146), .CLK(clk), .Q(\mem<155> ) );
  DFFPOSX1 \mem_reg<156>  ( .D(n1147), .CLK(clk), .Q(\mem<156> ) );
  DFFPOSX1 \mem_reg<157>  ( .D(n1148), .CLK(clk), .Q(\mem<157> ) );
  DFFPOSX1 \mem_reg<158>  ( .D(n1149), .CLK(clk), .Q(\mem<158> ) );
  DFFPOSX1 \mem_reg<159>  ( .D(n1150), .CLK(clk), .Q(\mem<159> ) );
  DFFPOSX1 \mem_reg<160>  ( .D(n1151), .CLK(clk), .Q(\mem<160> ) );
  DFFPOSX1 \mem_reg<161>  ( .D(n1152), .CLK(clk), .Q(\mem<161> ) );
  DFFPOSX1 \mem_reg<162>  ( .D(n1153), .CLK(clk), .Q(\mem<162> ) );
  DFFPOSX1 \mem_reg<163>  ( .D(n1154), .CLK(clk), .Q(\mem<163> ) );
  DFFPOSX1 \mem_reg<164>  ( .D(n1155), .CLK(clk), .Q(\mem<164> ) );
  DFFPOSX1 \mem_reg<165>  ( .D(n1156), .CLK(clk), .Q(\mem<165> ) );
  DFFPOSX1 \mem_reg<166>  ( .D(n1157), .CLK(clk), .Q(\mem<166> ) );
  DFFPOSX1 \mem_reg<167>  ( .D(n1158), .CLK(clk), .Q(\mem<167> ) );
  DFFPOSX1 \mem_reg<168>  ( .D(n1159), .CLK(clk), .Q(\mem<168> ) );
  DFFPOSX1 \mem_reg<169>  ( .D(n1160), .CLK(clk), .Q(\mem<169> ) );
  DFFPOSX1 \mem_reg<170>  ( .D(n1161), .CLK(clk), .Q(\mem<170> ) );
  DFFPOSX1 \mem_reg<171>  ( .D(n1162), .CLK(clk), .Q(\mem<171> ) );
  DFFPOSX1 \mem_reg<172>  ( .D(n1163), .CLK(clk), .Q(\mem<172> ) );
  DFFPOSX1 \mem_reg<173>  ( .D(n1164), .CLK(clk), .Q(\mem<173> ) );
  DFFPOSX1 \mem_reg<174>  ( .D(n1165), .CLK(clk), .Q(\mem<174> ) );
  DFFPOSX1 \mem_reg<175>  ( .D(n1166), .CLK(clk), .Q(\mem<175> ) );
  DFFPOSX1 \mem_reg<176>  ( .D(n1167), .CLK(clk), .Q(\mem<176> ) );
  DFFPOSX1 \mem_reg<177>  ( .D(n1168), .CLK(clk), .Q(\mem<177> ) );
  DFFPOSX1 \mem_reg<178>  ( .D(n1169), .CLK(clk), .Q(\mem<178> ) );
  DFFPOSX1 \mem_reg<179>  ( .D(n1170), .CLK(clk), .Q(\mem<179> ) );
  DFFPOSX1 \mem_reg<180>  ( .D(n1171), .CLK(clk), .Q(\mem<180> ) );
  DFFPOSX1 \mem_reg<181>  ( .D(n1172), .CLK(clk), .Q(\mem<181> ) );
  DFFPOSX1 \mem_reg<182>  ( .D(n1173), .CLK(clk), .Q(\mem<182> ) );
  DFFPOSX1 \mem_reg<183>  ( .D(n1174), .CLK(clk), .Q(\mem<183> ) );
  DFFPOSX1 \mem_reg<184>  ( .D(n1175), .CLK(clk), .Q(\mem<184> ) );
  DFFPOSX1 \mem_reg<185>  ( .D(n1176), .CLK(clk), .Q(\mem<185> ) );
  DFFPOSX1 \mem_reg<186>  ( .D(n1177), .CLK(clk), .Q(\mem<186> ) );
  DFFPOSX1 \mem_reg<187>  ( .D(n1178), .CLK(clk), .Q(\mem<187> ) );
  DFFPOSX1 \mem_reg<188>  ( .D(n1179), .CLK(clk), .Q(\mem<188> ) );
  DFFPOSX1 \mem_reg<189>  ( .D(n1180), .CLK(clk), .Q(\mem<189> ) );
  DFFPOSX1 \mem_reg<190>  ( .D(n1181), .CLK(clk), .Q(\mem<190> ) );
  DFFPOSX1 \mem_reg<191>  ( .D(n1182), .CLK(clk), .Q(\mem<191> ) );
  DFFPOSX1 \mem_reg<192>  ( .D(n1183), .CLK(clk), .Q(\mem<192> ) );
  DFFPOSX1 \mem_reg<193>  ( .D(n1184), .CLK(clk), .Q(\mem<193> ) );
  DFFPOSX1 \mem_reg<194>  ( .D(n1185), .CLK(clk), .Q(\mem<194> ) );
  DFFPOSX1 \mem_reg<195>  ( .D(n1186), .CLK(clk), .Q(\mem<195> ) );
  DFFPOSX1 \mem_reg<196>  ( .D(n1187), .CLK(clk), .Q(\mem<196> ) );
  DFFPOSX1 \mem_reg<197>  ( .D(n1188), .CLK(clk), .Q(\mem<197> ) );
  DFFPOSX1 \mem_reg<198>  ( .D(n1189), .CLK(clk), .Q(\mem<198> ) );
  DFFPOSX1 \mem_reg<199>  ( .D(n1190), .CLK(clk), .Q(\mem<199> ) );
  DFFPOSX1 \mem_reg<200>  ( .D(n1191), .CLK(clk), .Q(\mem<200> ) );
  DFFPOSX1 \mem_reg<201>  ( .D(n1192), .CLK(clk), .Q(\mem<201> ) );
  DFFPOSX1 \mem_reg<202>  ( .D(n1193), .CLK(clk), .Q(\mem<202> ) );
  DFFPOSX1 \mem_reg<203>  ( .D(n1194), .CLK(clk), .Q(\mem<203> ) );
  DFFPOSX1 \mem_reg<204>  ( .D(n1195), .CLK(clk), .Q(\mem<204> ) );
  DFFPOSX1 \mem_reg<205>  ( .D(n1196), .CLK(clk), .Q(\mem<205> ) );
  DFFPOSX1 \mem_reg<206>  ( .D(n1197), .CLK(clk), .Q(\mem<206> ) );
  DFFPOSX1 \mem_reg<207>  ( .D(n1198), .CLK(clk), .Q(\mem<207> ) );
  DFFPOSX1 \mem_reg<208>  ( .D(n1199), .CLK(clk), .Q(\mem<208> ) );
  DFFPOSX1 \mem_reg<209>  ( .D(n1200), .CLK(clk), .Q(\mem<209> ) );
  DFFPOSX1 \mem_reg<210>  ( .D(n1201), .CLK(clk), .Q(\mem<210> ) );
  DFFPOSX1 \mem_reg<211>  ( .D(n1202), .CLK(clk), .Q(\mem<211> ) );
  DFFPOSX1 \mem_reg<212>  ( .D(n1203), .CLK(clk), .Q(\mem<212> ) );
  DFFPOSX1 \mem_reg<213>  ( .D(n1204), .CLK(clk), .Q(\mem<213> ) );
  DFFPOSX1 \mem_reg<214>  ( .D(n1205), .CLK(clk), .Q(\mem<214> ) );
  DFFPOSX1 \mem_reg<215>  ( .D(n1206), .CLK(clk), .Q(\mem<215> ) );
  DFFPOSX1 \mem_reg<216>  ( .D(n1207), .CLK(clk), .Q(\mem<216> ) );
  DFFPOSX1 \mem_reg<217>  ( .D(n1208), .CLK(clk), .Q(\mem<217> ) );
  DFFPOSX1 \mem_reg<218>  ( .D(n1209), .CLK(clk), .Q(\mem<218> ) );
  DFFPOSX1 \mem_reg<219>  ( .D(n1210), .CLK(clk), .Q(\mem<219> ) );
  DFFPOSX1 \mem_reg<220>  ( .D(n1211), .CLK(clk), .Q(\mem<220> ) );
  DFFPOSX1 \mem_reg<221>  ( .D(n1212), .CLK(clk), .Q(\mem<221> ) );
  DFFPOSX1 \mem_reg<222>  ( .D(n1213), .CLK(clk), .Q(\mem<222> ) );
  DFFPOSX1 \mem_reg<223>  ( .D(n1214), .CLK(clk), .Q(\mem<223> ) );
  DFFPOSX1 \mem_reg<224>  ( .D(n1215), .CLK(clk), .Q(\mem<224> ) );
  DFFPOSX1 \mem_reg<225>  ( .D(n1216), .CLK(clk), .Q(\mem<225> ) );
  DFFPOSX1 \mem_reg<226>  ( .D(n1217), .CLK(clk), .Q(\mem<226> ) );
  DFFPOSX1 \mem_reg<227>  ( .D(n1218), .CLK(clk), .Q(\mem<227> ) );
  DFFPOSX1 \mem_reg<228>  ( .D(n1219), .CLK(clk), .Q(\mem<228> ) );
  DFFPOSX1 \mem_reg<229>  ( .D(n1220), .CLK(clk), .Q(\mem<229> ) );
  DFFPOSX1 \mem_reg<230>  ( .D(n1221), .CLK(clk), .Q(\mem<230> ) );
  DFFPOSX1 \mem_reg<231>  ( .D(n1222), .CLK(clk), .Q(\mem<231> ) );
  DFFPOSX1 \mem_reg<232>  ( .D(n1223), .CLK(clk), .Q(\mem<232> ) );
  DFFPOSX1 \mem_reg<233>  ( .D(n1224), .CLK(clk), .Q(\mem<233> ) );
  DFFPOSX1 \mem_reg<234>  ( .D(n1225), .CLK(clk), .Q(\mem<234> ) );
  DFFPOSX1 \mem_reg<235>  ( .D(n1226), .CLK(clk), .Q(\mem<235> ) );
  DFFPOSX1 \mem_reg<236>  ( .D(n1227), .CLK(clk), .Q(\mem<236> ) );
  DFFPOSX1 \mem_reg<237>  ( .D(n1228), .CLK(clk), .Q(\mem<237> ) );
  DFFPOSX1 \mem_reg<238>  ( .D(n1229), .CLK(clk), .Q(\mem<238> ) );
  DFFPOSX1 \mem_reg<239>  ( .D(n1230), .CLK(clk), .Q(\mem<239> ) );
  DFFPOSX1 \mem_reg<240>  ( .D(n1231), .CLK(clk), .Q(\mem<240> ) );
  DFFPOSX1 \mem_reg<241>  ( .D(n1232), .CLK(clk), .Q(\mem<241> ) );
  DFFPOSX1 \mem_reg<242>  ( .D(n1233), .CLK(clk), .Q(\mem<242> ) );
  DFFPOSX1 \mem_reg<243>  ( .D(n1234), .CLK(clk), .Q(\mem<243> ) );
  DFFPOSX1 \mem_reg<244>  ( .D(n1235), .CLK(clk), .Q(\mem<244> ) );
  DFFPOSX1 \mem_reg<245>  ( .D(n1236), .CLK(clk), .Q(\mem<245> ) );
  DFFPOSX1 \mem_reg<246>  ( .D(n1237), .CLK(clk), .Q(\mem<246> ) );
  DFFPOSX1 \mem_reg<247>  ( .D(n1238), .CLK(clk), .Q(\mem<247> ) );
  DFFPOSX1 \mem_reg<248>  ( .D(n1239), .CLK(clk), .Q(\mem<248> ) );
  DFFPOSX1 \mem_reg<249>  ( .D(n1240), .CLK(clk), .Q(\mem<249> ) );
  DFFPOSX1 \mem_reg<250>  ( .D(n1241), .CLK(clk), .Q(\mem<250> ) );
  DFFPOSX1 \mem_reg<251>  ( .D(n1242), .CLK(clk), .Q(\mem<251> ) );
  DFFPOSX1 \mem_reg<252>  ( .D(n1243), .CLK(clk), .Q(\mem<252> ) );
  DFFPOSX1 \mem_reg<253>  ( .D(n1244), .CLK(clk), .Q(\mem<253> ) );
  DFFPOSX1 \mem_reg<254>  ( .D(n1245), .CLK(clk), .Q(\mem<254> ) );
  DFFPOSX1 \mem_reg<255>  ( .D(n1246), .CLK(clk), .Q(\mem<255> ) );
  AND2X2 U6 ( .A(N21), .B(n984), .Y(n1265) );
  AND2X2 U7 ( .A(N21), .B(n985), .Y(n1258) );
  AND2X2 U8 ( .A(n982), .B(n980), .Y(n1264) );
  AND2X2 U9 ( .A(n982), .B(n981), .Y(n1262) );
  AND2X2 U10 ( .A(data_in), .B(n68), .Y(n1495) );
  OAI21X1 U49 ( .A(n958), .B(n636), .C(n1511), .Y(n1246) );
  OAI21X1 U50 ( .A(n37), .B(n978), .C(\mem<255> ), .Y(n1511) );
  OAI21X1 U51 ( .A(n636), .B(n955), .C(n1510), .Y(n1245) );
  OAI21X1 U52 ( .A(n979), .B(n35), .C(\mem<254> ), .Y(n1510) );
  OAI21X1 U53 ( .A(n636), .B(n954), .C(n1509), .Y(n1244) );
  OAI21X1 U54 ( .A(n979), .B(n33), .C(\mem<253> ), .Y(n1509) );
  OAI21X1 U55 ( .A(n636), .B(n953), .C(n1508), .Y(n1243) );
  OAI21X1 U56 ( .A(n979), .B(n31), .C(\mem<252> ), .Y(n1508) );
  OAI21X1 U57 ( .A(n636), .B(n951), .C(n1507), .Y(n1242) );
  OAI21X1 U58 ( .A(n979), .B(n29), .C(\mem<251> ), .Y(n1507) );
  OAI21X1 U59 ( .A(n636), .B(n949), .C(n1506), .Y(n1241) );
  OAI21X1 U60 ( .A(n979), .B(n27), .C(\mem<250> ), .Y(n1506) );
  OAI21X1 U61 ( .A(n636), .B(n947), .C(n1505), .Y(n1240) );
  OAI21X1 U62 ( .A(n979), .B(n25), .C(\mem<249> ), .Y(n1505) );
  OAI21X1 U63 ( .A(n636), .B(n945), .C(n1504), .Y(n1239) );
  OAI21X1 U64 ( .A(n979), .B(n23), .C(\mem<248> ), .Y(n1504) );
  OAI21X1 U65 ( .A(n636), .B(n944), .C(n1503), .Y(n1238) );
  OAI21X1 U66 ( .A(n979), .B(n21), .C(\mem<247> ), .Y(n1503) );
  OAI21X1 U67 ( .A(n636), .B(n943), .C(n1502), .Y(n1237) );
  OAI21X1 U68 ( .A(n978), .B(n19), .C(\mem<246> ), .Y(n1502) );
  OAI21X1 U69 ( .A(n636), .B(n942), .C(n1501), .Y(n1236) );
  OAI21X1 U70 ( .A(n978), .B(n17), .C(\mem<245> ), .Y(n1501) );
  OAI21X1 U71 ( .A(n636), .B(n941), .C(n1500), .Y(n1235) );
  OAI21X1 U72 ( .A(n978), .B(n15), .C(\mem<244> ), .Y(n1500) );
  OAI21X1 U73 ( .A(n636), .B(n940), .C(n1499), .Y(n1234) );
  OAI21X1 U74 ( .A(n978), .B(n13), .C(\mem<243> ), .Y(n1499) );
  OAI21X1 U75 ( .A(n636), .B(n939), .C(n1498), .Y(n1233) );
  OAI21X1 U76 ( .A(n978), .B(n11), .C(\mem<242> ), .Y(n1498) );
  OAI21X1 U77 ( .A(n636), .B(n938), .C(n1497), .Y(n1232) );
  OAI21X1 U78 ( .A(n978), .B(n9), .C(\mem<241> ), .Y(n1497) );
  OAI21X1 U79 ( .A(n636), .B(n936), .C(n1496), .Y(n1231) );
  OAI21X1 U80 ( .A(n978), .B(n7), .C(\mem<240> ), .Y(n1496) );
  OAI21X1 U83 ( .A(n958), .B(n369), .C(n1492), .Y(n1230) );
  OAI21X1 U84 ( .A(n37), .B(n977), .C(\mem<239> ), .Y(n1492) );
  OAI21X1 U85 ( .A(n956), .B(n369), .C(n1491), .Y(n1229) );
  OAI21X1 U86 ( .A(n35), .B(n977), .C(\mem<238> ), .Y(n1491) );
  OAI21X1 U87 ( .A(n954), .B(n369), .C(n1490), .Y(n1228) );
  OAI21X1 U88 ( .A(n33), .B(n977), .C(\mem<237> ), .Y(n1490) );
  OAI21X1 U89 ( .A(n953), .B(n369), .C(n1489), .Y(n1227) );
  OAI21X1 U90 ( .A(n31), .B(n977), .C(\mem<236> ), .Y(n1489) );
  OAI21X1 U91 ( .A(n952), .B(n369), .C(n1488), .Y(n1226) );
  OAI21X1 U92 ( .A(n29), .B(n977), .C(\mem<235> ), .Y(n1488) );
  OAI21X1 U93 ( .A(n950), .B(n369), .C(n1487), .Y(n1225) );
  OAI21X1 U94 ( .A(n27), .B(n977), .C(\mem<234> ), .Y(n1487) );
  OAI21X1 U95 ( .A(n948), .B(n369), .C(n1486), .Y(n1224) );
  OAI21X1 U96 ( .A(n25), .B(n977), .C(\mem<233> ), .Y(n1486) );
  OAI21X1 U97 ( .A(n946), .B(n369), .C(n1485), .Y(n1223) );
  OAI21X1 U98 ( .A(n23), .B(n977), .C(\mem<232> ), .Y(n1485) );
  OAI21X1 U99 ( .A(n944), .B(n369), .C(n1484), .Y(n1222) );
  OAI21X1 U100 ( .A(n21), .B(n976), .C(\mem<231> ), .Y(n1484) );
  OAI21X1 U101 ( .A(n943), .B(n369), .C(n1483), .Y(n1221) );
  OAI21X1 U102 ( .A(n19), .B(n976), .C(\mem<230> ), .Y(n1483) );
  OAI21X1 U103 ( .A(n942), .B(n369), .C(n1482), .Y(n1220) );
  OAI21X1 U104 ( .A(n17), .B(n976), .C(\mem<229> ), .Y(n1482) );
  OAI21X1 U105 ( .A(n941), .B(n369), .C(n1481), .Y(n1219) );
  OAI21X1 U106 ( .A(n15), .B(n976), .C(\mem<228> ), .Y(n1481) );
  OAI21X1 U107 ( .A(n940), .B(n369), .C(n1480), .Y(n1218) );
  OAI21X1 U108 ( .A(n13), .B(n976), .C(\mem<227> ), .Y(n1480) );
  OAI21X1 U109 ( .A(n939), .B(n369), .C(n1479), .Y(n1217) );
  OAI21X1 U110 ( .A(n11), .B(n976), .C(\mem<226> ), .Y(n1479) );
  OAI21X1 U111 ( .A(n938), .B(n369), .C(n1478), .Y(n1216) );
  OAI21X1 U112 ( .A(n9), .B(n976), .C(\mem<225> ), .Y(n1478) );
  OAI21X1 U113 ( .A(n936), .B(n369), .C(n1477), .Y(n1215) );
  OAI21X1 U114 ( .A(n7), .B(n976), .C(\mem<224> ), .Y(n1477) );
  OAI21X1 U117 ( .A(n958), .B(n353), .C(n1475), .Y(n1214) );
  OAI21X1 U118 ( .A(n37), .B(n975), .C(\mem<223> ), .Y(n1475) );
  OAI21X1 U119 ( .A(n956), .B(n353), .C(n1474), .Y(n1213) );
  OAI21X1 U120 ( .A(n35), .B(n975), .C(\mem<222> ), .Y(n1474) );
  OAI21X1 U121 ( .A(n954), .B(n353), .C(n1473), .Y(n1212) );
  OAI21X1 U122 ( .A(n33), .B(n975), .C(\mem<221> ), .Y(n1473) );
  OAI21X1 U123 ( .A(n953), .B(n353), .C(n1472), .Y(n1211) );
  OAI21X1 U124 ( .A(n31), .B(n975), .C(\mem<220> ), .Y(n1472) );
  OAI21X1 U125 ( .A(n952), .B(n353), .C(n1471), .Y(n1210) );
  OAI21X1 U126 ( .A(n29), .B(n975), .C(\mem<219> ), .Y(n1471) );
  OAI21X1 U127 ( .A(n950), .B(n353), .C(n1470), .Y(n1209) );
  OAI21X1 U128 ( .A(n27), .B(n975), .C(\mem<218> ), .Y(n1470) );
  OAI21X1 U129 ( .A(n948), .B(n353), .C(n1469), .Y(n1208) );
  OAI21X1 U130 ( .A(n25), .B(n975), .C(\mem<217> ), .Y(n1469) );
  OAI21X1 U131 ( .A(n946), .B(n353), .C(n1468), .Y(n1207) );
  OAI21X1 U132 ( .A(n23), .B(n975), .C(\mem<216> ), .Y(n1468) );
  OAI21X1 U133 ( .A(n944), .B(n353), .C(n1467), .Y(n1206) );
  OAI21X1 U134 ( .A(n21), .B(n975), .C(\mem<215> ), .Y(n1467) );
  OAI21X1 U135 ( .A(n943), .B(n353), .C(n1466), .Y(n1205) );
  OAI21X1 U136 ( .A(n19), .B(n975), .C(\mem<214> ), .Y(n1466) );
  OAI21X1 U137 ( .A(n942), .B(n353), .C(n1465), .Y(n1204) );
  OAI21X1 U138 ( .A(n17), .B(n975), .C(\mem<213> ), .Y(n1465) );
  OAI21X1 U139 ( .A(n941), .B(n353), .C(n1464), .Y(n1203) );
  OAI21X1 U140 ( .A(n15), .B(n975), .C(\mem<212> ), .Y(n1464) );
  OAI21X1 U141 ( .A(n940), .B(n353), .C(n1463), .Y(n1202) );
  OAI21X1 U142 ( .A(n13), .B(n975), .C(\mem<211> ), .Y(n1463) );
  OAI21X1 U143 ( .A(n939), .B(n353), .C(n1462), .Y(n1201) );
  OAI21X1 U144 ( .A(n11), .B(n975), .C(\mem<210> ), .Y(n1462) );
  OAI21X1 U145 ( .A(n938), .B(n353), .C(n1461), .Y(n1200) );
  OAI21X1 U146 ( .A(n9), .B(n975), .C(\mem<209> ), .Y(n1461) );
  OAI21X1 U147 ( .A(n936), .B(n353), .C(n1460), .Y(n1199) );
  OAI21X1 U148 ( .A(n7), .B(n975), .C(\mem<208> ), .Y(n1460) );
  OAI21X1 U151 ( .A(n958), .B(n335), .C(n1459), .Y(n1198) );
  OAI21X1 U152 ( .A(n37), .B(n974), .C(\mem<207> ), .Y(n1459) );
  OAI21X1 U153 ( .A(n956), .B(n335), .C(n1458), .Y(n1197) );
  OAI21X1 U154 ( .A(n35), .B(n974), .C(\mem<206> ), .Y(n1458) );
  OAI21X1 U155 ( .A(n954), .B(n335), .C(n1457), .Y(n1196) );
  OAI21X1 U156 ( .A(n33), .B(n974), .C(\mem<205> ), .Y(n1457) );
  OAI21X1 U157 ( .A(n953), .B(n335), .C(n1456), .Y(n1195) );
  OAI21X1 U158 ( .A(n31), .B(n974), .C(\mem<204> ), .Y(n1456) );
  OAI21X1 U159 ( .A(n952), .B(n335), .C(n1455), .Y(n1194) );
  OAI21X1 U160 ( .A(n29), .B(n974), .C(\mem<203> ), .Y(n1455) );
  OAI21X1 U161 ( .A(n950), .B(n335), .C(n1454), .Y(n1193) );
  OAI21X1 U162 ( .A(n27), .B(n974), .C(\mem<202> ), .Y(n1454) );
  OAI21X1 U163 ( .A(n948), .B(n335), .C(n1453), .Y(n1192) );
  OAI21X1 U164 ( .A(n25), .B(n974), .C(\mem<201> ), .Y(n1453) );
  OAI21X1 U165 ( .A(n946), .B(n335), .C(n1452), .Y(n1191) );
  OAI21X1 U166 ( .A(n23), .B(n974), .C(\mem<200> ), .Y(n1452) );
  OAI21X1 U167 ( .A(n944), .B(n335), .C(n1451), .Y(n1190) );
  OAI21X1 U168 ( .A(n21), .B(n974), .C(\mem<199> ), .Y(n1451) );
  OAI21X1 U169 ( .A(n943), .B(n335), .C(n1450), .Y(n1189) );
  OAI21X1 U170 ( .A(n19), .B(n974), .C(\mem<198> ), .Y(n1450) );
  OAI21X1 U171 ( .A(n942), .B(n335), .C(n1449), .Y(n1188) );
  OAI21X1 U172 ( .A(n17), .B(n974), .C(\mem<197> ), .Y(n1449) );
  OAI21X1 U173 ( .A(n941), .B(n335), .C(n1448), .Y(n1187) );
  OAI21X1 U174 ( .A(n15), .B(n974), .C(\mem<196> ), .Y(n1448) );
  OAI21X1 U175 ( .A(n940), .B(n335), .C(n1447), .Y(n1186) );
  OAI21X1 U176 ( .A(n13), .B(n974), .C(\mem<195> ), .Y(n1447) );
  OAI21X1 U177 ( .A(n939), .B(n335), .C(n1446), .Y(n1185) );
  OAI21X1 U178 ( .A(n11), .B(n974), .C(\mem<194> ), .Y(n1446) );
  OAI21X1 U179 ( .A(n938), .B(n335), .C(n1445), .Y(n1184) );
  OAI21X1 U180 ( .A(n9), .B(n974), .C(\mem<193> ), .Y(n1445) );
  OAI21X1 U181 ( .A(n936), .B(n335), .C(n1444), .Y(n1183) );
  OAI21X1 U182 ( .A(n7), .B(n974), .C(\mem<192> ), .Y(n1444) );
  OAI21X1 U185 ( .A(n958), .B(n317), .C(n1443), .Y(n1182) );
  OAI21X1 U186 ( .A(n37), .B(n973), .C(\mem<191> ), .Y(n1443) );
  OAI21X1 U187 ( .A(n956), .B(n317), .C(n1442), .Y(n1181) );
  OAI21X1 U188 ( .A(n35), .B(n973), .C(\mem<190> ), .Y(n1442) );
  OAI21X1 U189 ( .A(n954), .B(n317), .C(n1441), .Y(n1180) );
  OAI21X1 U190 ( .A(n33), .B(n973), .C(\mem<189> ), .Y(n1441) );
  OAI21X1 U191 ( .A(n953), .B(n317), .C(n1440), .Y(n1179) );
  OAI21X1 U192 ( .A(n31), .B(n973), .C(\mem<188> ), .Y(n1440) );
  OAI21X1 U193 ( .A(n952), .B(n317), .C(n1439), .Y(n1178) );
  OAI21X1 U194 ( .A(n29), .B(n973), .C(\mem<187> ), .Y(n1439) );
  OAI21X1 U195 ( .A(n950), .B(n317), .C(n1438), .Y(n1177) );
  OAI21X1 U196 ( .A(n27), .B(n973), .C(\mem<186> ), .Y(n1438) );
  OAI21X1 U197 ( .A(n948), .B(n317), .C(n1437), .Y(n1176) );
  OAI21X1 U198 ( .A(n25), .B(n973), .C(\mem<185> ), .Y(n1437) );
  OAI21X1 U199 ( .A(n946), .B(n317), .C(n1436), .Y(n1175) );
  OAI21X1 U200 ( .A(n23), .B(n973), .C(\mem<184> ), .Y(n1436) );
  OAI21X1 U201 ( .A(n944), .B(n317), .C(n1435), .Y(n1174) );
  OAI21X1 U202 ( .A(n21), .B(n972), .C(\mem<183> ), .Y(n1435) );
  OAI21X1 U203 ( .A(n943), .B(n317), .C(n1434), .Y(n1173) );
  OAI21X1 U204 ( .A(n19), .B(n972), .C(\mem<182> ), .Y(n1434) );
  OAI21X1 U205 ( .A(n942), .B(n317), .C(n1433), .Y(n1172) );
  OAI21X1 U206 ( .A(n17), .B(n972), .C(\mem<181> ), .Y(n1433) );
  OAI21X1 U207 ( .A(n941), .B(n317), .C(n1432), .Y(n1171) );
  OAI21X1 U208 ( .A(n15), .B(n972), .C(\mem<180> ), .Y(n1432) );
  OAI21X1 U209 ( .A(n940), .B(n317), .C(n1431), .Y(n1170) );
  OAI21X1 U210 ( .A(n13), .B(n972), .C(\mem<179> ), .Y(n1431) );
  OAI21X1 U211 ( .A(n939), .B(n317), .C(n1430), .Y(n1169) );
  OAI21X1 U212 ( .A(n11), .B(n972), .C(\mem<178> ), .Y(n1430) );
  OAI21X1 U213 ( .A(n938), .B(n317), .C(n1429), .Y(n1168) );
  OAI21X1 U214 ( .A(n9), .B(n972), .C(\mem<177> ), .Y(n1429) );
  OAI21X1 U215 ( .A(n936), .B(n317), .C(n1428), .Y(n1167) );
  OAI21X1 U216 ( .A(n7), .B(n972), .C(\mem<176> ), .Y(n1428) );
  OAI21X1 U219 ( .A(n958), .B(n296), .C(n1426), .Y(n1166) );
  OAI21X1 U220 ( .A(n37), .B(n971), .C(\mem<175> ), .Y(n1426) );
  OAI21X1 U221 ( .A(n956), .B(n296), .C(n1425), .Y(n1165) );
  OAI21X1 U222 ( .A(n35), .B(n971), .C(\mem<174> ), .Y(n1425) );
  OAI21X1 U223 ( .A(n954), .B(n296), .C(n1424), .Y(n1164) );
  OAI21X1 U224 ( .A(n33), .B(n971), .C(\mem<173> ), .Y(n1424) );
  OAI21X1 U225 ( .A(n953), .B(n296), .C(n1423), .Y(n1163) );
  OAI21X1 U226 ( .A(n31), .B(n971), .C(\mem<172> ), .Y(n1423) );
  OAI21X1 U227 ( .A(n952), .B(n296), .C(n1422), .Y(n1162) );
  OAI21X1 U228 ( .A(n29), .B(n971), .C(\mem<171> ), .Y(n1422) );
  OAI21X1 U229 ( .A(n950), .B(n296), .C(n1421), .Y(n1161) );
  OAI21X1 U230 ( .A(n27), .B(n971), .C(\mem<170> ), .Y(n1421) );
  OAI21X1 U231 ( .A(n948), .B(n296), .C(n1420), .Y(n1160) );
  OAI21X1 U232 ( .A(n25), .B(n971), .C(\mem<169> ), .Y(n1420) );
  OAI21X1 U233 ( .A(n946), .B(n296), .C(n1419), .Y(n1159) );
  OAI21X1 U234 ( .A(n23), .B(n971), .C(\mem<168> ), .Y(n1419) );
  OAI21X1 U235 ( .A(n944), .B(n296), .C(n1418), .Y(n1158) );
  OAI21X1 U236 ( .A(n21), .B(n970), .C(\mem<167> ), .Y(n1418) );
  OAI21X1 U237 ( .A(n943), .B(n296), .C(n1417), .Y(n1157) );
  OAI21X1 U238 ( .A(n19), .B(n970), .C(\mem<166> ), .Y(n1417) );
  OAI21X1 U239 ( .A(n942), .B(n296), .C(n1416), .Y(n1156) );
  OAI21X1 U240 ( .A(n17), .B(n970), .C(\mem<165> ), .Y(n1416) );
  OAI21X1 U241 ( .A(n941), .B(n296), .C(n1415), .Y(n1155) );
  OAI21X1 U242 ( .A(n15), .B(n970), .C(\mem<164> ), .Y(n1415) );
  OAI21X1 U243 ( .A(n940), .B(n296), .C(n1414), .Y(n1154) );
  OAI21X1 U244 ( .A(n13), .B(n970), .C(\mem<163> ), .Y(n1414) );
  OAI21X1 U245 ( .A(n939), .B(n296), .C(n1413), .Y(n1153) );
  OAI21X1 U246 ( .A(n11), .B(n970), .C(\mem<162> ), .Y(n1413) );
  OAI21X1 U247 ( .A(n938), .B(n296), .C(n1412), .Y(n1152) );
  OAI21X1 U248 ( .A(n9), .B(n970), .C(\mem<161> ), .Y(n1412) );
  OAI21X1 U249 ( .A(n936), .B(n296), .C(n1411), .Y(n1151) );
  OAI21X1 U250 ( .A(n7), .B(n970), .C(\mem<160> ), .Y(n1411) );
  OAI21X1 U253 ( .A(n958), .B(n260), .C(n1410), .Y(n1150) );
  OAI21X1 U254 ( .A(n37), .B(n969), .C(\mem<159> ), .Y(n1410) );
  OAI21X1 U255 ( .A(n956), .B(n260), .C(n1409), .Y(n1149) );
  OAI21X1 U256 ( .A(n35), .B(n969), .C(\mem<158> ), .Y(n1409) );
  OAI21X1 U257 ( .A(n954), .B(n260), .C(n1408), .Y(n1148) );
  OAI21X1 U258 ( .A(n33), .B(n969), .C(\mem<157> ), .Y(n1408) );
  OAI21X1 U259 ( .A(n953), .B(n260), .C(n1407), .Y(n1147) );
  OAI21X1 U260 ( .A(n31), .B(n969), .C(\mem<156> ), .Y(n1407) );
  OAI21X1 U261 ( .A(n952), .B(n260), .C(n1406), .Y(n1146) );
  OAI21X1 U262 ( .A(n29), .B(n969), .C(\mem<155> ), .Y(n1406) );
  OAI21X1 U263 ( .A(n950), .B(n260), .C(n1405), .Y(n1145) );
  OAI21X1 U264 ( .A(n27), .B(n969), .C(\mem<154> ), .Y(n1405) );
  OAI21X1 U265 ( .A(n948), .B(n260), .C(n1404), .Y(n1144) );
  OAI21X1 U266 ( .A(n25), .B(n969), .C(\mem<153> ), .Y(n1404) );
  OAI21X1 U267 ( .A(n946), .B(n260), .C(n1403), .Y(n1143) );
  OAI21X1 U268 ( .A(n23), .B(n969), .C(\mem<152> ), .Y(n1403) );
  OAI21X1 U269 ( .A(n944), .B(n260), .C(n1402), .Y(n1142) );
  OAI21X1 U270 ( .A(n21), .B(n968), .C(\mem<151> ), .Y(n1402) );
  OAI21X1 U271 ( .A(n943), .B(n260), .C(n1401), .Y(n1141) );
  OAI21X1 U272 ( .A(n19), .B(n968), .C(\mem<150> ), .Y(n1401) );
  OAI21X1 U273 ( .A(n942), .B(n260), .C(n1400), .Y(n1140) );
  OAI21X1 U274 ( .A(n17), .B(n968), .C(\mem<149> ), .Y(n1400) );
  OAI21X1 U275 ( .A(n941), .B(n260), .C(n1399), .Y(n1139) );
  OAI21X1 U276 ( .A(n15), .B(n968), .C(\mem<148> ), .Y(n1399) );
  OAI21X1 U277 ( .A(n940), .B(n260), .C(n1398), .Y(n1138) );
  OAI21X1 U278 ( .A(n13), .B(n968), .C(\mem<147> ), .Y(n1398) );
  OAI21X1 U279 ( .A(n939), .B(n260), .C(n1397), .Y(n1137) );
  OAI21X1 U280 ( .A(n11), .B(n968), .C(\mem<146> ), .Y(n1397) );
  OAI21X1 U281 ( .A(n938), .B(n260), .C(n1396), .Y(n1136) );
  OAI21X1 U282 ( .A(n9), .B(n968), .C(\mem<145> ), .Y(n1396) );
  OAI21X1 U283 ( .A(n936), .B(n260), .C(n1395), .Y(n1135) );
  OAI21X1 U284 ( .A(n7), .B(n968), .C(\mem<144> ), .Y(n1395) );
  OAI21X1 U287 ( .A(n958), .B(n225), .C(n1394), .Y(n1134) );
  OAI21X1 U288 ( .A(n37), .B(n967), .C(\mem<143> ), .Y(n1394) );
  OAI21X1 U289 ( .A(n956), .B(n225), .C(n1393), .Y(n1133) );
  OAI21X1 U290 ( .A(n35), .B(n967), .C(\mem<142> ), .Y(n1393) );
  OAI21X1 U291 ( .A(n954), .B(n225), .C(n1392), .Y(n1132) );
  OAI21X1 U292 ( .A(n33), .B(n967), .C(\mem<141> ), .Y(n1392) );
  OAI21X1 U293 ( .A(n953), .B(n225), .C(n1391), .Y(n1131) );
  OAI21X1 U294 ( .A(n31), .B(n967), .C(\mem<140> ), .Y(n1391) );
  OAI21X1 U295 ( .A(n952), .B(n225), .C(n1390), .Y(n1130) );
  OAI21X1 U296 ( .A(n29), .B(n967), .C(\mem<139> ), .Y(n1390) );
  OAI21X1 U297 ( .A(n950), .B(n225), .C(n1389), .Y(n1129) );
  OAI21X1 U298 ( .A(n27), .B(n967), .C(\mem<138> ), .Y(n1389) );
  OAI21X1 U299 ( .A(n948), .B(n225), .C(n1388), .Y(n1128) );
  OAI21X1 U300 ( .A(n25), .B(n967), .C(\mem<137> ), .Y(n1388) );
  OAI21X1 U301 ( .A(n946), .B(n225), .C(n1387), .Y(n1127) );
  OAI21X1 U302 ( .A(n23), .B(n967), .C(\mem<136> ), .Y(n1387) );
  OAI21X1 U303 ( .A(n944), .B(n225), .C(n1386), .Y(n1126) );
  OAI21X1 U304 ( .A(n21), .B(n966), .C(\mem<135> ), .Y(n1386) );
  OAI21X1 U305 ( .A(n943), .B(n225), .C(n1385), .Y(n1125) );
  OAI21X1 U306 ( .A(n19), .B(n966), .C(\mem<134> ), .Y(n1385) );
  OAI21X1 U307 ( .A(n942), .B(n225), .C(n1384), .Y(n1124) );
  OAI21X1 U308 ( .A(n17), .B(n966), .C(\mem<133> ), .Y(n1384) );
  OAI21X1 U309 ( .A(n941), .B(n225), .C(n1383), .Y(n1123) );
  OAI21X1 U310 ( .A(n15), .B(n966), .C(\mem<132> ), .Y(n1383) );
  OAI21X1 U311 ( .A(n940), .B(n225), .C(n1382), .Y(n1122) );
  OAI21X1 U312 ( .A(n13), .B(n966), .C(\mem<131> ), .Y(n1382) );
  OAI21X1 U313 ( .A(n939), .B(n225), .C(n1381), .Y(n1121) );
  OAI21X1 U314 ( .A(n11), .B(n966), .C(\mem<130> ), .Y(n1381) );
  OAI21X1 U315 ( .A(n938), .B(n225), .C(n1380), .Y(n1120) );
  OAI21X1 U316 ( .A(n9), .B(n966), .C(\mem<129> ), .Y(n1380) );
  OAI21X1 U317 ( .A(n936), .B(n225), .C(n1379), .Y(n1119) );
  OAI21X1 U318 ( .A(n7), .B(n966), .C(\mem<128> ), .Y(n1379) );
  OAI21X1 U321 ( .A(n957), .B(n189), .C(n1378), .Y(n1118) );
  OAI21X1 U322 ( .A(n37), .B(n965), .C(\mem<127> ), .Y(n1378) );
  OAI21X1 U323 ( .A(n956), .B(n189), .C(n1377), .Y(n1117) );
  OAI21X1 U324 ( .A(n35), .B(n965), .C(\mem<126> ), .Y(n1377) );
  OAI21X1 U325 ( .A(n954), .B(n189), .C(n1376), .Y(n1116) );
  OAI21X1 U326 ( .A(n33), .B(n965), .C(\mem<125> ), .Y(n1376) );
  OAI21X1 U327 ( .A(n953), .B(n189), .C(n1375), .Y(n1115) );
  OAI21X1 U328 ( .A(n31), .B(n965), .C(\mem<124> ), .Y(n1375) );
  OAI21X1 U329 ( .A(n952), .B(n189), .C(n1374), .Y(n1114) );
  OAI21X1 U330 ( .A(n29), .B(n965), .C(\mem<123> ), .Y(n1374) );
  OAI21X1 U331 ( .A(n950), .B(n189), .C(n1373), .Y(n1113) );
  OAI21X1 U332 ( .A(n27), .B(n965), .C(\mem<122> ), .Y(n1373) );
  OAI21X1 U333 ( .A(n948), .B(n189), .C(n1372), .Y(n1112) );
  OAI21X1 U334 ( .A(n25), .B(n965), .C(\mem<121> ), .Y(n1372) );
  OAI21X1 U335 ( .A(n946), .B(n189), .C(n1371), .Y(n1111) );
  OAI21X1 U336 ( .A(n23), .B(n965), .C(\mem<120> ), .Y(n1371) );
  OAI21X1 U337 ( .A(n944), .B(n189), .C(n1370), .Y(n1110) );
  OAI21X1 U338 ( .A(n21), .B(n965), .C(\mem<119> ), .Y(n1370) );
  OAI21X1 U339 ( .A(n943), .B(n189), .C(n1369), .Y(n1109) );
  OAI21X1 U340 ( .A(n19), .B(n965), .C(\mem<118> ), .Y(n1369) );
  OAI21X1 U341 ( .A(n942), .B(n189), .C(n1368), .Y(n1108) );
  OAI21X1 U342 ( .A(n17), .B(n965), .C(\mem<117> ), .Y(n1368) );
  OAI21X1 U343 ( .A(n941), .B(n189), .C(n1367), .Y(n1107) );
  OAI21X1 U344 ( .A(n15), .B(n965), .C(\mem<116> ), .Y(n1367) );
  OAI21X1 U345 ( .A(n940), .B(n189), .C(n1366), .Y(n1106) );
  OAI21X1 U346 ( .A(n13), .B(n965), .C(\mem<115> ), .Y(n1366) );
  OAI21X1 U347 ( .A(n939), .B(n189), .C(n1365), .Y(n1105) );
  OAI21X1 U348 ( .A(n11), .B(n965), .C(\mem<114> ), .Y(n1365) );
  OAI21X1 U349 ( .A(n938), .B(n189), .C(n1364), .Y(n1104) );
  OAI21X1 U350 ( .A(n9), .B(n965), .C(\mem<113> ), .Y(n1364) );
  OAI21X1 U351 ( .A(n936), .B(n189), .C(n1363), .Y(n1103) );
  OAI21X1 U352 ( .A(n7), .B(n965), .C(\mem<112> ), .Y(n1363) );
  OAI21X1 U355 ( .A(n957), .B(n171), .C(n1362), .Y(n1102) );
  OAI21X1 U356 ( .A(n37), .B(n964), .C(\mem<111> ), .Y(n1362) );
  OAI21X1 U357 ( .A(n955), .B(n171), .C(n1361), .Y(n1101) );
  OAI21X1 U358 ( .A(n35), .B(n964), .C(\mem<110> ), .Y(n1361) );
  OAI21X1 U359 ( .A(n954), .B(n171), .C(n1360), .Y(n1100) );
  OAI21X1 U360 ( .A(n33), .B(n964), .C(\mem<109> ), .Y(n1360) );
  OAI21X1 U361 ( .A(n953), .B(n171), .C(n1359), .Y(n1099) );
  OAI21X1 U362 ( .A(n31), .B(n964), .C(\mem<108> ), .Y(n1359) );
  OAI21X1 U363 ( .A(n951), .B(n171), .C(n1358), .Y(n1098) );
  OAI21X1 U364 ( .A(n29), .B(n964), .C(\mem<107> ), .Y(n1358) );
  OAI21X1 U365 ( .A(n949), .B(n171), .C(n1357), .Y(n1097) );
  OAI21X1 U366 ( .A(n27), .B(n964), .C(\mem<106> ), .Y(n1357) );
  OAI21X1 U367 ( .A(n947), .B(n171), .C(n1356), .Y(n1096) );
  OAI21X1 U368 ( .A(n25), .B(n964), .C(\mem<105> ), .Y(n1356) );
  OAI21X1 U369 ( .A(n945), .B(n171), .C(n1355), .Y(n1095) );
  OAI21X1 U370 ( .A(n23), .B(n964), .C(\mem<104> ), .Y(n1355) );
  OAI21X1 U371 ( .A(n944), .B(n171), .C(n1354), .Y(n1094) );
  OAI21X1 U372 ( .A(n21), .B(n964), .C(\mem<103> ), .Y(n1354) );
  OAI21X1 U373 ( .A(n943), .B(n171), .C(n1353), .Y(n1093) );
  OAI21X1 U374 ( .A(n19), .B(n964), .C(\mem<102> ), .Y(n1353) );
  OAI21X1 U375 ( .A(n942), .B(n171), .C(n1352), .Y(n1092) );
  OAI21X1 U376 ( .A(n17), .B(n964), .C(\mem<101> ), .Y(n1352) );
  OAI21X1 U377 ( .A(n941), .B(n171), .C(n1351), .Y(n1091) );
  OAI21X1 U378 ( .A(n15), .B(n964), .C(\mem<100> ), .Y(n1351) );
  OAI21X1 U379 ( .A(n940), .B(n171), .C(n1350), .Y(n1090) );
  OAI21X1 U380 ( .A(n13), .B(n964), .C(\mem<99> ), .Y(n1350) );
  OAI21X1 U381 ( .A(n939), .B(n171), .C(n1349), .Y(n1089) );
  OAI21X1 U382 ( .A(n11), .B(n964), .C(\mem<98> ), .Y(n1349) );
  OAI21X1 U383 ( .A(n938), .B(n171), .C(n1348), .Y(n1088) );
  OAI21X1 U384 ( .A(n9), .B(n964), .C(\mem<97> ), .Y(n1348) );
  OAI21X1 U385 ( .A(n936), .B(n171), .C(n1347), .Y(n1087) );
  OAI21X1 U386 ( .A(n7), .B(n964), .C(\mem<96> ), .Y(n1347) );
  OAI21X1 U389 ( .A(n957), .B(n152), .C(n1346), .Y(n1086) );
  OAI21X1 U390 ( .A(n37), .B(n963), .C(\mem<95> ), .Y(n1346) );
  OAI21X1 U391 ( .A(n955), .B(n152), .C(n1345), .Y(n1085) );
  OAI21X1 U392 ( .A(n35), .B(n963), .C(\mem<94> ), .Y(n1345) );
  OAI21X1 U393 ( .A(n954), .B(n152), .C(n1344), .Y(n1084) );
  OAI21X1 U394 ( .A(n33), .B(n963), .C(\mem<93> ), .Y(n1344) );
  OAI21X1 U395 ( .A(n953), .B(n152), .C(n1343), .Y(n1083) );
  OAI21X1 U396 ( .A(n31), .B(n963), .C(\mem<92> ), .Y(n1343) );
  OAI21X1 U397 ( .A(n951), .B(n152), .C(n1342), .Y(n1082) );
  OAI21X1 U398 ( .A(n29), .B(n963), .C(\mem<91> ), .Y(n1342) );
  OAI21X1 U399 ( .A(n949), .B(n152), .C(n1341), .Y(n1081) );
  OAI21X1 U400 ( .A(n27), .B(n963), .C(\mem<90> ), .Y(n1341) );
  OAI21X1 U401 ( .A(n947), .B(n152), .C(n1340), .Y(n1080) );
  OAI21X1 U402 ( .A(n25), .B(n963), .C(\mem<89> ), .Y(n1340) );
  OAI21X1 U403 ( .A(n945), .B(n152), .C(n1339), .Y(n1079) );
  OAI21X1 U404 ( .A(n23), .B(n963), .C(\mem<88> ), .Y(n1339) );
  OAI21X1 U405 ( .A(n944), .B(n152), .C(n1338), .Y(n1078) );
  OAI21X1 U406 ( .A(n21), .B(n963), .C(\mem<87> ), .Y(n1338) );
  OAI21X1 U407 ( .A(n943), .B(n152), .C(n1337), .Y(n1077) );
  OAI21X1 U408 ( .A(n19), .B(n963), .C(\mem<86> ), .Y(n1337) );
  OAI21X1 U409 ( .A(n942), .B(n152), .C(n1336), .Y(n1076) );
  OAI21X1 U410 ( .A(n17), .B(n963), .C(\mem<85> ), .Y(n1336) );
  OAI21X1 U411 ( .A(n941), .B(n152), .C(n1335), .Y(n1075) );
  OAI21X1 U412 ( .A(n15), .B(n963), .C(\mem<84> ), .Y(n1335) );
  OAI21X1 U413 ( .A(n940), .B(n152), .C(n1334), .Y(n1074) );
  OAI21X1 U414 ( .A(n13), .B(n963), .C(\mem<83> ), .Y(n1334) );
  OAI21X1 U415 ( .A(n939), .B(n152), .C(n1333), .Y(n1073) );
  OAI21X1 U416 ( .A(n11), .B(n963), .C(\mem<82> ), .Y(n1333) );
  OAI21X1 U417 ( .A(n938), .B(n152), .C(n1332), .Y(n1072) );
  OAI21X1 U418 ( .A(n9), .B(n963), .C(\mem<81> ), .Y(n1332) );
  OAI21X1 U419 ( .A(n936), .B(n152), .C(n1331), .Y(n1071) );
  OAI21X1 U420 ( .A(n7), .B(n963), .C(\mem<80> ), .Y(n1331) );
  OAI21X1 U423 ( .A(n957), .B(n149), .C(n1330), .Y(n1070) );
  OAI21X1 U424 ( .A(n37), .B(n962), .C(\mem<79> ), .Y(n1330) );
  OAI21X1 U425 ( .A(n955), .B(n149), .C(n1329), .Y(n1069) );
  OAI21X1 U426 ( .A(n35), .B(n962), .C(\mem<78> ), .Y(n1329) );
  OAI21X1 U427 ( .A(n954), .B(n149), .C(n1328), .Y(n1068) );
  OAI21X1 U428 ( .A(n33), .B(n962), .C(\mem<77> ), .Y(n1328) );
  OAI21X1 U429 ( .A(n953), .B(n149), .C(n1327), .Y(n1067) );
  OAI21X1 U430 ( .A(n31), .B(n962), .C(\mem<76> ), .Y(n1327) );
  OAI21X1 U431 ( .A(n951), .B(n149), .C(n1326), .Y(n1066) );
  OAI21X1 U432 ( .A(n29), .B(n962), .C(\mem<75> ), .Y(n1326) );
  OAI21X1 U433 ( .A(n949), .B(n149), .C(n1325), .Y(n1065) );
  OAI21X1 U434 ( .A(n27), .B(n962), .C(\mem<74> ), .Y(n1325) );
  OAI21X1 U435 ( .A(n947), .B(n149), .C(n1324), .Y(n1064) );
  OAI21X1 U436 ( .A(n25), .B(n962), .C(\mem<73> ), .Y(n1324) );
  OAI21X1 U437 ( .A(n945), .B(n149), .C(n1323), .Y(n1063) );
  OAI21X1 U438 ( .A(n23), .B(n962), .C(\mem<72> ), .Y(n1323) );
  OAI21X1 U439 ( .A(n944), .B(n149), .C(n1322), .Y(n1062) );
  OAI21X1 U440 ( .A(n21), .B(n962), .C(\mem<71> ), .Y(n1322) );
  OAI21X1 U441 ( .A(n943), .B(n149), .C(n1321), .Y(n1061) );
  OAI21X1 U442 ( .A(n19), .B(n962), .C(\mem<70> ), .Y(n1321) );
  OAI21X1 U443 ( .A(n942), .B(n149), .C(n1320), .Y(n1060) );
  OAI21X1 U444 ( .A(n17), .B(n962), .C(\mem<69> ), .Y(n1320) );
  OAI21X1 U445 ( .A(n941), .B(n149), .C(n1319), .Y(n1059) );
  OAI21X1 U446 ( .A(n15), .B(n962), .C(\mem<68> ), .Y(n1319) );
  OAI21X1 U447 ( .A(n940), .B(n149), .C(n1318), .Y(n1058) );
  OAI21X1 U448 ( .A(n13), .B(n962), .C(\mem<67> ), .Y(n1318) );
  OAI21X1 U449 ( .A(n939), .B(n149), .C(n1317), .Y(n1057) );
  OAI21X1 U450 ( .A(n11), .B(n962), .C(\mem<66> ), .Y(n1317) );
  OAI21X1 U451 ( .A(n938), .B(n149), .C(n1316), .Y(n1056) );
  OAI21X1 U452 ( .A(n9), .B(n962), .C(\mem<65> ), .Y(n1316) );
  OAI21X1 U453 ( .A(n936), .B(n149), .C(n1315), .Y(n1055) );
  OAI21X1 U454 ( .A(n7), .B(n962), .C(\mem<64> ), .Y(n1315) );
  OAI21X1 U458 ( .A(n957), .B(n131), .C(n1314), .Y(n1054) );
  OAI21X1 U459 ( .A(n37), .B(n961), .C(\mem<63> ), .Y(n1314) );
  OAI21X1 U460 ( .A(n955), .B(n131), .C(n1313), .Y(n1053) );
  OAI21X1 U461 ( .A(n35), .B(n961), .C(\mem<62> ), .Y(n1313) );
  OAI21X1 U462 ( .A(n954), .B(n131), .C(n1312), .Y(n1052) );
  OAI21X1 U463 ( .A(n33), .B(n961), .C(\mem<61> ), .Y(n1312) );
  OAI21X1 U464 ( .A(n953), .B(n131), .C(n1311), .Y(n1051) );
  OAI21X1 U465 ( .A(n31), .B(n961), .C(\mem<60> ), .Y(n1311) );
  OAI21X1 U466 ( .A(n951), .B(n131), .C(n1310), .Y(n1050) );
  OAI21X1 U467 ( .A(n29), .B(n961), .C(\mem<59> ), .Y(n1310) );
  OAI21X1 U468 ( .A(n949), .B(n131), .C(n1309), .Y(n1049) );
  OAI21X1 U469 ( .A(n27), .B(n961), .C(\mem<58> ), .Y(n1309) );
  OAI21X1 U470 ( .A(n947), .B(n131), .C(n1308), .Y(n1048) );
  OAI21X1 U471 ( .A(n25), .B(n961), .C(\mem<57> ), .Y(n1308) );
  OAI21X1 U472 ( .A(n945), .B(n131), .C(n1307), .Y(n1047) );
  OAI21X1 U473 ( .A(n23), .B(n961), .C(\mem<56> ), .Y(n1307) );
  OAI21X1 U474 ( .A(n944), .B(n131), .C(n1306), .Y(n1046) );
  OAI21X1 U475 ( .A(n21), .B(n961), .C(\mem<55> ), .Y(n1306) );
  OAI21X1 U476 ( .A(n943), .B(n131), .C(n1305), .Y(n1045) );
  OAI21X1 U477 ( .A(n19), .B(n961), .C(\mem<54> ), .Y(n1305) );
  OAI21X1 U478 ( .A(n942), .B(n131), .C(n1304), .Y(n1044) );
  OAI21X1 U479 ( .A(n17), .B(n961), .C(\mem<53> ), .Y(n1304) );
  OAI21X1 U480 ( .A(n941), .B(n131), .C(n1303), .Y(n1043) );
  OAI21X1 U481 ( .A(n15), .B(n961), .C(\mem<52> ), .Y(n1303) );
  OAI21X1 U482 ( .A(n940), .B(n131), .C(n1302), .Y(n1042) );
  OAI21X1 U483 ( .A(n13), .B(n961), .C(\mem<51> ), .Y(n1302) );
  OAI21X1 U484 ( .A(n939), .B(n131), .C(n1301), .Y(n1041) );
  OAI21X1 U485 ( .A(n11), .B(n961), .C(\mem<50> ), .Y(n1301) );
  OAI21X1 U486 ( .A(n938), .B(n131), .C(n1300), .Y(n1040) );
  OAI21X1 U487 ( .A(n9), .B(n961), .C(\mem<49> ), .Y(n1300) );
  OAI21X1 U488 ( .A(n936), .B(n131), .C(n1299), .Y(n1039) );
  OAI21X1 U489 ( .A(n7), .B(n961), .C(\mem<48> ), .Y(n1299) );
  OAI21X1 U492 ( .A(n957), .B(n114), .C(n1298), .Y(n1038) );
  OAI21X1 U493 ( .A(n37), .B(n960), .C(\mem<47> ), .Y(n1298) );
  OAI21X1 U494 ( .A(n955), .B(n114), .C(n1297), .Y(n1037) );
  OAI21X1 U495 ( .A(n35), .B(n960), .C(\mem<46> ), .Y(n1297) );
  OAI21X1 U496 ( .A(n954), .B(n114), .C(n1296), .Y(n1036) );
  OAI21X1 U497 ( .A(n33), .B(n960), .C(\mem<45> ), .Y(n1296) );
  OAI21X1 U498 ( .A(n953), .B(n114), .C(n1295), .Y(n1035) );
  OAI21X1 U499 ( .A(n31), .B(n960), .C(\mem<44> ), .Y(n1295) );
  OAI21X1 U500 ( .A(n951), .B(n114), .C(n1294), .Y(n1034) );
  OAI21X1 U501 ( .A(n29), .B(n960), .C(\mem<43> ), .Y(n1294) );
  OAI21X1 U502 ( .A(n949), .B(n114), .C(n1293), .Y(n1033) );
  OAI21X1 U503 ( .A(n27), .B(n960), .C(\mem<42> ), .Y(n1293) );
  OAI21X1 U504 ( .A(n947), .B(n114), .C(n1292), .Y(n1032) );
  OAI21X1 U505 ( .A(n25), .B(n960), .C(\mem<41> ), .Y(n1292) );
  OAI21X1 U506 ( .A(n945), .B(n114), .C(n1291), .Y(n1031) );
  OAI21X1 U507 ( .A(n23), .B(n960), .C(\mem<40> ), .Y(n1291) );
  OAI21X1 U508 ( .A(n944), .B(n114), .C(n1290), .Y(n1030) );
  OAI21X1 U509 ( .A(n21), .B(n960), .C(\mem<39> ), .Y(n1290) );
  OAI21X1 U510 ( .A(n943), .B(n114), .C(n1289), .Y(n1029) );
  OAI21X1 U511 ( .A(n19), .B(n960), .C(\mem<38> ), .Y(n1289) );
  OAI21X1 U512 ( .A(n942), .B(n114), .C(n1288), .Y(n1028) );
  OAI21X1 U513 ( .A(n17), .B(n960), .C(\mem<37> ), .Y(n1288) );
  OAI21X1 U514 ( .A(n941), .B(n114), .C(n1287), .Y(n1027) );
  OAI21X1 U515 ( .A(n15), .B(n960), .C(\mem<36> ), .Y(n1287) );
  OAI21X1 U516 ( .A(n940), .B(n114), .C(n1286), .Y(n1026) );
  OAI21X1 U517 ( .A(n13), .B(n960), .C(\mem<35> ), .Y(n1286) );
  OAI21X1 U518 ( .A(n939), .B(n114), .C(n1285), .Y(n1025) );
  OAI21X1 U519 ( .A(n11), .B(n960), .C(\mem<34> ), .Y(n1285) );
  OAI21X1 U520 ( .A(n938), .B(n114), .C(n1284), .Y(n1024) );
  OAI21X1 U521 ( .A(n9), .B(n960), .C(\mem<33> ), .Y(n1284) );
  OAI21X1 U522 ( .A(n936), .B(n114), .C(n1283), .Y(n1023) );
  OAI21X1 U523 ( .A(n7), .B(n960), .C(\mem<32> ), .Y(n1283) );
  OAI21X1 U526 ( .A(n957), .B(n95), .C(n1282), .Y(n1022) );
  OAI21X1 U527 ( .A(n37), .B(n959), .C(\mem<31> ), .Y(n1282) );
  OAI21X1 U528 ( .A(n955), .B(n95), .C(n1281), .Y(n1021) );
  OAI21X1 U529 ( .A(n35), .B(n959), .C(\mem<30> ), .Y(n1281) );
  OAI21X1 U530 ( .A(n954), .B(n95), .C(n1280), .Y(n1020) );
  OAI21X1 U531 ( .A(n33), .B(n959), .C(\mem<29> ), .Y(n1280) );
  OAI21X1 U532 ( .A(n953), .B(n95), .C(n1279), .Y(n1019) );
  OAI21X1 U533 ( .A(n31), .B(n959), .C(\mem<28> ), .Y(n1279) );
  OAI21X1 U534 ( .A(n951), .B(n95), .C(n1278), .Y(n1018) );
  OAI21X1 U535 ( .A(n29), .B(n959), .C(\mem<27> ), .Y(n1278) );
  OAI21X1 U536 ( .A(n949), .B(n95), .C(n1277), .Y(n1017) );
  OAI21X1 U537 ( .A(n27), .B(n959), .C(\mem<26> ), .Y(n1277) );
  OAI21X1 U538 ( .A(n947), .B(n95), .C(n1276), .Y(n1016) );
  OAI21X1 U539 ( .A(n25), .B(n959), .C(\mem<25> ), .Y(n1276) );
  OAI21X1 U540 ( .A(n945), .B(n95), .C(n1275), .Y(n1015) );
  OAI21X1 U541 ( .A(n23), .B(n959), .C(\mem<24> ), .Y(n1275) );
  OAI21X1 U542 ( .A(n944), .B(n95), .C(n1274), .Y(n1014) );
  OAI21X1 U543 ( .A(n21), .B(n959), .C(\mem<23> ), .Y(n1274) );
  OAI21X1 U544 ( .A(n943), .B(n95), .C(n1273), .Y(n1013) );
  OAI21X1 U545 ( .A(n19), .B(n959), .C(\mem<22> ), .Y(n1273) );
  OAI21X1 U546 ( .A(n942), .B(n95), .C(n1272), .Y(n1012) );
  OAI21X1 U547 ( .A(n17), .B(n959), .C(\mem<21> ), .Y(n1272) );
  OAI21X1 U548 ( .A(n941), .B(n95), .C(n1271), .Y(n1011) );
  OAI21X1 U549 ( .A(n15), .B(n959), .C(\mem<20> ), .Y(n1271) );
  OAI21X1 U550 ( .A(n940), .B(n95), .C(n1270), .Y(n1010) );
  OAI21X1 U551 ( .A(n13), .B(n959), .C(\mem<19> ), .Y(n1270) );
  OAI21X1 U552 ( .A(n939), .B(n95), .C(n1269), .Y(n1009) );
  OAI21X1 U553 ( .A(n11), .B(n959), .C(\mem<18> ), .Y(n1269) );
  OAI21X1 U554 ( .A(n938), .B(n95), .C(n1268), .Y(n1008) );
  OAI21X1 U555 ( .A(n9), .B(n959), .C(\mem<17> ), .Y(n1268) );
  OAI21X1 U556 ( .A(n936), .B(n95), .C(n1267), .Y(n1007) );
  OAI21X1 U557 ( .A(n7), .B(n959), .C(\mem<16> ), .Y(n1267) );
  OAI21X1 U561 ( .A(n957), .B(n71), .C(n1266), .Y(n1006) );
  OAI21X1 U562 ( .A(n37), .B(n937), .C(\mem<15> ), .Y(n1266) );
  OAI21X1 U565 ( .A(n955), .B(n71), .C(n1263), .Y(n1005) );
  OAI21X1 U566 ( .A(n35), .B(n937), .C(\mem<14> ), .Y(n1263) );
  OAI21X1 U569 ( .A(n954), .B(n71), .C(n1261), .Y(n1004) );
  OAI21X1 U570 ( .A(n33), .B(n937), .C(\mem<13> ), .Y(n1261) );
  OAI21X1 U573 ( .A(n953), .B(n71), .C(n1260), .Y(n1003) );
  OAI21X1 U574 ( .A(n31), .B(n937), .C(\mem<12> ), .Y(n1260) );
  OAI21X1 U577 ( .A(n951), .B(n71), .C(n1259), .Y(n1002) );
  OAI21X1 U578 ( .A(n29), .B(n937), .C(\mem<11> ), .Y(n1259) );
  OAI21X1 U581 ( .A(n949), .B(n71), .C(n1257), .Y(n1001) );
  OAI21X1 U582 ( .A(n27), .B(n937), .C(\mem<10> ), .Y(n1257) );
  OAI21X1 U585 ( .A(n947), .B(n71), .C(n1256), .Y(n1000) );
  OAI21X1 U586 ( .A(n25), .B(n937), .C(\mem<9> ), .Y(n1256) );
  OAI21X1 U589 ( .A(n945), .B(n71), .C(n1255), .Y(n999) );
  OAI21X1 U590 ( .A(n23), .B(n937), .C(\mem<8> ), .Y(n1255) );
  OAI21X1 U593 ( .A(n944), .B(n71), .C(n1254), .Y(n998) );
  OAI21X1 U594 ( .A(n21), .B(n937), .C(\mem<7> ), .Y(n1254) );
  OAI21X1 U597 ( .A(n943), .B(n71), .C(n1253), .Y(n997) );
  OAI21X1 U598 ( .A(n19), .B(n937), .C(\mem<6> ), .Y(n1253) );
  OAI21X1 U601 ( .A(n942), .B(n71), .C(n1252), .Y(n996) );
  OAI21X1 U602 ( .A(n17), .B(n937), .C(\mem<5> ), .Y(n1252) );
  OAI21X1 U605 ( .A(n941), .B(n71), .C(n1251), .Y(n995) );
  OAI21X1 U606 ( .A(n15), .B(n937), .C(\mem<4> ), .Y(n1251) );
  OAI21X1 U610 ( .A(n940), .B(n71), .C(n1250), .Y(n994) );
  OAI21X1 U611 ( .A(n13), .B(n937), .C(\mem<3> ), .Y(n1250) );
  OAI21X1 U614 ( .A(n939), .B(n71), .C(n1249), .Y(n993) );
  OAI21X1 U615 ( .A(n11), .B(n937), .C(\mem<2> ), .Y(n1249) );
  OAI21X1 U618 ( .A(n938), .B(n71), .C(n1248), .Y(n992) );
  OAI21X1 U619 ( .A(n9), .B(n937), .C(\mem<1> ), .Y(n1248) );
  OAI21X1 U623 ( .A(n936), .B(n71), .C(n1247), .Y(n991) );
  OAI21X1 U624 ( .A(n7), .B(n937), .C(\mem<0> ), .Y(n1247) );
  INVX2 U2 ( .A(n66), .Y(n68) );
  INVX2 U3 ( .A(n187), .Y(n189) );
  INVX2 U4 ( .A(N21), .Y(n907) );
  INVX2 U5 ( .A(n907), .Y(n908) );
  AND2X1 U11 ( .A(N25), .B(n988), .Y(n1427) );
  INVX1 U12 ( .A(N22), .Y(n987) );
  AND2X1 U13 ( .A(N25), .B(N24), .Y(n1494) );
  AND2X1 U14 ( .A(N23), .B(n986), .Y(n1493) );
  AND2X1 U15 ( .A(N23), .B(n987), .Y(n1476) );
  BUFX2 U16 ( .A(n634), .Y(n978) );
  BUFX2 U17 ( .A(n360), .Y(n976) );
  BUFX2 U18 ( .A(n314), .Y(n972) );
  BUFX2 U19 ( .A(n278), .Y(n970) );
  BUFX2 U20 ( .A(n242), .Y(n968) );
  BUFX2 U21 ( .A(n207), .Y(n966) );
  BUFX2 U22 ( .A(n89), .Y(n957) );
  BUFX2 U23 ( .A(n86), .Y(n955) );
  BUFX2 U24 ( .A(n83), .Y(n951) );
  BUFX2 U25 ( .A(n80), .Y(n949) );
  BUFX2 U26 ( .A(n77), .Y(n947) );
  BUFX2 U27 ( .A(n74), .Y(n945) );
  INVX1 U28 ( .A(n935), .Y(n921) );
  INVX2 U29 ( .A(n987), .Y(n986) );
  INVX1 U30 ( .A(n39), .Y(n937) );
  INVX1 U31 ( .A(n53), .Y(n959) );
  INVX1 U32 ( .A(n54), .Y(n960) );
  INVX1 U33 ( .A(n56), .Y(n961) );
  INVX4 U34 ( .A(n980), .Y(n934) );
  INVX1 U35 ( .A(n57), .Y(n962) );
  INVX1 U36 ( .A(n59), .Y(n963) );
  INVX1 U37 ( .A(n60), .Y(n964) );
  INVX1 U38 ( .A(n62), .Y(n965) );
  INVX1 U39 ( .A(n63), .Y(n974) );
  INVX1 U40 ( .A(n65), .Y(n975) );
  INVX1 U41 ( .A(n50), .Y(n953) );
  INVX1 U42 ( .A(n51), .Y(n954) );
  BUFX2 U43 ( .A(n83), .Y(n952) );
  BUFX2 U44 ( .A(n86), .Y(n956) );
  BUFX2 U45 ( .A(n89), .Y(n958) );
  BUFX2 U46 ( .A(n74), .Y(n946) );
  INVX1 U47 ( .A(n985), .Y(n984) );
  BUFX2 U48 ( .A(n207), .Y(n967) );
  BUFX2 U81 ( .A(n242), .Y(n969) );
  BUFX2 U82 ( .A(n278), .Y(n971) );
  BUFX2 U115 ( .A(n314), .Y(n973) );
  BUFX2 U116 ( .A(n360), .Y(n977) );
  BUFX2 U149 ( .A(n634), .Y(n979) );
  BUFX2 U150 ( .A(n77), .Y(n948) );
  BUFX2 U183 ( .A(n80), .Y(n950) );
  INVX1 U184 ( .A(n38), .Y(n936) );
  INVX1 U217 ( .A(n40), .Y(n938) );
  INVX1 U218 ( .A(n41), .Y(n939) );
  INVX1 U251 ( .A(n43), .Y(n940) );
  INVX1 U252 ( .A(n44), .Y(n941) );
  INVX1 U285 ( .A(n45), .Y(n942) );
  INVX1 U286 ( .A(n47), .Y(n943) );
  INVX1 U319 ( .A(n48), .Y(n944) );
  INVX1 U320 ( .A(N24), .Y(n988) );
  AND2X2 U353 ( .A(n5), .B(n3), .Y(n1) );
  AND2X1 U354 ( .A(n787), .B(n918), .Y(n2) );
  INVX1 U387 ( .A(n2), .Y(n3) );
  AND2X1 U388 ( .A(n786), .B(n653), .Y(n4) );
  INVX1 U421 ( .A(n4), .Y(n5) );
  AND2X1 U422 ( .A(n38), .B(n68), .Y(n6) );
  INVX1 U455 ( .A(n6), .Y(n7) );
  AND2X1 U456 ( .A(n40), .B(n68), .Y(n8) );
  INVX1 U457 ( .A(n8), .Y(n9) );
  AND2X1 U490 ( .A(n41), .B(n68), .Y(n10) );
  INVX1 U491 ( .A(n10), .Y(n11) );
  AND2X1 U524 ( .A(n43), .B(n68), .Y(n12) );
  INVX1 U525 ( .A(n12), .Y(n13) );
  AND2X1 U558 ( .A(n44), .B(n68), .Y(n14) );
  INVX1 U559 ( .A(n14), .Y(n15) );
  AND2X1 U560 ( .A(n45), .B(n68), .Y(n16) );
  INVX1 U563 ( .A(n16), .Y(n17) );
  AND2X1 U564 ( .A(n47), .B(n68), .Y(n18) );
  INVX1 U567 ( .A(n18), .Y(n19) );
  AND2X1 U568 ( .A(n48), .B(n68), .Y(n20) );
  INVX1 U571 ( .A(n20), .Y(n21) );
  AND2X1 U572 ( .A(n72), .B(n68), .Y(n22) );
  INVX1 U575 ( .A(n22), .Y(n23) );
  AND2X1 U576 ( .A(n75), .B(n68), .Y(n24) );
  INVX1 U579 ( .A(n24), .Y(n25) );
  AND2X1 U580 ( .A(n78), .B(n68), .Y(n26) );
  INVX1 U583 ( .A(n26), .Y(n27) );
  AND2X1 U584 ( .A(n81), .B(n68), .Y(n28) );
  INVX1 U587 ( .A(n28), .Y(n29) );
  AND2X1 U588 ( .A(n50), .B(n68), .Y(n30) );
  INVX1 U591 ( .A(n30), .Y(n31) );
  AND2X1 U592 ( .A(n51), .B(n68), .Y(n32) );
  INVX1 U595 ( .A(n32), .Y(n33) );
  AND2X1 U596 ( .A(n84), .B(n68), .Y(n34) );
  INVX1 U599 ( .A(n34), .Y(n35) );
  AND2X1 U600 ( .A(n87), .B(n68), .Y(n36) );
  INVX1 U603 ( .A(n36), .Y(n37) );
  AND2X1 U604 ( .A(n646), .B(n638), .Y(n38) );
  AND2X1 U607 ( .A(n648), .B(n640), .Y(n39) );
  AND2X1 U608 ( .A(n646), .B(n642), .Y(n40) );
  AND2X1 U609 ( .A(n646), .B(n1262), .Y(n41) );
  AND2X1 U612 ( .A(n646), .B(n1264), .Y(n43) );
  AND2X1 U613 ( .A(n650), .B(n638), .Y(n44) );
  AND2X1 U616 ( .A(n650), .B(n642), .Y(n45) );
  AND2X1 U617 ( .A(n650), .B(n1262), .Y(n47) );
  AND2X1 U620 ( .A(n650), .B(n1264), .Y(n48) );
  AND2X1 U621 ( .A(n638), .B(n1265), .Y(n50) );
  AND2X1 U622 ( .A(n642), .B(n1265), .Y(n51) );
  AND2X1 U625 ( .A(n648), .B(n644), .Y(n53) );
  AND2X1 U626 ( .A(n648), .B(n1476), .Y(n54) );
  AND2X1 U627 ( .A(n648), .B(n1493), .Y(n56) );
  AND2X1 U628 ( .A(n652), .B(n640), .Y(n57) );
  AND2X1 U629 ( .A(n652), .B(n644), .Y(n59) );
  AND2X1 U630 ( .A(n652), .B(n1476), .Y(n60) );
  AND2X1 U631 ( .A(n652), .B(n1493), .Y(n62) );
  AND2X1 U632 ( .A(n640), .B(n1494), .Y(n63) );
  AND2X1 U633 ( .A(n644), .B(n1494), .Y(n65) );
  OR2X1 U634 ( .A(n990), .B(rst), .Y(n66) );
  AND2X1 U635 ( .A(n39), .B(n1495), .Y(n69) );
  INVX1 U636 ( .A(n69), .Y(n71) );
  AND2X1 U637 ( .A(n1258), .B(n638), .Y(n72) );
  INVX1 U638 ( .A(n72), .Y(n74) );
  AND2X1 U639 ( .A(n1258), .B(n642), .Y(n75) );
  INVX1 U640 ( .A(n75), .Y(n77) );
  AND2X1 U641 ( .A(n1258), .B(n1262), .Y(n78) );
  INVX1 U642 ( .A(n78), .Y(n80) );
  AND2X1 U643 ( .A(n1258), .B(n1264), .Y(n81) );
  INVX1 U644 ( .A(n81), .Y(n83) );
  AND2X1 U645 ( .A(n1262), .B(n1265), .Y(n84) );
  INVX1 U646 ( .A(n84), .Y(n86) );
  AND2X1 U647 ( .A(n1265), .B(n1264), .Y(n87) );
  INVX1 U648 ( .A(n87), .Y(n89) );
  AND2X1 U649 ( .A(n53), .B(n1495), .Y(n93) );
  INVX1 U650 ( .A(n93), .Y(n95) );
  AND2X1 U651 ( .A(n54), .B(n1495), .Y(n112) );
  INVX1 U652 ( .A(n112), .Y(n114) );
  AND2X1 U653 ( .A(n56), .B(n1495), .Y(n130) );
  INVX1 U654 ( .A(n130), .Y(n131) );
  AND2X1 U655 ( .A(n57), .B(n1495), .Y(n133) );
  INVX1 U656 ( .A(n133), .Y(n149) );
  AND2X1 U657 ( .A(n59), .B(n1495), .Y(n150) );
  INVX1 U658 ( .A(n150), .Y(n152) );
  AND2X1 U659 ( .A(n60), .B(n1495), .Y(n169) );
  INVX1 U660 ( .A(n169), .Y(n171) );
  AND2X1 U661 ( .A(n62), .B(n1495), .Y(n187) );
  AND2X1 U662 ( .A(n1427), .B(n640), .Y(n205) );
  INVX1 U663 ( .A(n205), .Y(n207) );
  AND2X1 U664 ( .A(n205), .B(n1495), .Y(n223) );
  INVX1 U665 ( .A(n223), .Y(n225) );
  AND2X1 U666 ( .A(n1427), .B(n644), .Y(n241) );
  INVX1 U667 ( .A(n241), .Y(n242) );
  AND2X1 U668 ( .A(n241), .B(n1495), .Y(n244) );
  INVX1 U669 ( .A(n244), .Y(n260) );
  AND2X1 U670 ( .A(n1427), .B(n1476), .Y(n262) );
  INVX1 U671 ( .A(n262), .Y(n278) );
  AND2X1 U672 ( .A(n262), .B(n1495), .Y(n280) );
  INVX1 U673 ( .A(n280), .Y(n296) );
  AND2X1 U674 ( .A(n1427), .B(n1493), .Y(n298) );
  INVX1 U675 ( .A(n298), .Y(n314) );
  AND2X1 U676 ( .A(n298), .B(n1495), .Y(n315) );
  INVX1 U677 ( .A(n315), .Y(n317) );
  AND2X1 U678 ( .A(n63), .B(n1495), .Y(n333) );
  INVX1 U679 ( .A(n333), .Y(n335) );
  AND2X1 U680 ( .A(n65), .B(n1495), .Y(n351) );
  INVX1 U681 ( .A(n351), .Y(n353) );
  AND2X1 U682 ( .A(n1476), .B(n1494), .Y(n354) );
  INVX1 U683 ( .A(n354), .Y(n360) );
  AND2X1 U684 ( .A(n354), .B(n1495), .Y(n362) );
  INVX1 U685 ( .A(n362), .Y(n369) );
  AND2X1 U686 ( .A(n1494), .B(n1493), .Y(n374) );
  INVX1 U687 ( .A(n374), .Y(n634) );
  AND2X1 U688 ( .A(n1495), .B(n374), .Y(n635) );
  INVX1 U689 ( .A(n635), .Y(n636) );
  OR2X1 U690 ( .A(n980), .B(n982), .Y(n637) );
  INVX1 U691 ( .A(n637), .Y(n638) );
  OR2X1 U692 ( .A(n986), .B(N23), .Y(n639) );
  INVX1 U693 ( .A(n639), .Y(n640) );
  OR2X1 U694 ( .A(n981), .B(n982), .Y(n641) );
  INVX1 U695 ( .A(n641), .Y(n642) );
  OR2X1 U696 ( .A(n987), .B(N23), .Y(n643) );
  INVX1 U697 ( .A(n643), .Y(n644) );
  OR2X1 U698 ( .A(n984), .B(N21), .Y(n645) );
  INVX1 U699 ( .A(n645), .Y(n646) );
  OR2X1 U700 ( .A(N24), .B(N25), .Y(n647) );
  INVX1 U701 ( .A(n647), .Y(n648) );
  OR2X1 U702 ( .A(n985), .B(N21), .Y(n649) );
  INVX1 U703 ( .A(n649), .Y(n650) );
  OR2X1 U704 ( .A(n988), .B(N25), .Y(n651) );
  INVX1 U705 ( .A(n651), .Y(n652) );
  INVX1 U706 ( .A(n918), .Y(n653) );
  MUX2X1 U707 ( .B(\mem<65> ), .A(\mem<64> ), .S(n922), .Y(n834) );
  MUX2X1 U708 ( .B(\mem<81> ), .A(\mem<80> ), .S(n922), .Y(n819) );
  MUX2X1 U709 ( .B(\mem<69> ), .A(\mem<68> ), .S(n922), .Y(n831) );
  MUX2X1 U710 ( .B(\mem<85> ), .A(\mem<84> ), .S(n922), .Y(n816) );
  INVX1 U711 ( .A(N19), .Y(n983) );
  MUX2X1 U712 ( .B(n655), .A(n656), .S(n920), .Y(n654) );
  MUX2X1 U713 ( .B(n658), .A(n659), .S(n920), .Y(n657) );
  MUX2X1 U714 ( .B(n661), .A(n662), .S(n920), .Y(n660) );
  MUX2X1 U715 ( .B(n664), .A(n665), .S(n920), .Y(n663) );
  MUX2X1 U716 ( .B(n667), .A(n668), .S(n909), .Y(n666) );
  MUX2X1 U717 ( .B(n670), .A(n671), .S(n920), .Y(n669) );
  MUX2X1 U718 ( .B(n673), .A(n674), .S(n920), .Y(n672) );
  MUX2X1 U719 ( .B(n676), .A(n677), .S(n920), .Y(n675) );
  MUX2X1 U720 ( .B(n679), .A(n680), .S(n920), .Y(n678) );
  MUX2X1 U721 ( .B(n682), .A(n683), .S(n909), .Y(n681) );
  MUX2X1 U722 ( .B(n685), .A(n686), .S(n920), .Y(n684) );
  MUX2X1 U723 ( .B(n688), .A(n689), .S(n920), .Y(n687) );
  MUX2X1 U724 ( .B(n691), .A(n692), .S(n920), .Y(n690) );
  MUX2X1 U725 ( .B(n694), .A(n695), .S(n920), .Y(n693) );
  MUX2X1 U726 ( .B(n697), .A(n698), .S(n909), .Y(n696) );
  MUX2X1 U727 ( .B(n700), .A(n701), .S(n919), .Y(n699) );
  MUX2X1 U728 ( .B(n703), .A(n704), .S(n919), .Y(n702) );
  MUX2X1 U729 ( .B(n706), .A(n707), .S(n919), .Y(n705) );
  MUX2X1 U730 ( .B(n709), .A(n710), .S(n919), .Y(n708) );
  MUX2X1 U731 ( .B(n712), .A(n713), .S(n909), .Y(n711) );
  MUX2X1 U732 ( .B(n715), .A(n716), .S(N23), .Y(n714) );
  MUX2X1 U733 ( .B(n718), .A(n719), .S(n919), .Y(n717) );
  MUX2X1 U734 ( .B(n721), .A(n722), .S(n919), .Y(n720) );
  MUX2X1 U735 ( .B(n724), .A(n725), .S(n919), .Y(n723) );
  MUX2X1 U736 ( .B(n727), .A(n728), .S(n919), .Y(n726) );
  MUX2X1 U737 ( .B(n730), .A(n731), .S(n909), .Y(n729) );
  MUX2X1 U738 ( .B(n733), .A(n734), .S(n919), .Y(n732) );
  MUX2X1 U739 ( .B(n736), .A(n737), .S(n919), .Y(n735) );
  MUX2X1 U740 ( .B(n739), .A(n740), .S(n919), .Y(n738) );
  MUX2X1 U741 ( .B(n742), .A(n743), .S(n919), .Y(n741) );
  MUX2X1 U742 ( .B(n745), .A(n746), .S(n909), .Y(n744) );
  MUX2X1 U743 ( .B(n748), .A(n749), .S(n918), .Y(n747) );
  MUX2X1 U744 ( .B(n751), .A(n752), .S(n918), .Y(n750) );
  MUX2X1 U745 ( .B(n754), .A(n755), .S(n918), .Y(n753) );
  MUX2X1 U746 ( .B(n757), .A(n758), .S(n918), .Y(n756) );
  MUX2X1 U747 ( .B(n760), .A(n761), .S(n909), .Y(n759) );
  MUX2X1 U748 ( .B(n763), .A(n764), .S(n918), .Y(n762) );
  MUX2X1 U749 ( .B(n766), .A(n767), .S(n918), .Y(n765) );
  MUX2X1 U750 ( .B(n769), .A(n770), .S(n918), .Y(n768) );
  MUX2X1 U751 ( .B(n772), .A(n773), .S(n918), .Y(n771) );
  MUX2X1 U752 ( .B(n775), .A(n776), .S(n909), .Y(n774) );
  MUX2X1 U753 ( .B(n778), .A(n779), .S(N23), .Y(n777) );
  MUX2X1 U754 ( .B(n781), .A(n782), .S(n918), .Y(n780) );
  MUX2X1 U755 ( .B(n784), .A(n785), .S(n918), .Y(n783) );
  MUX2X1 U756 ( .B(n789), .A(n790), .S(n918), .Y(n788) );
  MUX2X1 U757 ( .B(n792), .A(n793), .S(n909), .Y(n791) );
  MUX2X1 U758 ( .B(n795), .A(n796), .S(n917), .Y(n794) );
  MUX2X1 U759 ( .B(n798), .A(n799), .S(n917), .Y(n797) );
  MUX2X1 U760 ( .B(n801), .A(n802), .S(n917), .Y(n800) );
  MUX2X1 U761 ( .B(n804), .A(n805), .S(n917), .Y(n803) );
  MUX2X1 U762 ( .B(n807), .A(n808), .S(n909), .Y(n806) );
  MUX2X1 U763 ( .B(n810), .A(n811), .S(n917), .Y(n809) );
  MUX2X1 U764 ( .B(n813), .A(n814), .S(n917), .Y(n812) );
  MUX2X1 U765 ( .B(n816), .A(n817), .S(n917), .Y(n815) );
  MUX2X1 U766 ( .B(n819), .A(n820), .S(n917), .Y(n818) );
  MUX2X1 U767 ( .B(n822), .A(n823), .S(n909), .Y(n821) );
  MUX2X1 U768 ( .B(n825), .A(n826), .S(n917), .Y(n824) );
  MUX2X1 U769 ( .B(n828), .A(n829), .S(n917), .Y(n827) );
  MUX2X1 U770 ( .B(n831), .A(n832), .S(n917), .Y(n830) );
  MUX2X1 U771 ( .B(n834), .A(n835), .S(n917), .Y(n833) );
  MUX2X1 U772 ( .B(n837), .A(n838), .S(n909), .Y(n836) );
  MUX2X1 U773 ( .B(n840), .A(n841), .S(N23), .Y(n839) );
  MUX2X1 U774 ( .B(n843), .A(n844), .S(n916), .Y(n842) );
  MUX2X1 U775 ( .B(n846), .A(n847), .S(n916), .Y(n845) );
  MUX2X1 U776 ( .B(n849), .A(n850), .S(n916), .Y(n848) );
  MUX2X1 U777 ( .B(n852), .A(n853), .S(n916), .Y(n851) );
  MUX2X1 U778 ( .B(n855), .A(n856), .S(n908), .Y(n854) );
  MUX2X1 U779 ( .B(n858), .A(n859), .S(n916), .Y(n857) );
  MUX2X1 U780 ( .B(n861), .A(n862), .S(n916), .Y(n860) );
  MUX2X1 U781 ( .B(n864), .A(n865), .S(n916), .Y(n863) );
  MUX2X1 U782 ( .B(n867), .A(n868), .S(n916), .Y(n866) );
  MUX2X1 U783 ( .B(n870), .A(n871), .S(n908), .Y(n869) );
  MUX2X1 U784 ( .B(n873), .A(n874), .S(n916), .Y(n872) );
  MUX2X1 U785 ( .B(n876), .A(n877), .S(n916), .Y(n875) );
  MUX2X1 U786 ( .B(n879), .A(n880), .S(n916), .Y(n878) );
  MUX2X1 U787 ( .B(n882), .A(n883), .S(n916), .Y(n881) );
  MUX2X1 U788 ( .B(n885), .A(n886), .S(n908), .Y(n884) );
  MUX2X1 U789 ( .B(n888), .A(n889), .S(n915), .Y(n887) );
  MUX2X1 U790 ( .B(n891), .A(n892), .S(n915), .Y(n890) );
  MUX2X1 U791 ( .B(n894), .A(n895), .S(n915), .Y(n893) );
  MUX2X1 U792 ( .B(n897), .A(n898), .S(n915), .Y(n896) );
  MUX2X1 U793 ( .B(n900), .A(n901), .S(n908), .Y(n899) );
  MUX2X1 U794 ( .B(n903), .A(n904), .S(N23), .Y(n902) );
  MUX2X1 U795 ( .B(n905), .A(n906), .S(N25), .Y(N28) );
  MUX2X1 U796 ( .B(\mem<254> ), .A(\mem<255> ), .S(n929), .Y(n656) );
  MUX2X1 U797 ( .B(\mem<252> ), .A(\mem<253> ), .S(n927), .Y(n655) );
  MUX2X1 U798 ( .B(\mem<250> ), .A(\mem<251> ), .S(n927), .Y(n659) );
  MUX2X1 U799 ( .B(\mem<248> ), .A(\mem<249> ), .S(n929), .Y(n658) );
  MUX2X1 U800 ( .B(n657), .A(n654), .S(n912), .Y(n668) );
  MUX2X1 U801 ( .B(\mem<246> ), .A(\mem<247> ), .S(n927), .Y(n662) );
  MUX2X1 U802 ( .B(\mem<244> ), .A(\mem<245> ), .S(n927), .Y(n661) );
  MUX2X1 U803 ( .B(\mem<242> ), .A(\mem<243> ), .S(n927), .Y(n665) );
  MUX2X1 U804 ( .B(\mem<240> ), .A(\mem<241> ), .S(n927), .Y(n664) );
  MUX2X1 U805 ( .B(n663), .A(n660), .S(n912), .Y(n667) );
  MUX2X1 U806 ( .B(\mem<238> ), .A(\mem<239> ), .S(n925), .Y(n671) );
  MUX2X1 U807 ( .B(\mem<236> ), .A(\mem<237> ), .S(n925), .Y(n670) );
  MUX2X1 U808 ( .B(\mem<234> ), .A(\mem<235> ), .S(n925), .Y(n674) );
  MUX2X1 U809 ( .B(\mem<232> ), .A(\mem<233> ), .S(n925), .Y(n673) );
  MUX2X1 U810 ( .B(n672), .A(n669), .S(n912), .Y(n683) );
  MUX2X1 U811 ( .B(\mem<230> ), .A(\mem<231> ), .S(n925), .Y(n677) );
  MUX2X1 U812 ( .B(\mem<228> ), .A(\mem<229> ), .S(n925), .Y(n676) );
  MUX2X1 U813 ( .B(\mem<226> ), .A(\mem<227> ), .S(n925), .Y(n680) );
  MUX2X1 U814 ( .B(\mem<224> ), .A(\mem<225> ), .S(n925), .Y(n679) );
  MUX2X1 U815 ( .B(n678), .A(n675), .S(n912), .Y(n682) );
  MUX2X1 U816 ( .B(n681), .A(n666), .S(n986), .Y(n716) );
  MUX2X1 U817 ( .B(\mem<222> ), .A(\mem<223> ), .S(n925), .Y(n686) );
  MUX2X1 U818 ( .B(\mem<220> ), .A(\mem<221> ), .S(n925), .Y(n685) );
  MUX2X1 U819 ( .B(\mem<218> ), .A(\mem<219> ), .S(n925), .Y(n689) );
  MUX2X1 U820 ( .B(\mem<216> ), .A(\mem<217> ), .S(n925), .Y(n688) );
  MUX2X1 U821 ( .B(n687), .A(n684), .S(n912), .Y(n698) );
  MUX2X1 U822 ( .B(\mem<214> ), .A(\mem<215> ), .S(n926), .Y(n692) );
  MUX2X1 U823 ( .B(\mem<212> ), .A(\mem<213> ), .S(n926), .Y(n691) );
  MUX2X1 U824 ( .B(\mem<210> ), .A(\mem<211> ), .S(n926), .Y(n695) );
  MUX2X1 U825 ( .B(\mem<208> ), .A(\mem<209> ), .S(n926), .Y(n694) );
  MUX2X1 U826 ( .B(n693), .A(n690), .S(n912), .Y(n697) );
  MUX2X1 U827 ( .B(\mem<206> ), .A(\mem<207> ), .S(n926), .Y(n701) );
  MUX2X1 U828 ( .B(\mem<204> ), .A(\mem<205> ), .S(n926), .Y(n700) );
  MUX2X1 U829 ( .B(\mem<202> ), .A(\mem<203> ), .S(n926), .Y(n704) );
  MUX2X1 U830 ( .B(\mem<200> ), .A(\mem<201> ), .S(n926), .Y(n703) );
  MUX2X1 U831 ( .B(n702), .A(n699), .S(n912), .Y(n713) );
  MUX2X1 U832 ( .B(\mem<198> ), .A(\mem<199> ), .S(n926), .Y(n707) );
  MUX2X1 U833 ( .B(\mem<196> ), .A(\mem<197> ), .S(n926), .Y(n706) );
  MUX2X1 U834 ( .B(\mem<194> ), .A(\mem<195> ), .S(n926), .Y(n710) );
  MUX2X1 U835 ( .B(\mem<192> ), .A(\mem<193> ), .S(n926), .Y(n709) );
  MUX2X1 U836 ( .B(n708), .A(n705), .S(n912), .Y(n712) );
  MUX2X1 U837 ( .B(n711), .A(n696), .S(n986), .Y(n715) );
  MUX2X1 U838 ( .B(\mem<190> ), .A(\mem<191> ), .S(n927), .Y(n719) );
  MUX2X1 U839 ( .B(\mem<188> ), .A(\mem<189> ), .S(n927), .Y(n718) );
  MUX2X1 U840 ( .B(\mem<186> ), .A(\mem<187> ), .S(n927), .Y(n722) );
  MUX2X1 U841 ( .B(\mem<184> ), .A(\mem<185> ), .S(n927), .Y(n721) );
  MUX2X1 U842 ( .B(n720), .A(n717), .S(n912), .Y(n731) );
  MUX2X1 U843 ( .B(\mem<182> ), .A(\mem<183> ), .S(n927), .Y(n725) );
  MUX2X1 U844 ( .B(\mem<180> ), .A(\mem<181> ), .S(n927), .Y(n724) );
  MUX2X1 U845 ( .B(\mem<178> ), .A(\mem<179> ), .S(n927), .Y(n728) );
  MUX2X1 U846 ( .B(\mem<176> ), .A(\mem<177> ), .S(n927), .Y(n727) );
  MUX2X1 U847 ( .B(n726), .A(n723), .S(n912), .Y(n730) );
  MUX2X1 U848 ( .B(\mem<174> ), .A(\mem<175> ), .S(n927), .Y(n734) );
  MUX2X1 U849 ( .B(\mem<172> ), .A(\mem<173> ), .S(n927), .Y(n733) );
  MUX2X1 U850 ( .B(\mem<170> ), .A(\mem<171> ), .S(n927), .Y(n737) );
  MUX2X1 U851 ( .B(\mem<168> ), .A(\mem<169> ), .S(n927), .Y(n736) );
  MUX2X1 U852 ( .B(n735), .A(n732), .S(n912), .Y(n746) );
  MUX2X1 U853 ( .B(\mem<166> ), .A(\mem<167> ), .S(n928), .Y(n740) );
  MUX2X1 U854 ( .B(\mem<164> ), .A(\mem<165> ), .S(n928), .Y(n739) );
  MUX2X1 U855 ( .B(\mem<162> ), .A(\mem<163> ), .S(n928), .Y(n743) );
  MUX2X1 U856 ( .B(\mem<160> ), .A(\mem<161> ), .S(n928), .Y(n742) );
  MUX2X1 U857 ( .B(n741), .A(n738), .S(n912), .Y(n745) );
  MUX2X1 U858 ( .B(n744), .A(n729), .S(n986), .Y(n779) );
  MUX2X1 U859 ( .B(\mem<158> ), .A(\mem<159> ), .S(n928), .Y(n749) );
  MUX2X1 U860 ( .B(\mem<156> ), .A(\mem<157> ), .S(n928), .Y(n748) );
  MUX2X1 U861 ( .B(\mem<154> ), .A(\mem<155> ), .S(n928), .Y(n752) );
  MUX2X1 U862 ( .B(\mem<152> ), .A(\mem<153> ), .S(n928), .Y(n751) );
  MUX2X1 U863 ( .B(n750), .A(n747), .S(n911), .Y(n761) );
  MUX2X1 U864 ( .B(\mem<150> ), .A(\mem<151> ), .S(n928), .Y(n755) );
  MUX2X1 U865 ( .B(\mem<148> ), .A(\mem<149> ), .S(n928), .Y(n754) );
  MUX2X1 U866 ( .B(\mem<146> ), .A(\mem<147> ), .S(n928), .Y(n758) );
  MUX2X1 U867 ( .B(\mem<144> ), .A(\mem<145> ), .S(n928), .Y(n757) );
  MUX2X1 U868 ( .B(n756), .A(n753), .S(n911), .Y(n760) );
  MUX2X1 U869 ( .B(\mem<142> ), .A(\mem<143> ), .S(n929), .Y(n764) );
  MUX2X1 U870 ( .B(\mem<140> ), .A(\mem<141> ), .S(n929), .Y(n763) );
  MUX2X1 U871 ( .B(\mem<138> ), .A(\mem<139> ), .S(n929), .Y(n767) );
  MUX2X1 U872 ( .B(\mem<136> ), .A(\mem<137> ), .S(n929), .Y(n766) );
  MUX2X1 U873 ( .B(n765), .A(n762), .S(n911), .Y(n776) );
  MUX2X1 U874 ( .B(\mem<134> ), .A(\mem<135> ), .S(n929), .Y(n770) );
  MUX2X1 U875 ( .B(\mem<132> ), .A(\mem<133> ), .S(n929), .Y(n769) );
  MUX2X1 U876 ( .B(\mem<130> ), .A(\mem<131> ), .S(n929), .Y(n773) );
  MUX2X1 U877 ( .B(\mem<128> ), .A(\mem<129> ), .S(n929), .Y(n772) );
  MUX2X1 U878 ( .B(n771), .A(n768), .S(n911), .Y(n775) );
  MUX2X1 U879 ( .B(n774), .A(n759), .S(n986), .Y(n778) );
  MUX2X1 U880 ( .B(n777), .A(n714), .S(N24), .Y(n906) );
  MUX2X1 U881 ( .B(\mem<126> ), .A(\mem<127> ), .S(n929), .Y(n782) );
  MUX2X1 U882 ( .B(\mem<124> ), .A(\mem<125> ), .S(n929), .Y(n781) );
  MUX2X1 U883 ( .B(\mem<122> ), .A(\mem<123> ), .S(n929), .Y(n785) );
  MUX2X1 U884 ( .B(\mem<120> ), .A(\mem<121> ), .S(n929), .Y(n784) );
  MUX2X1 U885 ( .B(n783), .A(n780), .S(n911), .Y(n793) );
  MUX2X1 U886 ( .B(\mem<118> ), .A(\mem<119> ), .S(n930), .Y(n787) );
  MUX2X1 U887 ( .B(\mem<116> ), .A(\mem<117> ), .S(n930), .Y(n786) );
  MUX2X1 U888 ( .B(\mem<114> ), .A(\mem<115> ), .S(n930), .Y(n790) );
  MUX2X1 U889 ( .B(\mem<112> ), .A(\mem<113> ), .S(n930), .Y(n789) );
  MUX2X1 U890 ( .B(n788), .A(n1), .S(n911), .Y(n792) );
  MUX2X1 U891 ( .B(\mem<110> ), .A(\mem<111> ), .S(n930), .Y(n796) );
  MUX2X1 U892 ( .B(\mem<108> ), .A(\mem<109> ), .S(n930), .Y(n795) );
  MUX2X1 U893 ( .B(\mem<106> ), .A(\mem<107> ), .S(n930), .Y(n799) );
  MUX2X1 U894 ( .B(\mem<104> ), .A(\mem<105> ), .S(n930), .Y(n798) );
  MUX2X1 U895 ( .B(n797), .A(n794), .S(n911), .Y(n808) );
  MUX2X1 U896 ( .B(\mem<102> ), .A(\mem<103> ), .S(n930), .Y(n802) );
  MUX2X1 U897 ( .B(\mem<100> ), .A(\mem<101> ), .S(n930), .Y(n801) );
  MUX2X1 U898 ( .B(\mem<98> ), .A(\mem<99> ), .S(n930), .Y(n805) );
  MUX2X1 U899 ( .B(\mem<96> ), .A(\mem<97> ), .S(n930), .Y(n804) );
  MUX2X1 U900 ( .B(n803), .A(n800), .S(n911), .Y(n807) );
  MUX2X1 U901 ( .B(n806), .A(n791), .S(n986), .Y(n841) );
  MUX2X1 U902 ( .B(\mem<94> ), .A(\mem<95> ), .S(n931), .Y(n811) );
  MUX2X1 U903 ( .B(\mem<92> ), .A(\mem<93> ), .S(n931), .Y(n810) );
  MUX2X1 U904 ( .B(\mem<90> ), .A(\mem<91> ), .S(n931), .Y(n814) );
  MUX2X1 U905 ( .B(\mem<88> ), .A(\mem<89> ), .S(n931), .Y(n813) );
  MUX2X1 U906 ( .B(n812), .A(n809), .S(n911), .Y(n823) );
  MUX2X1 U907 ( .B(\mem<86> ), .A(\mem<87> ), .S(n931), .Y(n817) );
  MUX2X1 U908 ( .B(\mem<82> ), .A(\mem<83> ), .S(n931), .Y(n820) );
  MUX2X1 U909 ( .B(n818), .A(n815), .S(n911), .Y(n822) );
  MUX2X1 U910 ( .B(\mem<78> ), .A(\mem<79> ), .S(n931), .Y(n826) );
  MUX2X1 U911 ( .B(\mem<76> ), .A(\mem<77> ), .S(n931), .Y(n825) );
  MUX2X1 U912 ( .B(\mem<74> ), .A(\mem<75> ), .S(n931), .Y(n829) );
  MUX2X1 U913 ( .B(\mem<72> ), .A(\mem<73> ), .S(n931), .Y(n828) );
  MUX2X1 U914 ( .B(n827), .A(n824), .S(n911), .Y(n838) );
  MUX2X1 U915 ( .B(\mem<70> ), .A(\mem<71> ), .S(n932), .Y(n832) );
  MUX2X1 U916 ( .B(\mem<66> ), .A(\mem<67> ), .S(n932), .Y(n835) );
  MUX2X1 U917 ( .B(n833), .A(n830), .S(n911), .Y(n837) );
  MUX2X1 U918 ( .B(n836), .A(n821), .S(n986), .Y(n840) );
  MUX2X1 U919 ( .B(\mem<62> ), .A(\mem<63> ), .S(n932), .Y(n844) );
  MUX2X1 U920 ( .B(\mem<60> ), .A(\mem<61> ), .S(n932), .Y(n843) );
  MUX2X1 U921 ( .B(\mem<58> ), .A(\mem<59> ), .S(n932), .Y(n847) );
  MUX2X1 U922 ( .B(\mem<56> ), .A(\mem<57> ), .S(n932), .Y(n846) );
  MUX2X1 U923 ( .B(n845), .A(n842), .S(n910), .Y(n856) );
  MUX2X1 U924 ( .B(\mem<54> ), .A(\mem<55> ), .S(n932), .Y(n850) );
  MUX2X1 U925 ( .B(\mem<52> ), .A(\mem<53> ), .S(n932), .Y(n849) );
  MUX2X1 U926 ( .B(\mem<50> ), .A(\mem<51> ), .S(n932), .Y(n853) );
  MUX2X1 U927 ( .B(\mem<48> ), .A(\mem<49> ), .S(n932), .Y(n852) );
  MUX2X1 U928 ( .B(n851), .A(n848), .S(n910), .Y(n855) );
  MUX2X1 U929 ( .B(\mem<46> ), .A(\mem<47> ), .S(n933), .Y(n859) );
  MUX2X1 U930 ( .B(\mem<44> ), .A(\mem<45> ), .S(n933), .Y(n858) );
  MUX2X1 U931 ( .B(\mem<42> ), .A(\mem<43> ), .S(n933), .Y(n862) );
  MUX2X1 U932 ( .B(\mem<40> ), .A(\mem<41> ), .S(n933), .Y(n861) );
  MUX2X1 U933 ( .B(n860), .A(n857), .S(n910), .Y(n871) );
  MUX2X1 U934 ( .B(\mem<38> ), .A(\mem<39> ), .S(n933), .Y(n865) );
  MUX2X1 U935 ( .B(\mem<36> ), .A(\mem<37> ), .S(n933), .Y(n864) );
  MUX2X1 U936 ( .B(\mem<34> ), .A(\mem<35> ), .S(n933), .Y(n868) );
  MUX2X1 U937 ( .B(\mem<32> ), .A(\mem<33> ), .S(n933), .Y(n867) );
  MUX2X1 U938 ( .B(n866), .A(n863), .S(n910), .Y(n870) );
  MUX2X1 U939 ( .B(n869), .A(n854), .S(n986), .Y(n904) );
  MUX2X1 U940 ( .B(\mem<30> ), .A(\mem<31> ), .S(n933), .Y(n874) );
  MUX2X1 U941 ( .B(\mem<28> ), .A(\mem<29> ), .S(n933), .Y(n873) );
  MUX2X1 U942 ( .B(\mem<26> ), .A(\mem<27> ), .S(n933), .Y(n877) );
  MUX2X1 U943 ( .B(\mem<24> ), .A(\mem<25> ), .S(n933), .Y(n876) );
  MUX2X1 U944 ( .B(n875), .A(n872), .S(n910), .Y(n886) );
  MUX2X1 U945 ( .B(\mem<22> ), .A(\mem<23> ), .S(n929), .Y(n880) );
  MUX2X1 U946 ( .B(\mem<20> ), .A(\mem<21> ), .S(n928), .Y(n879) );
  MUX2X1 U947 ( .B(\mem<18> ), .A(\mem<19> ), .S(n927), .Y(n883) );
  MUX2X1 U948 ( .B(\mem<16> ), .A(\mem<17> ), .S(n931), .Y(n882) );
  MUX2X1 U949 ( .B(n881), .A(n878), .S(n910), .Y(n885) );
  MUX2X1 U950 ( .B(\mem<14> ), .A(\mem<15> ), .S(n927), .Y(n889) );
  MUX2X1 U951 ( .B(\mem<12> ), .A(\mem<13> ), .S(n927), .Y(n888) );
  MUX2X1 U952 ( .B(\mem<10> ), .A(\mem<11> ), .S(n928), .Y(n892) );
  MUX2X1 U953 ( .B(\mem<8> ), .A(\mem<9> ), .S(n932), .Y(n891) );
  MUX2X1 U954 ( .B(n890), .A(n887), .S(n910), .Y(n901) );
  MUX2X1 U955 ( .B(\mem<6> ), .A(\mem<7> ), .S(n929), .Y(n895) );
  MUX2X1 U956 ( .B(\mem<4> ), .A(\mem<5> ), .S(n932), .Y(n894) );
  MUX2X1 U957 ( .B(\mem<2> ), .A(\mem<3> ), .S(n931), .Y(n898) );
  MUX2X1 U958 ( .B(\mem<0> ), .A(\mem<1> ), .S(n929), .Y(n897) );
  MUX2X1 U959 ( .B(n896), .A(n893), .S(n910), .Y(n900) );
  MUX2X1 U960 ( .B(n899), .A(n884), .S(n986), .Y(n903) );
  MUX2X1 U961 ( .B(n902), .A(n839), .S(N24), .Y(n905) );
  INVX8 U962 ( .A(n907), .Y(n909) );
  INVX8 U963 ( .A(n985), .Y(n910) );
  INVX8 U964 ( .A(n985), .Y(n911) );
  INVX8 U965 ( .A(n985), .Y(n912) );
  INVX8 U966 ( .A(n982), .Y(n913) );
  INVX8 U967 ( .A(n982), .Y(n914) );
  INVX8 U968 ( .A(n914), .Y(n915) );
  INVX8 U969 ( .A(n914), .Y(n916) );
  INVX8 U970 ( .A(n914), .Y(n917) );
  INVX8 U971 ( .A(n913), .Y(n918) );
  INVX8 U972 ( .A(n913), .Y(n919) );
  INVX8 U973 ( .A(n913), .Y(n920) );
  INVX8 U974 ( .A(n980), .Y(n922) );
  INVX8 U975 ( .A(n980), .Y(n923) );
  INVX8 U976 ( .A(n935), .Y(n924) );
  INVX8 U977 ( .A(n924), .Y(n925) );
  INVX8 U978 ( .A(n924), .Y(n926) );
  INVX8 U979 ( .A(n923), .Y(n927) );
  INVX8 U980 ( .A(n923), .Y(n928) );
  INVX8 U981 ( .A(n923), .Y(n929) );
  INVX8 U982 ( .A(n922), .Y(n930) );
  INVX8 U983 ( .A(n922), .Y(n931) );
  INVX8 U984 ( .A(n922), .Y(n932) );
  INVX8 U985 ( .A(n921), .Y(n933) );
  INVX8 U986 ( .A(n934), .Y(n935) );
  INVX1 U987 ( .A(N28), .Y(n989) );
  INVX4 U988 ( .A(n981), .Y(n980) );
  INVX1 U989 ( .A(write), .Y(n990) );
  INVX1 U990 ( .A(N18), .Y(n981) );
  INVX8 U991 ( .A(n983), .Y(n982) );
  INVX8 U992 ( .A(N20), .Y(n985) );
  NOR3X1 U993 ( .A(write), .B(rst), .C(n989), .Y(data_out) );
endmodule


module final_memory_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1046, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n373, n374, n375, n376, n377, n378, n380,
         n382, n383, n384, n385, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n403, n404, n405, n406, n407,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n584, n585, n586, n587,
         n588, n589, n590, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n50, n150, n189, n289, n348, n372, n379, n381, n386, n387,
         n401, n402, n409, n421, n422, n434, n435, n447, n448, n460, n461,
         n473, n474, n486, n487, n507, n508, n522, n523, n537, n538, n552,
         n553, n567, n568, n582, n583, n591, n592, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n870), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n869), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n868), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n867), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n866), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n865), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n864), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n863), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n862), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n861), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n860), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n859), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n858), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n857), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n856), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n855), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n854), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n853), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n852), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n851), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n850), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n849), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n848), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n847), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n846), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n845), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n844), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n843), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n842), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n841), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n840), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n839), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n838), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n837), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n836), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n835), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n834), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n833), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n832), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n831), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n830), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n829), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n828), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n827), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n826), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n825), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n824), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n823), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n822), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n821), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n820), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n819), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n818), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n817), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n816), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n815), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n814), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n813), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n812), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n811), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n810), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n809), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n808), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n807), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n806), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n805), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n804), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n803), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n802), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n801), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n800), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n799), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n798), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n797), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n796), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n795), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n794), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n793), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n792), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n791), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n790), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n789), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n788), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n787), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n786), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n785), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n784), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n783), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n782), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n781), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n780), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n779), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n778), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n777), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n776), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n775), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n774), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n773), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n772), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n771), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n770), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n769), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n768), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n767), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n766), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n765), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n764), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n763), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n762), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n761), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n760), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n759), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n758), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n757), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n756), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n755), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n754), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n753), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n752), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n751), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n750), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n749), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n748), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n747), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n746), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n745), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n744), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n743), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n742), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n741), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n740), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n739), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n738), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n737), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n736), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n735), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n734), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n733), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n732), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n731), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n730), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n729), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n728), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n727), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n726), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n725), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n724), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n723), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n722), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n721), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n720), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n719), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n718), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n717), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n716), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n715), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n714), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n713), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n712), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n711), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n710), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n709), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n708), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n707), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n706), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n705), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n704), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n703), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n702), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n701), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n700), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n699), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n698), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n697), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n696), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n695), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n694), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n693), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n692), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n691), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n690), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n689), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n688), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n687), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n686), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n685), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n684), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n683), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n682), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n681), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n680), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n679), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n678), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n677), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n676), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n675), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n674), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n673), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n672), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n671), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n670), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n669), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n668), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n667), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n666), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n665), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n664), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n663), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n662), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n661), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n660), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n659), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n658), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n657), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n656), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n655), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n654), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n653), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n652), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n651), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n650), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n649), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n648), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n647), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n646), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n645), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n644), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n643), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n642), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n641), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n640), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n639), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n638), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n637), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n636), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n635), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n634), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n633), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n632), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n631), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n630), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n629), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n628), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n627), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n626), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n625), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n624), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n623), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n622), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n621), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n620), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n619), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n618), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n617), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n616), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n615), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n614), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n613), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n612), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n611), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n610), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n609), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n608), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n607), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n413), .B(n414), .Y(n412) );
  AND2X2 U10 ( .A(n418), .B(n419), .Y(n417) );
  AND2X2 U11 ( .A(n426), .B(n427), .Y(n425) );
  AND2X2 U12 ( .A(n431), .B(n432), .Y(n430) );
  AND2X2 U13 ( .A(n439), .B(n440), .Y(n438) );
  AND2X2 U14 ( .A(n444), .B(n445), .Y(n443) );
  AND2X2 U15 ( .A(n452), .B(n453), .Y(n451) );
  AND2X2 U16 ( .A(n457), .B(n458), .Y(n456) );
  AND2X2 U17 ( .A(n465), .B(n466), .Y(n464) );
  AND2X2 U18 ( .A(n470), .B(n471), .Y(n469) );
  AND2X2 U19 ( .A(n478), .B(n479), .Y(n477) );
  AND2X2 U20 ( .A(n483), .B(n484), .Y(n482) );
  AND2X2 U21 ( .A(n491), .B(n492), .Y(n490) );
  AND2X2 U22 ( .A(n496), .B(n497), .Y(n495) );
  AND2X2 U30 ( .A(n588), .B(n1026), .Y(n248) );
  AND2X2 U31 ( .A(n589), .B(n1026), .Y(n91) );
  AND2X2 U32 ( .A(n588), .B(\addr_1c<0> ), .Y(n228) );
  AND2X2 U33 ( .A(n589), .B(\addr_1c<0> ), .Y(n71) );
  AND2X2 U34 ( .A(n596), .B(n597), .Y(n595) );
  AND2X2 U45 ( .A(n603), .B(n604), .Y(n602) );
  NOR3X1 U94 ( .A(n1014), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1015), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1038), .C(n40), .Y(n607) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n40) );
  OAI21X1 U98 ( .A(n1011), .B(n1039), .C(n41), .Y(n608) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n41) );
  OAI21X1 U100 ( .A(n1011), .B(n1040), .C(n42), .Y(n609) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n42) );
  OAI21X1 U102 ( .A(n1011), .B(n1041), .C(n43), .Y(n610) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n43) );
  OAI21X1 U104 ( .A(n1011), .B(n1042), .C(n44), .Y(n611) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n44) );
  OAI21X1 U106 ( .A(n1011), .B(n1043), .C(n45), .Y(n612) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n45) );
  OAI21X1 U108 ( .A(n1011), .B(n1044), .C(n46), .Y(n613) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n46) );
  OAI21X1 U110 ( .A(n1011), .B(n1045), .C(n47), .Y(n614) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n47) );
  NAND3X1 U112 ( .A(n48), .B(n49), .C(n965), .Y(n39) );
  OAI21X1 U113 ( .A(n6), .B(n1030), .C(n51), .Y(n615) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n51) );
  OAI21X1 U115 ( .A(n6), .B(n1031), .C(n52), .Y(n616) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n52) );
  OAI21X1 U117 ( .A(n6), .B(n1032), .C(n53), .Y(n617) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n53) );
  OAI21X1 U119 ( .A(n6), .B(n1033), .C(n54), .Y(n618) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n54) );
  OAI21X1 U121 ( .A(n6), .B(n1034), .C(n55), .Y(n619) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n55) );
  OAI21X1 U123 ( .A(n6), .B(n1035), .C(n56), .Y(n620) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n56) );
  OAI21X1 U125 ( .A(n6), .B(n1036), .C(n57), .Y(n621) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n57) );
  OAI21X1 U127 ( .A(n6), .B(n1037), .C(n58), .Y(n622) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n58) );
  OAI21X1 U130 ( .A(n1038), .B(n1010), .C(n62), .Y(n623) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n62) );
  OAI21X1 U132 ( .A(n1039), .B(n1009), .C(n63), .Y(n624) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n63) );
  OAI21X1 U134 ( .A(n1040), .B(n1009), .C(n64), .Y(n625) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n64) );
  OAI21X1 U136 ( .A(n1041), .B(n1009), .C(n65), .Y(n626) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n65) );
  OAI21X1 U138 ( .A(n1042), .B(n1009), .C(n66), .Y(n627) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n66) );
  OAI21X1 U140 ( .A(n1043), .B(n1009), .C(n67), .Y(n628) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n67) );
  OAI21X1 U142 ( .A(n1044), .B(n1009), .C(n68), .Y(n629) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n68) );
  OAI21X1 U144 ( .A(n1045), .B(n1009), .C(n69), .Y(n630) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n69) );
  NAND3X1 U146 ( .A(n70), .B(n48), .C(n71), .Y(n61) );
  OAI21X1 U147 ( .A(n1030), .B(n1008), .C(n73), .Y(n631) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n73) );
  OAI21X1 U149 ( .A(n1031), .B(n1008), .C(n74), .Y(n632) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n74) );
  OAI21X1 U151 ( .A(n1032), .B(n1008), .C(n75), .Y(n633) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n75) );
  OAI21X1 U153 ( .A(n1033), .B(n1008), .C(n76), .Y(n634) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n76) );
  OAI21X1 U155 ( .A(n1034), .B(n1008), .C(n77), .Y(n635) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n77) );
  OAI21X1 U157 ( .A(n1035), .B(n1008), .C(n78), .Y(n636) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n78) );
  OAI21X1 U159 ( .A(n1036), .B(n1008), .C(n79), .Y(n637) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n79) );
  OAI21X1 U161 ( .A(n1037), .B(n1008), .C(n80), .Y(n638) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n80) );
  NAND3X1 U163 ( .A(n973), .B(n48), .C(n81), .Y(n72) );
  OAI21X1 U164 ( .A(n1038), .B(n1007), .C(n83), .Y(n639) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n83) );
  OAI21X1 U166 ( .A(n1039), .B(n1006), .C(n84), .Y(n640) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n84) );
  OAI21X1 U168 ( .A(n1040), .B(n1006), .C(n85), .Y(n641) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n85) );
  OAI21X1 U170 ( .A(n1041), .B(n1006), .C(n86), .Y(n642) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n86) );
  OAI21X1 U172 ( .A(n1042), .B(n1006), .C(n87), .Y(n643) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n87) );
  OAI21X1 U174 ( .A(n1043), .B(n1006), .C(n88), .Y(n644) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n88) );
  OAI21X1 U176 ( .A(n1044), .B(n1006), .C(n89), .Y(n645) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n89) );
  OAI21X1 U178 ( .A(n1045), .B(n1006), .C(n90), .Y(n646) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n90) );
  NAND3X1 U180 ( .A(n70), .B(n48), .C(n91), .Y(n82) );
  OAI21X1 U181 ( .A(n1030), .B(n1005), .C(n93), .Y(n647) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n93) );
  OAI21X1 U183 ( .A(n1031), .B(n1005), .C(n94), .Y(n648) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n94) );
  OAI21X1 U185 ( .A(n1032), .B(n1005), .C(n95), .Y(n649) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n95) );
  OAI21X1 U187 ( .A(n1033), .B(n1005), .C(n96), .Y(n650) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n96) );
  OAI21X1 U189 ( .A(n1034), .B(n1005), .C(n97), .Y(n651) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n97) );
  OAI21X1 U191 ( .A(n1035), .B(n1005), .C(n98), .Y(n652) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n98) );
  OAI21X1 U193 ( .A(n1036), .B(n1005), .C(n99), .Y(n653) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n99) );
  OAI21X1 U195 ( .A(n1037), .B(n1005), .C(n100), .Y(n654) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n100) );
  NAND3X1 U197 ( .A(n973), .B(n48), .C(n101), .Y(n92) );
  OAI21X1 U198 ( .A(n1038), .B(n1004), .C(n103), .Y(n655) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n103) );
  OAI21X1 U200 ( .A(n1039), .B(n1003), .C(n104), .Y(n656) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n104) );
  OAI21X1 U202 ( .A(n1040), .B(n1003), .C(n105), .Y(n657) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n105) );
  OAI21X1 U204 ( .A(n1041), .B(n1003), .C(n106), .Y(n658) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n106) );
  OAI21X1 U206 ( .A(n1042), .B(n1003), .C(n107), .Y(n659) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n107) );
  OAI21X1 U208 ( .A(n1043), .B(n1003), .C(n108), .Y(n660) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n108) );
  OAI21X1 U210 ( .A(n1044), .B(n1003), .C(n109), .Y(n661) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n109) );
  OAI21X1 U212 ( .A(n1045), .B(n1003), .C(n110), .Y(n662) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n110) );
  NAND3X1 U214 ( .A(n71), .B(n48), .C(n111), .Y(n102) );
  OAI21X1 U215 ( .A(n1030), .B(n1002), .C(n113), .Y(n663) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n113) );
  OAI21X1 U217 ( .A(n1031), .B(n1002), .C(n114), .Y(n664) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n114) );
  OAI21X1 U219 ( .A(n1032), .B(n1002), .C(n115), .Y(n665) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n115) );
  OAI21X1 U221 ( .A(n1033), .B(n1002), .C(n116), .Y(n666) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n116) );
  OAI21X1 U223 ( .A(n1034), .B(n1002), .C(n117), .Y(n667) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n117) );
  OAI21X1 U225 ( .A(n1035), .B(n1002), .C(n118), .Y(n668) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n118) );
  OAI21X1 U227 ( .A(n1036), .B(n1002), .C(n119), .Y(n669) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n119) );
  OAI21X1 U229 ( .A(n1037), .B(n1002), .C(n120), .Y(n670) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n120) );
  NAND3X1 U231 ( .A(n973), .B(n48), .C(n121), .Y(n112) );
  OAI21X1 U232 ( .A(n1038), .B(n1001), .C(n123), .Y(n671) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n123) );
  OAI21X1 U234 ( .A(n1039), .B(n1000), .C(n124), .Y(n672) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n124) );
  OAI21X1 U236 ( .A(n1040), .B(n1000), .C(n125), .Y(n673) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n125) );
  OAI21X1 U238 ( .A(n1041), .B(n1000), .C(n126), .Y(n674) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n126) );
  OAI21X1 U240 ( .A(n1042), .B(n1000), .C(n127), .Y(n675) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n127) );
  OAI21X1 U242 ( .A(n1043), .B(n1000), .C(n128), .Y(n676) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n128) );
  OAI21X1 U244 ( .A(n1044), .B(n1000), .C(n129), .Y(n677) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n129) );
  OAI21X1 U246 ( .A(n1045), .B(n1000), .C(n130), .Y(n678) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n130) );
  NAND3X1 U248 ( .A(n91), .B(n48), .C(n111), .Y(n122) );
  OAI21X1 U249 ( .A(n1030), .B(n999), .C(n132), .Y(n679) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n132) );
  OAI21X1 U251 ( .A(n1031), .B(n999), .C(n133), .Y(n680) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n133) );
  OAI21X1 U253 ( .A(n1032), .B(n999), .C(n134), .Y(n681) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n134) );
  OAI21X1 U255 ( .A(n1033), .B(n999), .C(n135), .Y(n682) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n135) );
  OAI21X1 U257 ( .A(n1034), .B(n999), .C(n136), .Y(n683) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n136) );
  OAI21X1 U259 ( .A(n1035), .B(n999), .C(n137), .Y(n684) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n137) );
  OAI21X1 U261 ( .A(n1036), .B(n999), .C(n138), .Y(n685) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n138) );
  OAI21X1 U263 ( .A(n1037), .B(n999), .C(n139), .Y(n686) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n139) );
  NAND3X1 U265 ( .A(n973), .B(n48), .C(n140), .Y(n131) );
  OAI21X1 U266 ( .A(n1038), .B(n998), .C(n142), .Y(n687) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n142) );
  OAI21X1 U268 ( .A(n1039), .B(n998), .C(n143), .Y(n688) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n143) );
  OAI21X1 U270 ( .A(n1040), .B(n998), .C(n144), .Y(n689) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n144) );
  OAI21X1 U272 ( .A(n1041), .B(n998), .C(n145), .Y(n690) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n145) );
  OAI21X1 U274 ( .A(n1042), .B(n998), .C(n146), .Y(n691) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n146) );
  OAI21X1 U276 ( .A(n1043), .B(n998), .C(n147), .Y(n692) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n147) );
  OAI21X1 U278 ( .A(n1044), .B(n998), .C(n148), .Y(n693) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n148) );
  OAI21X1 U280 ( .A(n1045), .B(n998), .C(n149), .Y(n694) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n149) );
  NAND3X1 U282 ( .A(n71), .B(n48), .C(n969), .Y(n141) );
  OAI21X1 U283 ( .A(n1030), .B(n997), .C(n152), .Y(n695) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n152) );
  OAI21X1 U285 ( .A(n1031), .B(n997), .C(n153), .Y(n696) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n153) );
  OAI21X1 U287 ( .A(n1032), .B(n997), .C(n154), .Y(n697) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n154) );
  OAI21X1 U289 ( .A(n1033), .B(n997), .C(n155), .Y(n698) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n155) );
  OAI21X1 U291 ( .A(n1034), .B(n997), .C(n156), .Y(n699) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n156) );
  OAI21X1 U293 ( .A(n1035), .B(n997), .C(n157), .Y(n700) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n157) );
  OAI21X1 U295 ( .A(n1036), .B(n997), .C(n158), .Y(n701) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n158) );
  OAI21X1 U297 ( .A(n1037), .B(n997), .C(n159), .Y(n702) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n159) );
  NAND3X1 U299 ( .A(n973), .B(n48), .C(n160), .Y(n151) );
  OAI21X1 U300 ( .A(n1038), .B(n996), .C(n162), .Y(n703) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n162) );
  OAI21X1 U302 ( .A(n1039), .B(n996), .C(n163), .Y(n704) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n163) );
  OAI21X1 U304 ( .A(n1040), .B(n996), .C(n164), .Y(n705) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n164) );
  OAI21X1 U306 ( .A(n1041), .B(n996), .C(n165), .Y(n706) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n165) );
  OAI21X1 U308 ( .A(n1042), .B(n996), .C(n166), .Y(n707) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n166) );
  OAI21X1 U310 ( .A(n1043), .B(n996), .C(n167), .Y(n708) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n167) );
  OAI21X1 U312 ( .A(n1044), .B(n996), .C(n168), .Y(n709) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n168) );
  OAI21X1 U314 ( .A(n1045), .B(n996), .C(n169), .Y(n710) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n169) );
  NAND3X1 U316 ( .A(n91), .B(n48), .C(n969), .Y(n161) );
  OAI21X1 U317 ( .A(n1030), .B(n995), .C(n171), .Y(n711) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n171) );
  OAI21X1 U319 ( .A(n1031), .B(n995), .C(n172), .Y(n712) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n172) );
  OAI21X1 U321 ( .A(n1032), .B(n995), .C(n173), .Y(n713) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n173) );
  OAI21X1 U323 ( .A(n1033), .B(n995), .C(n174), .Y(n714) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n174) );
  OAI21X1 U325 ( .A(n1034), .B(n995), .C(n175), .Y(n715) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n175) );
  OAI21X1 U327 ( .A(n1035), .B(n995), .C(n176), .Y(n716) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n176) );
  OAI21X1 U329 ( .A(n1036), .B(n995), .C(n177), .Y(n717) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n177) );
  OAI21X1 U331 ( .A(n1037), .B(n995), .C(n178), .Y(n718) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n178) );
  NAND3X1 U333 ( .A(n973), .B(n48), .C(n179), .Y(n170) );
  OAI21X1 U334 ( .A(n1038), .B(n994), .C(n181), .Y(n719) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n181) );
  OAI21X1 U336 ( .A(n1039), .B(n994), .C(n182), .Y(n720) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n182) );
  OAI21X1 U338 ( .A(n1040), .B(n994), .C(n183), .Y(n721) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n183) );
  OAI21X1 U340 ( .A(n1041), .B(n994), .C(n184), .Y(n722) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n184) );
  OAI21X1 U342 ( .A(n1042), .B(n994), .C(n185), .Y(n723) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n185) );
  OAI21X1 U344 ( .A(n1043), .B(n994), .C(n186), .Y(n724) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n186) );
  OAI21X1 U346 ( .A(n1044), .B(n994), .C(n187), .Y(n725) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n187) );
  OAI21X1 U348 ( .A(n1045), .B(n994), .C(n188), .Y(n726) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n188) );
  NAND3X1 U350 ( .A(n71), .B(n48), .C(n967), .Y(n180) );
  OAI21X1 U351 ( .A(n1030), .B(n993), .C(n191), .Y(n727) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n191) );
  OAI21X1 U353 ( .A(n1031), .B(n993), .C(n192), .Y(n728) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n192) );
  OAI21X1 U355 ( .A(n1032), .B(n993), .C(n193), .Y(n729) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n193) );
  OAI21X1 U357 ( .A(n1033), .B(n993), .C(n194), .Y(n730) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n194) );
  OAI21X1 U359 ( .A(n1034), .B(n993), .C(n195), .Y(n731) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n195) );
  OAI21X1 U361 ( .A(n1035), .B(n993), .C(n196), .Y(n732) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n196) );
  OAI21X1 U363 ( .A(n1036), .B(n993), .C(n197), .Y(n733) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n197) );
  OAI21X1 U365 ( .A(n1037), .B(n993), .C(n198), .Y(n734) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n198) );
  NAND3X1 U367 ( .A(n973), .B(n48), .C(n199), .Y(n190) );
  OAI21X1 U368 ( .A(n1038), .B(n992), .C(n201), .Y(n735) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n201) );
  OAI21X1 U370 ( .A(n1039), .B(n992), .C(n202), .Y(n736) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n202) );
  OAI21X1 U372 ( .A(n1040), .B(n992), .C(n203), .Y(n737) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n203) );
  OAI21X1 U374 ( .A(n1041), .B(n992), .C(n204), .Y(n738) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n204) );
  OAI21X1 U376 ( .A(n1042), .B(n992), .C(n205), .Y(n739) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n205) );
  OAI21X1 U378 ( .A(n1043), .B(n992), .C(n206), .Y(n740) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n206) );
  OAI21X1 U380 ( .A(n1044), .B(n992), .C(n207), .Y(n741) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n207) );
  OAI21X1 U382 ( .A(n1045), .B(n992), .C(n208), .Y(n742) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n208) );
  NAND3X1 U384 ( .A(n91), .B(n48), .C(n967), .Y(n200) );
  OAI21X1 U385 ( .A(n1030), .B(n991), .C(n210), .Y(n743) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n210) );
  OAI21X1 U387 ( .A(n1031), .B(n991), .C(n211), .Y(n744) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n211) );
  OAI21X1 U389 ( .A(n1032), .B(n991), .C(n212), .Y(n745) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n212) );
  OAI21X1 U391 ( .A(n1033), .B(n991), .C(n213), .Y(n746) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n213) );
  OAI21X1 U393 ( .A(n1034), .B(n991), .C(n214), .Y(n747) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n214) );
  OAI21X1 U395 ( .A(n1035), .B(n991), .C(n215), .Y(n748) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n215) );
  OAI21X1 U397 ( .A(n1036), .B(n991), .C(n216), .Y(n749) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n216) );
  OAI21X1 U399 ( .A(n1037), .B(n991), .C(n217), .Y(n750) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n217) );
  NAND3X1 U401 ( .A(n973), .B(n48), .C(n218), .Y(n209) );
  OAI21X1 U402 ( .A(n1038), .B(n990), .C(n220), .Y(n751) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n220) );
  OAI21X1 U404 ( .A(n1039), .B(n989), .C(n221), .Y(n752) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n221) );
  OAI21X1 U406 ( .A(n1040), .B(n989), .C(n222), .Y(n753) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n222) );
  OAI21X1 U408 ( .A(n1041), .B(n989), .C(n223), .Y(n754) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n223) );
  OAI21X1 U410 ( .A(n1042), .B(n989), .C(n224), .Y(n755) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n224) );
  OAI21X1 U412 ( .A(n1043), .B(n989), .C(n225), .Y(n756) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n225) );
  OAI21X1 U414 ( .A(n1044), .B(n989), .C(n226), .Y(n757) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n226) );
  OAI21X1 U416 ( .A(n1045), .B(n989), .C(n227), .Y(n758) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n227) );
  NAND3X1 U418 ( .A(n70), .B(n48), .C(n228), .Y(n219) );
  OAI21X1 U419 ( .A(n1030), .B(n988), .C(n230), .Y(n759) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n230) );
  OAI21X1 U421 ( .A(n1031), .B(n988), .C(n231), .Y(n760) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n231) );
  OAI21X1 U423 ( .A(n1032), .B(n988), .C(n232), .Y(n761) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n232) );
  OAI21X1 U425 ( .A(n1033), .B(n988), .C(n233), .Y(n762) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n233) );
  OAI21X1 U427 ( .A(n1034), .B(n988), .C(n234), .Y(n763) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n234) );
  OAI21X1 U429 ( .A(n1035), .B(n988), .C(n235), .Y(n764) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n235) );
  OAI21X1 U431 ( .A(n1036), .B(n988), .C(n236), .Y(n765) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n236) );
  OAI21X1 U433 ( .A(n1037), .B(n988), .C(n237), .Y(n766) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n237) );
  NAND3X1 U435 ( .A(n973), .B(n48), .C(n238), .Y(n229) );
  OAI21X1 U436 ( .A(n1038), .B(n987), .C(n240), .Y(n767) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n240) );
  OAI21X1 U438 ( .A(n1039), .B(n986), .C(n241), .Y(n768) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n241) );
  OAI21X1 U440 ( .A(n1040), .B(n986), .C(n242), .Y(n769) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n242) );
  OAI21X1 U442 ( .A(n1041), .B(n986), .C(n243), .Y(n770) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n243) );
  OAI21X1 U444 ( .A(n1042), .B(n986), .C(n244), .Y(n771) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n244) );
  OAI21X1 U446 ( .A(n1043), .B(n986), .C(n245), .Y(n772) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n245) );
  OAI21X1 U448 ( .A(n1044), .B(n986), .C(n246), .Y(n773) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n246) );
  OAI21X1 U450 ( .A(n1045), .B(n986), .C(n247), .Y(n774) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n247) );
  NAND3X1 U452 ( .A(n70), .B(n48), .C(n248), .Y(n239) );
  OAI21X1 U453 ( .A(n1030), .B(n985), .C(n251), .Y(n775) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n251) );
  OAI21X1 U455 ( .A(n1031), .B(n985), .C(n252), .Y(n776) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n252) );
  OAI21X1 U457 ( .A(n1032), .B(n985), .C(n253), .Y(n777) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n253) );
  OAI21X1 U459 ( .A(n1033), .B(n985), .C(n254), .Y(n778) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n254) );
  OAI21X1 U461 ( .A(n1034), .B(n985), .C(n255), .Y(n779) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n255) );
  OAI21X1 U463 ( .A(n1035), .B(n985), .C(n256), .Y(n780) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n256) );
  OAI21X1 U465 ( .A(n1036), .B(n985), .C(n257), .Y(n781) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n257) );
  OAI21X1 U467 ( .A(n1037), .B(n985), .C(n258), .Y(n782) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n258) );
  NAND3X1 U469 ( .A(n973), .B(n48), .C(n259), .Y(n250) );
  OAI21X1 U470 ( .A(n1038), .B(n984), .C(n261), .Y(n783) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n261) );
  OAI21X1 U472 ( .A(n1039), .B(n983), .C(n262), .Y(n784) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n262) );
  OAI21X1 U474 ( .A(n1040), .B(n983), .C(n263), .Y(n785) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n263) );
  OAI21X1 U476 ( .A(n1041), .B(n983), .C(n264), .Y(n786) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n264) );
  OAI21X1 U478 ( .A(n1042), .B(n983), .C(n265), .Y(n787) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n265) );
  OAI21X1 U480 ( .A(n1043), .B(n983), .C(n266), .Y(n788) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n266) );
  OAI21X1 U482 ( .A(n1044), .B(n983), .C(n267), .Y(n789) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n267) );
  OAI21X1 U484 ( .A(n1045), .B(n983), .C(n268), .Y(n790) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n268) );
  NAND3X1 U486 ( .A(n111), .B(n48), .C(n228), .Y(n260) );
  OAI21X1 U487 ( .A(n1030), .B(n982), .C(n270), .Y(n791) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n270) );
  OAI21X1 U489 ( .A(n1031), .B(n982), .C(n271), .Y(n792) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n271) );
  OAI21X1 U491 ( .A(n1032), .B(n982), .C(n272), .Y(n793) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n272) );
  OAI21X1 U493 ( .A(n1033), .B(n982), .C(n273), .Y(n794) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n273) );
  OAI21X1 U495 ( .A(n1034), .B(n982), .C(n274), .Y(n795) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n274) );
  OAI21X1 U497 ( .A(n1035), .B(n982), .C(n275), .Y(n796) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n275) );
  OAI21X1 U499 ( .A(n1036), .B(n982), .C(n276), .Y(n797) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n276) );
  OAI21X1 U501 ( .A(n1037), .B(n982), .C(n277), .Y(n798) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n277) );
  NAND3X1 U503 ( .A(n973), .B(n48), .C(n278), .Y(n269) );
  OAI21X1 U504 ( .A(n1038), .B(n981), .C(n280), .Y(n799) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n280) );
  OAI21X1 U506 ( .A(n1039), .B(n980), .C(n281), .Y(n800) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n281) );
  OAI21X1 U508 ( .A(n1040), .B(n980), .C(n282), .Y(n801) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n282) );
  OAI21X1 U510 ( .A(n1041), .B(n980), .C(n283), .Y(n802) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n283) );
  OAI21X1 U512 ( .A(n1042), .B(n980), .C(n284), .Y(n803) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n284) );
  OAI21X1 U514 ( .A(n1043), .B(n980), .C(n285), .Y(n804) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n285) );
  OAI21X1 U516 ( .A(n1044), .B(n980), .C(n286), .Y(n805) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n286) );
  OAI21X1 U518 ( .A(n1045), .B(n980), .C(n287), .Y(n806) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n287) );
  NAND3X1 U520 ( .A(n111), .B(n48), .C(n248), .Y(n279) );
  OAI21X1 U521 ( .A(n1030), .B(n979), .C(n291), .Y(n807) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n291) );
  OAI21X1 U523 ( .A(n1031), .B(n979), .C(n292), .Y(n808) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n292) );
  OAI21X1 U525 ( .A(n1032), .B(n979), .C(n293), .Y(n809) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n293) );
  OAI21X1 U527 ( .A(n1033), .B(n979), .C(n294), .Y(n810) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n294) );
  OAI21X1 U529 ( .A(n1034), .B(n979), .C(n295), .Y(n811) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n295) );
  OAI21X1 U531 ( .A(n1035), .B(n979), .C(n296), .Y(n812) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n296) );
  OAI21X1 U533 ( .A(n1036), .B(n979), .C(n297), .Y(n813) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n297) );
  OAI21X1 U535 ( .A(n1037), .B(n979), .C(n298), .Y(n814) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n298) );
  NAND3X1 U537 ( .A(n973), .B(n48), .C(n299), .Y(n290) );
  OAI21X1 U538 ( .A(n1038), .B(n978), .C(n301), .Y(n815) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n301) );
  OAI21X1 U540 ( .A(n1039), .B(n978), .C(n302), .Y(n816) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n302) );
  OAI21X1 U542 ( .A(n1040), .B(n978), .C(n303), .Y(n817) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n303) );
  OAI21X1 U544 ( .A(n1041), .B(n978), .C(n304), .Y(n818) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n304) );
  OAI21X1 U546 ( .A(n1042), .B(n978), .C(n305), .Y(n819) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n305) );
  OAI21X1 U548 ( .A(n1043), .B(n978), .C(n306), .Y(n820) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n306) );
  OAI21X1 U550 ( .A(n1044), .B(n978), .C(n307), .Y(n821) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n307) );
  OAI21X1 U552 ( .A(n1045), .B(n978), .C(n308), .Y(n822) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n308) );
  NAND3X1 U554 ( .A(n969), .B(n48), .C(n228), .Y(n300) );
  OAI21X1 U555 ( .A(n1030), .B(n977), .C(n310), .Y(n823) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n310) );
  OAI21X1 U557 ( .A(n1031), .B(n977), .C(n311), .Y(n824) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n311) );
  OAI21X1 U559 ( .A(n1032), .B(n977), .C(n312), .Y(n825) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n312) );
  OAI21X1 U561 ( .A(n1033), .B(n977), .C(n313), .Y(n826) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n313) );
  OAI21X1 U563 ( .A(n1034), .B(n977), .C(n314), .Y(n827) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n314) );
  OAI21X1 U565 ( .A(n1035), .B(n977), .C(n315), .Y(n828) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n315) );
  OAI21X1 U567 ( .A(n1036), .B(n977), .C(n316), .Y(n829) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n316) );
  OAI21X1 U569 ( .A(n1037), .B(n977), .C(n317), .Y(n830) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n317) );
  NAND3X1 U571 ( .A(n973), .B(n48), .C(n318), .Y(n309) );
  OAI21X1 U572 ( .A(n1038), .B(n976), .C(n320), .Y(n831) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n320) );
  OAI21X1 U574 ( .A(n1039), .B(n976), .C(n321), .Y(n832) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n321) );
  OAI21X1 U576 ( .A(n1040), .B(n976), .C(n322), .Y(n833) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n322) );
  OAI21X1 U578 ( .A(n1041), .B(n976), .C(n323), .Y(n834) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n323) );
  OAI21X1 U580 ( .A(n1042), .B(n976), .C(n324), .Y(n835) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n324) );
  OAI21X1 U582 ( .A(n1043), .B(n976), .C(n325), .Y(n836) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n325) );
  OAI21X1 U584 ( .A(n1044), .B(n976), .C(n326), .Y(n837) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n326) );
  OAI21X1 U586 ( .A(n1045), .B(n976), .C(n327), .Y(n838) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n327) );
  NAND3X1 U588 ( .A(n969), .B(n48), .C(n248), .Y(n319) );
  OAI21X1 U590 ( .A(n1030), .B(n975), .C(n330), .Y(n839) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n330) );
  OAI21X1 U592 ( .A(n1031), .B(n975), .C(n331), .Y(n840) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n331) );
  OAI21X1 U594 ( .A(n1032), .B(n975), .C(n332), .Y(n841) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n332) );
  OAI21X1 U596 ( .A(n1033), .B(n975), .C(n333), .Y(n842) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n333) );
  OAI21X1 U598 ( .A(n1034), .B(n975), .C(n334), .Y(n843) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n334) );
  OAI21X1 U600 ( .A(n1035), .B(n975), .C(n335), .Y(n844) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n335) );
  OAI21X1 U602 ( .A(n1036), .B(n975), .C(n336), .Y(n845) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n336) );
  OAI21X1 U604 ( .A(n1037), .B(n975), .C(n337), .Y(n846) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n337) );
  NAND3X1 U606 ( .A(n973), .B(n48), .C(n338), .Y(n329) );
  OAI21X1 U607 ( .A(n1038), .B(n974), .C(n340), .Y(n847) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n340) );
  OAI21X1 U609 ( .A(n1039), .B(n974), .C(n341), .Y(n848) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n341) );
  OAI21X1 U611 ( .A(n1040), .B(n974), .C(n342), .Y(n849) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n342) );
  OAI21X1 U613 ( .A(n1041), .B(n974), .C(n343), .Y(n850) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n343) );
  OAI21X1 U615 ( .A(n1042), .B(n974), .C(n344), .Y(n851) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n344) );
  OAI21X1 U617 ( .A(n1043), .B(n974), .C(n345), .Y(n852) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n345) );
  OAI21X1 U619 ( .A(n1044), .B(n974), .C(n346), .Y(n853) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n346) );
  OAI21X1 U621 ( .A(n1045), .B(n974), .C(n347), .Y(n854) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n347) );
  NAND3X1 U623 ( .A(n967), .B(n48), .C(n228), .Y(n339) );
  OAI21X1 U624 ( .A(n1030), .B(n8), .C(n349), .Y(n855) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n349) );
  OAI21X1 U626 ( .A(n1031), .B(n8), .C(n350), .Y(n856) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n350) );
  OAI21X1 U628 ( .A(n1032), .B(n8), .C(n351), .Y(n857) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n351) );
  OAI21X1 U630 ( .A(n1033), .B(n8), .C(n352), .Y(n858) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n352) );
  OAI21X1 U632 ( .A(n1034), .B(n8), .C(n353), .Y(n859) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n353) );
  OAI21X1 U634 ( .A(n1035), .B(n8), .C(n354), .Y(n860) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n354) );
  OAI21X1 U636 ( .A(n1036), .B(n8), .C(n355), .Y(n861) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n355) );
  OAI21X1 U638 ( .A(n1037), .B(n8), .C(n356), .Y(n862) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n356) );
  NOR2X1 U641 ( .A(n964), .B(\addr_1c<4> ), .Y(n59) );
  OAI21X1 U642 ( .A(n1038), .B(n972), .C(n359), .Y(n863) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n359) );
  OAI21X1 U644 ( .A(n1039), .B(n972), .C(n360), .Y(n864) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n360) );
  OAI21X1 U646 ( .A(n1040), .B(n972), .C(n361), .Y(n865) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n361) );
  OAI21X1 U648 ( .A(n1041), .B(n972), .C(n362), .Y(n866) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n362) );
  OAI21X1 U650 ( .A(n1042), .B(n972), .C(n363), .Y(n867) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n363) );
  OAI21X1 U652 ( .A(n1043), .B(n972), .C(n364), .Y(n868) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n364) );
  OAI21X1 U654 ( .A(n1044), .B(n972), .C(n365), .Y(n869) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n365) );
  OAI21X1 U656 ( .A(n1045), .B(n972), .C(n366), .Y(n870) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n366) );
  NAND3X1 U658 ( .A(n967), .B(n48), .C(n248), .Y(n358) );
  NOR3X1 U661 ( .A(n370), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n369) );
  NOR3X1 U662 ( .A(n371), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n368) );
  AOI21X1 U663 ( .A(n473), .B(n373), .C(n963), .Y(n1046) );
  OAI21X1 U665 ( .A(rd), .B(n374), .C(wr), .Y(n373) );
  NAND3X1 U667 ( .A(n375), .B(n1025), .C(n376), .Y(n374) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n376) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n375) );
  AOI21X1 U670 ( .A(n460), .B(n378), .C(n1016), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n380), .C(n4), .Y(n378) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n91), .C(\mem<0><1> ), .D(n248), .Y(n383) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n71), .C(\mem<2><1> ), .D(n228), .Y(n382) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n91), .C(\mem<4><1> ), .D(n248), .Y(n385) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n71), .C(\mem<6><1> ), .D(n228), .Y(n384) );
  AOI22X1 U678 ( .A(n288), .B(n893), .C(n249), .D(n933), .Y(n377) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n91), .C(\mem<12><1> ), .D(n248), .Y(
        n389) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n71), .C(\mem<14><1> ), .D(n228), .Y(
        n388) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n91), .C(\mem<8><1> ), .D(n248), .Y(n391) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n71), .C(\mem<10><1> ), .D(n228), .Y(
        n390) );
  AOI21X1 U685 ( .A(n448), .B(n393), .C(n1016), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n940), .B(n395), .C(n950), .Y(n393) );
  AOI21X1 U687 ( .A(n397), .B(n398), .C(n971), .Y(n396) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n91), .C(\mem<0><0> ), .D(n248), .Y(n398) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n71), .C(\mem<2><0> ), .D(n228), .Y(n397) );
  AOI21X1 U690 ( .A(n399), .B(n400), .C(n970), .Y(n394) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n91), .C(\mem<4><0> ), .D(n248), .Y(n400) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n71), .C(\mem<6><0> ), .D(n228), .Y(n399) );
  AOI22X1 U693 ( .A(n288), .B(n891), .C(n249), .D(n931), .Y(n392) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n91), .C(\mem<12><0> ), .D(n248), .Y(
        n404) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n71), .C(\mem<14><0> ), .D(n228), .Y(
        n403) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n91), .C(\mem<8><0> ), .D(n248), .Y(n406) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n71), .C(\mem<10><0> ), .D(n228), .Y(
        n405) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n407) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n199), .C(\mem<19><7> ), .D(n179), .Y(
        n414) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n160), .C(\mem<23><7> ), .D(n140), .Y(
        n413) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n121), .C(\mem<27><7> ), .D(n101), .Y(
        n411) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n81), .C(\mem<31><7> ), .D(n60), .Y(n410) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n357), .C(\mem<3><7> ), .D(n338), .Y(n419) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n318), .C(\mem<7><7> ), .D(n299), .Y(n418) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n278), .C(\mem<11><7> ), .D(n259), .Y(
        n416) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n238), .C(\mem<15><7> ), .D(n218), .Y(
        n415) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n420) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n199), .C(\mem<19><6> ), .D(n179), .Y(
        n427) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n160), .C(\mem<23><6> ), .D(n140), .Y(
        n426) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n121), .C(\mem<27><6> ), .D(n101), .Y(
        n424) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n81), .C(\mem<31><6> ), .D(n60), .Y(n423) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n357), .C(\mem<3><6> ), .D(n338), .Y(n432) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n318), .C(\mem<7><6> ), .D(n299), .Y(n431) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n278), .C(\mem<11><6> ), .D(n259), .Y(
        n429) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n238), .C(\mem<15><6> ), .D(n218), .Y(
        n428) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n433) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n199), .C(\mem<19><5> ), .D(n179), .Y(
        n440) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n160), .C(\mem<23><5> ), .D(n140), .Y(
        n439) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n121), .C(\mem<27><5> ), .D(n101), .Y(
        n437) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n81), .C(\mem<31><5> ), .D(n60), .Y(n436) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n357), .C(\mem<3><5> ), .D(n338), .Y(n445) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n318), .C(\mem<7><5> ), .D(n299), .Y(n444) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n278), .C(\mem<11><5> ), .D(n259), .Y(
        n442) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n238), .C(\mem<15><5> ), .D(n218), .Y(
        n441) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n446) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n199), .C(\mem<19><4> ), .D(n179), .Y(
        n453) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n160), .C(\mem<23><4> ), .D(n140), .Y(
        n452) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n121), .C(\mem<27><4> ), .D(n101), .Y(
        n450) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n81), .C(\mem<31><4> ), .D(n60), .Y(n449) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n357), .C(\mem<3><4> ), .D(n338), .Y(n458) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n318), .C(\mem<7><4> ), .D(n299), .Y(n457) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n278), .C(\mem<11><4> ), .D(n259), .Y(
        n455) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n238), .C(\mem<15><4> ), .D(n218), .Y(
        n454) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n459) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n199), .C(\mem<19><3> ), .D(n179), .Y(
        n466) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n160), .C(\mem<23><3> ), .D(n140), .Y(
        n465) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n121), .C(\mem<27><3> ), .D(n101), .Y(
        n463) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n81), .C(\mem<31><3> ), .D(n60), .Y(n462) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n357), .C(\mem<3><3> ), .D(n338), .Y(n471) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n318), .C(\mem<7><3> ), .D(n299), .Y(n470) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n278), .C(\mem<11><3> ), .D(n259), .Y(
        n468) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n238), .C(\mem<15><3> ), .D(n218), .Y(
        n467) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n472) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n199), .C(\mem<19><2> ), .D(n179), .Y(
        n479) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n160), .C(\mem<23><2> ), .D(n140), .Y(
        n478) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n121), .C(\mem<27><2> ), .D(n101), .Y(
        n476) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n81), .C(\mem<31><2> ), .D(n60), .Y(n475) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n357), .C(\mem<3><2> ), .D(n338), .Y(n484) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n318), .C(\mem<7><2> ), .D(n299), .Y(n483) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n278), .C(\mem<11><2> ), .D(n259), .Y(
        n481) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n238), .C(\mem<15><2> ), .D(n218), .Y(
        n480) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n485) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n199), .C(\mem<19><1> ), .D(n179), .Y(
        n492) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n160), .C(\mem<23><1> ), .D(n140), .Y(
        n491) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n121), .C(\mem<27><1> ), .D(n101), .Y(
        n489) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n81), .C(\mem<31><1> ), .D(n60), .Y(n488) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n357), .C(\mem<3><1> ), .D(n338), .Y(n497) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n318), .C(\mem<7><1> ), .D(n299), .Y(n496) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n278), .C(\mem<11><1> ), .D(n259), .Y(
        n494) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n238), .C(\mem<15><1> ), .D(n218), .Y(
        n493) );
  AOI21X1 U777 ( .A(n447), .B(n499), .C(n1016), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n939), .B(n501), .C(n949), .Y(n499) );
  AOI21X1 U779 ( .A(n503), .B(n504), .C(n971), .Y(n502) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n91), .C(\mem<0><7> ), .D(n248), .Y(n504) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n71), .C(\mem<2><7> ), .D(n228), .Y(n503) );
  AOI21X1 U782 ( .A(n505), .B(n506), .C(n970), .Y(n500) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n91), .C(\mem<4><7> ), .D(n248), .Y(n506) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n71), .C(\mem<6><7> ), .D(n228), .Y(n505) );
  AOI22X1 U785 ( .A(n288), .B(n889), .C(n249), .D(n929), .Y(n498) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n91), .C(\mem<12><7> ), .D(n248), .Y(
        n510) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n71), .C(\mem<14><7> ), .D(n228), .Y(
        n509) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n91), .C(\mem<8><7> ), .D(n248), .Y(n512) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n71), .C(\mem<10><7> ), .D(n228), .Y(
        n511) );
  AOI21X1 U792 ( .A(n435), .B(n514), .C(n1016), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n938), .B(n516), .C(n948), .Y(n514) );
  AOI21X1 U794 ( .A(n518), .B(n519), .C(n971), .Y(n517) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n91), .C(\mem<0><6> ), .D(n248), .Y(n519) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n71), .C(\mem<2><6> ), .D(n228), .Y(n518) );
  AOI21X1 U797 ( .A(n520), .B(n521), .C(n970), .Y(n515) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n91), .C(\mem<4><6> ), .D(n248), .Y(n521) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n71), .C(\mem<6><6> ), .D(n228), .Y(n520) );
  AOI22X1 U800 ( .A(n288), .B(n887), .C(n249), .D(n927), .Y(n513) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n91), .C(\mem<12><6> ), .D(n248), .Y(
        n525) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n71), .C(\mem<14><6> ), .D(n228), .Y(
        n524) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n91), .C(\mem<8><6> ), .D(n248), .Y(n527) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n71), .C(\mem<10><6> ), .D(n228), .Y(
        n526) );
  AOI21X1 U807 ( .A(n434), .B(n529), .C(n1016), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n937), .B(n531), .C(n947), .Y(n529) );
  AOI21X1 U809 ( .A(n533), .B(n534), .C(n971), .Y(n532) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n91), .C(\mem<0><5> ), .D(n248), .Y(n534) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n71), .C(\mem<2><5> ), .D(n228), .Y(n533) );
  AOI21X1 U812 ( .A(n535), .B(n536), .C(n970), .Y(n530) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n91), .C(\mem<4><5> ), .D(n248), .Y(n536) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n71), .C(\mem<6><5> ), .D(n228), .Y(n535) );
  AOI22X1 U815 ( .A(n288), .B(n885), .C(n249), .D(n925), .Y(n528) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n91), .C(\mem<12><5> ), .D(n248), .Y(
        n540) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n71), .C(\mem<14><5> ), .D(n228), .Y(
        n539) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n91), .C(\mem<8><5> ), .D(n248), .Y(n542) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n71), .C(\mem<10><5> ), .D(n228), .Y(
        n541) );
  AOI21X1 U822 ( .A(n422), .B(n544), .C(n1016), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n936), .B(n546), .C(n946), .Y(n544) );
  AOI21X1 U824 ( .A(n548), .B(n549), .C(n971), .Y(n547) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n91), .C(\mem<0><4> ), .D(n248), .Y(n549) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n71), .C(\mem<2><4> ), .D(n228), .Y(n548) );
  AOI21X1 U827 ( .A(n550), .B(n551), .C(n970), .Y(n545) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n91), .C(\mem<4><4> ), .D(n248), .Y(n551) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n71), .C(\mem<6><4> ), .D(n228), .Y(n550) );
  AOI22X1 U830 ( .A(n288), .B(n883), .C(n249), .D(n923), .Y(n543) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n91), .C(\mem<12><4> ), .D(n248), .Y(
        n555) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n71), .C(\mem<14><4> ), .D(n228), .Y(
        n554) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n91), .C(\mem<8><4> ), .D(n248), .Y(n557) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n71), .C(\mem<10><4> ), .D(n228), .Y(
        n556) );
  AOI21X1 U837 ( .A(n421), .B(n559), .C(n1016), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n935), .B(n561), .C(n945), .Y(n559) );
  AOI21X1 U839 ( .A(n563), .B(n564), .C(n971), .Y(n562) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n91), .C(\mem<0><3> ), .D(n248), .Y(n564) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n71), .C(\mem<2><3> ), .D(n228), .Y(n563) );
  AOI21X1 U842 ( .A(n565), .B(n566), .C(n970), .Y(n560) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n91), .C(\mem<4><3> ), .D(n248), .Y(n566) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n71), .C(\mem<6><3> ), .D(n228), .Y(n565) );
  AOI22X1 U845 ( .A(n288), .B(n881), .C(n249), .D(n921), .Y(n558) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n91), .C(\mem<12><3> ), .D(n248), .Y(
        n570) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n71), .C(\mem<14><3> ), .D(n228), .Y(
        n569) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n91), .C(\mem<8><3> ), .D(n248), .Y(n572) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n71), .C(\mem<10><3> ), .D(n228), .Y(
        n571) );
  AOI21X1 U852 ( .A(n409), .B(n574), .C(n1016), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n934), .B(n576), .C(n944), .Y(n574) );
  AOI21X1 U854 ( .A(n578), .B(n579), .C(n971), .Y(n577) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n91), .C(\mem<0><2> ), .D(n248), .Y(n579) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n71), .C(\mem<2><2> ), .D(n228), .Y(n578) );
  AOI21X1 U857 ( .A(n580), .B(n581), .C(n970), .Y(n575) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n91), .C(\mem<4><2> ), .D(n248), .Y(n581) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n71), .C(\mem<6><2> ), .D(n228), .Y(n580) );
  AOI22X1 U860 ( .A(n288), .B(n879), .C(n249), .D(n919), .Y(n573) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n91), .C(\mem<12><2> ), .D(n248), .Y(
        n585) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n71), .C(\mem<14><2> ), .D(n228), .Y(
        n584) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n91), .C(\mem<8><2> ), .D(n248), .Y(n587) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n71), .C(\mem<10><2> ), .D(n228), .Y(
        n586) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n588) );
  NOR2X1 U868 ( .A(n1029), .B(\addr_1c<4> ), .Y(n589) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n590) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n199), .C(\mem<19><0> ), .D(n179), .Y(
        n597) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n160), .C(\mem<23><0> ), .D(n140), .Y(
        n596) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n121), .C(\mem<27><0> ), .D(n101), .Y(
        n594) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n81), .C(\mem<31><0> ), .D(n60), .Y(n593) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n357), .C(\mem<3><0> ), .D(n338), .Y(n604) );
  NAND2X1 U877 ( .A(n1027), .B(n1028), .Y(n367) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n318), .C(\mem<7><0> ), .D(n299), .Y(n603) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1028), .Y(n328) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n278), .C(\mem<11><0> ), .D(n259), .Y(
        n601) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n238), .C(\mem<15><0> ), .D(n218), .Y(
        n600) );
  dff_203 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_202 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_185 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_186 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_187 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_188 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_189 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_190 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_191 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_192 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_193 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_194 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_195 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1012) );
  dff_196 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1012) );
  dff_197 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1012) );
  dff_169 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_170 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_171 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_172 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_173 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_174 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_175 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_176 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_177 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_178 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_179 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_180 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_181 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_182 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_183 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_184 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_153 \reg2[0]  ( .q(\data_out<0> ), .d(n1024), .clk(clk), .rst(n1012) );
  dff_154 \reg2[1]  ( .q(\data_out<1> ), .d(n1023), .clk(clk), .rst(n1012) );
  dff_155 \reg2[2]  ( .q(\data_out<2> ), .d(n1022), .clk(clk), .rst(n1012) );
  dff_156 \reg2[3]  ( .q(\data_out<3> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_157 \reg2[4]  ( .q(\data_out<4> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_158 \reg2[5]  ( .q(\data_out<5> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_159 \reg2[6]  ( .q(\data_out<6> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_160 \reg2[7]  ( .q(\data_out<7> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_161 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1012) );
  dff_162 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1012) );
  dff_163 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_164 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_165 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_166 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_167 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_168 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_201 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_200 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_199 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_198 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  INVX1 U2 ( .A(rd), .Y(n1015) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n371) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n357), .Y(n49) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1029) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1028) );
  INVX1 U7 ( .A(\addr_1c<1> ), .Y(n1027) );
  OR2X1 U8 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n370) );
  AND2X1 U23 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n598) );
  AND2X1 U24 ( .A(\addr_1c<3> ), .B(n1026), .Y(n599) );
  AND2X1 U25 ( .A(n249), .B(n965), .Y(n70) );
  AND2X1 U26 ( .A(n288), .B(n965), .Y(n111) );
  AND2X1 U27 ( .A(\addr_1c<0> ), .B(n1029), .Y(n605) );
  AND2X1 U28 ( .A(n1026), .B(n1029), .Y(n606) );
  INVX1 U29 ( .A(\addr_1c<0> ), .Y(n1026) );
  INVX1 U35 ( .A(wr1), .Y(n1025) );
  AND2X1 U36 ( .A(\addr_1c<2> ), .B(n1027), .Y(n288) );
  AND2X1 U37 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n249) );
  AND2X1 U38 ( .A(n599), .B(n249), .Y(n81) );
  AND2X1 U39 ( .A(n288), .B(n598), .Y(n101) );
  AND2X1 U40 ( .A(n288), .B(n599), .Y(n121) );
  AND2X1 U41 ( .A(n941), .B(n598), .Y(n140) );
  AND2X1 U42 ( .A(n941), .B(n599), .Y(n160) );
  AND2X1 U43 ( .A(n598), .B(n951), .Y(n179) );
  AND2X1 U44 ( .A(n599), .B(n951), .Y(n199) );
  AND2X1 U46 ( .A(n605), .B(n249), .Y(n218) );
  AND2X1 U47 ( .A(n249), .B(n606), .Y(n238) );
  AND2X1 U48 ( .A(n605), .B(n288), .Y(n259) );
  AND2X1 U49 ( .A(n288), .B(n606), .Y(n278) );
  AND2X1 U50 ( .A(n605), .B(n941), .Y(n299) );
  AND2X1 U51 ( .A(n941), .B(n606), .Y(n318) );
  OR2X1 U52 ( .A(n970), .B(n964), .Y(n968) );
  AND2X1 U53 ( .A(n605), .B(n951), .Y(n338) );
  OR2X1 U54 ( .A(n964), .B(n971), .Y(n966) );
  AND2X1 U55 ( .A(n49), .B(\mem<32><0> ), .Y(n395) );
  AND2X1 U56 ( .A(n49), .B(\mem<32><1> ), .Y(n380) );
  AND2X1 U57 ( .A(n49), .B(\mem<32><2> ), .Y(n576) );
  AND2X1 U58 ( .A(n49), .B(\mem<32><3> ), .Y(n561) );
  AND2X1 U59 ( .A(n49), .B(\mem<32><4> ), .Y(n546) );
  AND2X1 U60 ( .A(n49), .B(\mem<32><5> ), .Y(n531) );
  AND2X1 U61 ( .A(n49), .B(\mem<32><6> ), .Y(n516) );
  AND2X1 U62 ( .A(n49), .B(\mem<32><7> ), .Y(n501) );
  INVX1 U63 ( .A(rd1), .Y(n1016) );
  BUFX2 U64 ( .A(n961), .Y(n1010) );
  BUFX2 U65 ( .A(n961), .Y(n1009) );
  BUFX2 U66 ( .A(n960), .Y(n1007) );
  BUFX2 U67 ( .A(n960), .Y(n1006) );
  BUFX2 U68 ( .A(n959), .Y(n1004) );
  BUFX2 U69 ( .A(n959), .Y(n1003) );
  BUFX2 U70 ( .A(n958), .Y(n1001) );
  BUFX2 U71 ( .A(n958), .Y(n1000) );
  BUFX2 U72 ( .A(n957), .Y(n990) );
  BUFX2 U73 ( .A(n957), .Y(n989) );
  BUFX2 U74 ( .A(n956), .Y(n987) );
  BUFX2 U75 ( .A(n956), .Y(n986) );
  BUFX2 U76 ( .A(n955), .Y(n984) );
  BUFX2 U77 ( .A(n955), .Y(n983) );
  BUFX2 U78 ( .A(n954), .Y(n981) );
  BUFX2 U79 ( .A(n954), .Y(n980) );
  INVX1 U80 ( .A(\data_in_1c<0> ), .Y(n1030) );
  INVX1 U81 ( .A(\data_in_1c<1> ), .Y(n1031) );
  INVX1 U82 ( .A(\data_in_1c<2> ), .Y(n1032) );
  INVX1 U83 ( .A(\data_in_1c<3> ), .Y(n1033) );
  INVX1 U84 ( .A(\data_in_1c<4> ), .Y(n1034) );
  INVX1 U85 ( .A(\data_in_1c<5> ), .Y(n1035) );
  INVX1 U86 ( .A(\data_in_1c<6> ), .Y(n1036) );
  INVX1 U87 ( .A(\data_in_1c<7> ), .Y(n1037) );
  INVX1 U88 ( .A(\data_in_1c<8> ), .Y(n1038) );
  INVX1 U89 ( .A(\data_in_1c<9> ), .Y(n1039) );
  INVX1 U90 ( .A(\data_in_1c<10> ), .Y(n1040) );
  INVX1 U91 ( .A(\data_in_1c<11> ), .Y(n1041) );
  INVX1 U92 ( .A(\data_in_1c<12> ), .Y(n1042) );
  INVX1 U93 ( .A(\data_in_1c<13> ), .Y(n1043) );
  INVX1 U129 ( .A(\data_in_1c<14> ), .Y(n1044) );
  INVX1 U589 ( .A(\data_in_1c<15> ), .Y(n1045) );
  INVX1 U640 ( .A(wr), .Y(n1014) );
  INVX1 U659 ( .A(n590), .Y(n1024) );
  INVX1 U660 ( .A(n485), .Y(n1023) );
  INVX1 U664 ( .A(n472), .Y(n1022) );
  INVX1 U666 ( .A(n459), .Y(n1021) );
  INVX1 U672 ( .A(n446), .Y(n1020) );
  INVX1 U675 ( .A(n433), .Y(n1019) );
  INVX1 U679 ( .A(n420), .Y(n1018) );
  INVX1 U682 ( .A(n407), .Y(n1017) );
  INVX1 U694 ( .A(rst), .Y(n1013) );
  INVX2 U697 ( .A(n1013), .Y(n1012) );
  AND2X1 U701 ( .A(wr1), .B(n1013), .Y(n48) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n60), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n487), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n474), .B(n486), .Y(n10) );
  OR2X1 U761 ( .A(n522), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n507), .B(n508), .Y(n12) );
  OR2X1 U772 ( .A(n538), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n523), .B(n537), .Y(n14) );
  OR2X1 U789 ( .A(n567), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n552), .B(n553), .Y(n16) );
  OR2X1 U804 ( .A(n583), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n568), .B(n582), .Y(n18) );
  OR2X1 U819 ( .A(n871), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n591), .B(n592), .Y(n20) );
  OR2X1 U834 ( .A(n874), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n872), .B(n873), .Y(n22) );
  OR2X1 U849 ( .A(n877), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n875), .B(n876), .Y(n24) );
  OR2X1 U864 ( .A(n896), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n894), .B(n895), .Y(n26) );
  OR2X1 U875 ( .A(n899), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n897), .B(n898), .Y(n28) );
  OR2X1 U883 ( .A(n902), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n900), .B(n901), .Y(n30) );
  OR2X1 U885 ( .A(n905), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n903), .B(n904), .Y(n32) );
  OR2X1 U887 ( .A(n908), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n906), .B(n907), .Y(n34) );
  OR2X1 U889 ( .A(n911), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n909), .B(n910), .Y(n36) );
  OR2X1 U891 ( .A(n914), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n912), .B(n913), .Y(n38) );
  OR2X1 U893 ( .A(n917), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n915), .B(n916), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n48), .Y(n189) );
  AND2X1 U896 ( .A(n48), .B(n357), .Y(n289) );
  AND2X1 U897 ( .A(n941), .B(n943), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n941), .B(n942), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1046), .Y(err) );
  BUFX2 U906 ( .A(n573), .Y(n409) );
  BUFX2 U907 ( .A(n558), .Y(n421) );
  BUFX2 U908 ( .A(n543), .Y(n422) );
  BUFX2 U909 ( .A(n528), .Y(n434) );
  BUFX2 U910 ( .A(n513), .Y(n435) );
  BUFX2 U911 ( .A(n498), .Y(n447) );
  BUFX2 U912 ( .A(n392), .Y(n448) );
  BUFX2 U913 ( .A(n377), .Y(n460) );
  AND2X2 U914 ( .A(rd), .B(n374), .Y(n461) );
  INVX1 U915 ( .A(n461), .Y(n473) );
  INVX1 U916 ( .A(n602), .Y(n474) );
  INVX1 U917 ( .A(n601), .Y(n486) );
  INVX1 U918 ( .A(n600), .Y(n487) );
  INVX1 U919 ( .A(n495), .Y(n507) );
  INVX1 U920 ( .A(n494), .Y(n508) );
  INVX1 U921 ( .A(n493), .Y(n522) );
  INVX1 U922 ( .A(n482), .Y(n523) );
  INVX1 U923 ( .A(n481), .Y(n537) );
  INVX1 U924 ( .A(n480), .Y(n538) );
  INVX1 U925 ( .A(n469), .Y(n552) );
  INVX1 U926 ( .A(n468), .Y(n553) );
  INVX1 U927 ( .A(n467), .Y(n567) );
  INVX1 U928 ( .A(n456), .Y(n568) );
  INVX1 U929 ( .A(n455), .Y(n582) );
  INVX1 U930 ( .A(n454), .Y(n583) );
  INVX1 U931 ( .A(n443), .Y(n591) );
  INVX1 U932 ( .A(n442), .Y(n592) );
  INVX1 U933 ( .A(n441), .Y(n871) );
  INVX1 U934 ( .A(n430), .Y(n872) );
  INVX1 U935 ( .A(n429), .Y(n873) );
  INVX1 U936 ( .A(n428), .Y(n874) );
  INVX1 U937 ( .A(n417), .Y(n875) );
  INVX1 U938 ( .A(n416), .Y(n876) );
  INVX1 U939 ( .A(n415), .Y(n877) );
  AND2X2 U940 ( .A(n586), .B(n587), .Y(n878) );
  INVX1 U941 ( .A(n878), .Y(n879) );
  AND2X2 U942 ( .A(n571), .B(n572), .Y(n880) );
  INVX1 U943 ( .A(n880), .Y(n881) );
  AND2X2 U944 ( .A(n556), .B(n557), .Y(n882) );
  INVX1 U945 ( .A(n882), .Y(n883) );
  AND2X2 U946 ( .A(n541), .B(n542), .Y(n884) );
  INVX1 U947 ( .A(n884), .Y(n885) );
  AND2X2 U948 ( .A(n526), .B(n527), .Y(n886) );
  INVX1 U949 ( .A(n886), .Y(n887) );
  AND2X2 U950 ( .A(n511), .B(n512), .Y(n888) );
  INVX1 U951 ( .A(n888), .Y(n889) );
  AND2X2 U952 ( .A(n405), .B(n406), .Y(n890) );
  INVX1 U953 ( .A(n890), .Y(n891) );
  AND2X2 U954 ( .A(n390), .B(n391), .Y(n892) );
  INVX1 U955 ( .A(n892), .Y(n893) );
  INVX1 U956 ( .A(n595), .Y(n894) );
  INVX1 U957 ( .A(n594), .Y(n895) );
  INVX1 U958 ( .A(n593), .Y(n896) );
  INVX1 U959 ( .A(n490), .Y(n897) );
  INVX1 U960 ( .A(n489), .Y(n898) );
  INVX1 U961 ( .A(n488), .Y(n899) );
  INVX1 U962 ( .A(n477), .Y(n900) );
  INVX1 U963 ( .A(n476), .Y(n901) );
  INVX1 U964 ( .A(n475), .Y(n902) );
  INVX1 U965 ( .A(n464), .Y(n903) );
  INVX1 U966 ( .A(n463), .Y(n904) );
  INVX1 U967 ( .A(n462), .Y(n905) );
  INVX1 U968 ( .A(n451), .Y(n906) );
  INVX1 U969 ( .A(n450), .Y(n907) );
  INVX1 U970 ( .A(n449), .Y(n908) );
  INVX1 U971 ( .A(n438), .Y(n909) );
  INVX1 U972 ( .A(n437), .Y(n910) );
  INVX1 U973 ( .A(n436), .Y(n911) );
  INVX1 U974 ( .A(n425), .Y(n912) );
  INVX1 U975 ( .A(n424), .Y(n913) );
  INVX1 U976 ( .A(n423), .Y(n914) );
  INVX1 U977 ( .A(n412), .Y(n915) );
  INVX1 U978 ( .A(n411), .Y(n916) );
  INVX1 U979 ( .A(n410), .Y(n917) );
  AND2X2 U980 ( .A(n584), .B(n585), .Y(n918) );
  INVX1 U981 ( .A(n918), .Y(n919) );
  AND2X2 U982 ( .A(n569), .B(n570), .Y(n920) );
  INVX1 U983 ( .A(n920), .Y(n921) );
  AND2X2 U984 ( .A(n554), .B(n555), .Y(n922) );
  INVX1 U985 ( .A(n922), .Y(n923) );
  AND2X2 U986 ( .A(n539), .B(n540), .Y(n924) );
  INVX1 U987 ( .A(n924), .Y(n925) );
  AND2X2 U988 ( .A(n524), .B(n525), .Y(n926) );
  INVX1 U989 ( .A(n926), .Y(n927) );
  AND2X2 U990 ( .A(n509), .B(n510), .Y(n928) );
  INVX1 U991 ( .A(n928), .Y(n929) );
  AND2X2 U992 ( .A(n403), .B(n404), .Y(n930) );
  INVX1 U993 ( .A(n930), .Y(n931) );
  AND2X2 U994 ( .A(n388), .B(n389), .Y(n932) );
  INVX1 U995 ( .A(n932), .Y(n933) );
  BUFX2 U996 ( .A(n575), .Y(n934) );
  BUFX2 U997 ( .A(n560), .Y(n935) );
  BUFX2 U998 ( .A(n545), .Y(n936) );
  BUFX2 U999 ( .A(n530), .Y(n937) );
  BUFX2 U1000 ( .A(n515), .Y(n938) );
  BUFX2 U1001 ( .A(n500), .Y(n939) );
  BUFX2 U1002 ( .A(n394), .Y(n940) );
  INVX1 U1003 ( .A(n970), .Y(n941) );
  INVX1 U1004 ( .A(n385), .Y(n942) );
  INVX1 U1005 ( .A(n384), .Y(n943) );
  BUFX2 U1006 ( .A(n328), .Y(n970) );
  BUFX2 U1007 ( .A(n577), .Y(n944) );
  BUFX2 U1008 ( .A(n562), .Y(n945) );
  BUFX2 U1009 ( .A(n547), .Y(n946) );
  BUFX2 U1010 ( .A(n532), .Y(n947) );
  BUFX2 U1011 ( .A(n517), .Y(n948) );
  BUFX2 U1012 ( .A(n502), .Y(n949) );
  BUFX2 U1013 ( .A(n396), .Y(n950) );
  INVX1 U1014 ( .A(n971), .Y(n951) );
  INVX1 U1015 ( .A(n383), .Y(n952) );
  INVX1 U1016 ( .A(n382), .Y(n953) );
  BUFX2 U1017 ( .A(n367), .Y(n971) );
  BUFX2 U1018 ( .A(n358), .Y(n972) );
  BUFX2 U1019 ( .A(n339), .Y(n974) );
  BUFX2 U1020 ( .A(n329), .Y(n975) );
  BUFX2 U1021 ( .A(n319), .Y(n976) );
  BUFX2 U1022 ( .A(n309), .Y(n977) );
  BUFX2 U1023 ( .A(n300), .Y(n978) );
  BUFX2 U1024 ( .A(n290), .Y(n979) );
  BUFX2 U1025 ( .A(n269), .Y(n982) );
  BUFX2 U1026 ( .A(n250), .Y(n985) );
  BUFX2 U1027 ( .A(n229), .Y(n988) );
  BUFX2 U1028 ( .A(n209), .Y(n991) );
  BUFX2 U1029 ( .A(n200), .Y(n992) );
  BUFX2 U1030 ( .A(n190), .Y(n993) );
  BUFX2 U1031 ( .A(n180), .Y(n994) );
  BUFX2 U1032 ( .A(n170), .Y(n995) );
  BUFX2 U1033 ( .A(n161), .Y(n996) );
  BUFX2 U1034 ( .A(n151), .Y(n997) );
  BUFX2 U1035 ( .A(n141), .Y(n998) );
  BUFX2 U1036 ( .A(n131), .Y(n999) );
  BUFX2 U1037 ( .A(n112), .Y(n1002) );
  BUFX2 U1038 ( .A(n92), .Y(n1005) );
  BUFX2 U1039 ( .A(n72), .Y(n1008) );
  BUFX2 U1040 ( .A(n59), .Y(n973) );
  AND2X1 U1041 ( .A(n249), .B(n598), .Y(n60) );
  BUFX2 U1042 ( .A(n39), .Y(n1011) );
  BUFX2 U1043 ( .A(n279), .Y(n954) );
  BUFX2 U1044 ( .A(n260), .Y(n955) );
  BUFX2 U1045 ( .A(n239), .Y(n956) );
  BUFX2 U1046 ( .A(n219), .Y(n957) );
  BUFX2 U1047 ( .A(n122), .Y(n958) );
  BUFX2 U1048 ( .A(n102), .Y(n959) );
  BUFX2 U1049 ( .A(n82), .Y(n960) );
  BUFX2 U1050 ( .A(n61), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  INVX1 U1053 ( .A(n965), .Y(n964) );
  AND2X1 U1054 ( .A(n368), .B(n369), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n951), .B(n606), .Y(n357) );
endmodule


module final_memory_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1838, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1046), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1047), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1048), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1049), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1050), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1051), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1052), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1053), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1054), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1055), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1056), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1057), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1058), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1059), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1060), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1061), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1062), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1063), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1064), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1065), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1066), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1067), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1068), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1069), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1070), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1071), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1072), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1073), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1074), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1075), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1076), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1077), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1078), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1079), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1080), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1081), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1082), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1083), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1085), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1086), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1087), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1088), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1089), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1090), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1091), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1092), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1093), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1094), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1095), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1096), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1097), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1098), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1099), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1100), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1101), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1102), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1103), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1104), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1105), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1106), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1107), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1108), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1109), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1110), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1111), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1112), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1113), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1114), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1115), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1116), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1117), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1118), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1119), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1120), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1121), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1122), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1123), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1124), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1125), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1126), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1127), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1128), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1129), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1130), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1131), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1132), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1133), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1134), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1135), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1136), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1137), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1138), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1139), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1140), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1141), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1142), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1143), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1144), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1145), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1146), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1147), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1148), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1149), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1150), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1151), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1152), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1153), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1154), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1155), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1156), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1157), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1166), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1167), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1168), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1169), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1170), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1171), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1172), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1173), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1174), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1175), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1176), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1177), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1178), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1179), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1180), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1181), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1182), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1183), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1184), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1185), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1186), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1187), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1188), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1189), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1190), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1191), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1192), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1193), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1194), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1195), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1196), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1197), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1198), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1199), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1200), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1201), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1202), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1203), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1204), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1205), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1214), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1215), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1216), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1217), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1218), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1219), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1220), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1221), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1222), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1223), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1224), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1225), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1226), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1227), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1228), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1229), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1230), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1231), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1232), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1233), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1234), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1235), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1236), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1238), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1239), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1240), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1241), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1242), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1243), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1244), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1245), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1246), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1247), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1248), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1249), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1250), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1251), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1252), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1253), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1254), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1255), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1256), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1257), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1258), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1259), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1260), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1261), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1262), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1263), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1264), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1265), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1266), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1267), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1268), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1269), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1270), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1271), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1272), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1273), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1274), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1275), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1276), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1277), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1278), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1279), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1280), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1281), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1282), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1283), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1284), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1285), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1286), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1287), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1288), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1289), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1290), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1291), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1292), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1294), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1295), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1296), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1297), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1298), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1299), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1300), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1301), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1302), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1303), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1304), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1305), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1306), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1307), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1308), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1309), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1477), .B(n1476), .Y(n1478) );
  AND2X2 U10 ( .A(n1472), .B(n1471), .Y(n1473) );
  AND2X2 U11 ( .A(n1466), .B(n1465), .Y(n1467) );
  AND2X2 U12 ( .A(n1461), .B(n1460), .Y(n1462) );
  AND2X2 U13 ( .A(n1455), .B(n1454), .Y(n1456) );
  AND2X2 U14 ( .A(n1450), .B(n1449), .Y(n1451) );
  AND2X2 U15 ( .A(n1444), .B(n1443), .Y(n1445) );
  AND2X2 U16 ( .A(n1439), .B(n1438), .Y(n1440) );
  AND2X2 U17 ( .A(n1433), .B(n1432), .Y(n1434) );
  AND2X2 U18 ( .A(n1428), .B(n1427), .Y(n1429) );
  AND2X2 U19 ( .A(n1422), .B(n1421), .Y(n1423) );
  AND2X2 U20 ( .A(n1417), .B(n1416), .Y(n1418) );
  AND2X2 U21 ( .A(n1411), .B(n1410), .Y(n1412) );
  AND2X2 U22 ( .A(n1406), .B(n1405), .Y(n1407) );
  AND2X2 U30 ( .A(n1326), .B(n1026), .Y(n1631) );
  AND2X2 U31 ( .A(n1325), .B(n1026), .Y(n1786) );
  AND2X2 U32 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1651) );
  AND2X2 U33 ( .A(n1325), .B(\addr_1c<0> ), .Y(n1806) );
  AND2X2 U34 ( .A(n1320), .B(n1319), .Y(n1321) );
  AND2X2 U45 ( .A(n1313), .B(n1312), .Y(n1314) );
  NOR3X1 U94 ( .A(n1022), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1023), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1038), .C(n1836), .Y(n1309) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1836) );
  OAI21X1 U98 ( .A(n1011), .B(n1039), .C(n1835), .Y(n1308) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1835) );
  OAI21X1 U100 ( .A(n1011), .B(n1040), .C(n1834), .Y(n1307) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1834) );
  OAI21X1 U102 ( .A(n1011), .B(n1041), .C(n1833), .Y(n1306) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1833) );
  OAI21X1 U104 ( .A(n1011), .B(n1042), .C(n1832), .Y(n1305) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1832) );
  OAI21X1 U106 ( .A(n1011), .B(n1043), .C(n1831), .Y(n1304) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1831) );
  OAI21X1 U108 ( .A(n1011), .B(n1044), .C(n1830), .Y(n1303) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1830) );
  OAI21X1 U110 ( .A(n1011), .B(n1045), .C(n1829), .Y(n1302) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1829) );
  NAND3X1 U112 ( .A(n1828), .B(n1827), .C(n965), .Y(n1837) );
  OAI21X1 U113 ( .A(n6), .B(n1030), .C(n1826), .Y(n1301) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1826) );
  OAI21X1 U115 ( .A(n6), .B(n1031), .C(n1825), .Y(n1300) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1825) );
  OAI21X1 U117 ( .A(n6), .B(n1032), .C(n1824), .Y(n1299) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1824) );
  OAI21X1 U119 ( .A(n6), .B(n1033), .C(n1823), .Y(n1298) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1823) );
  OAI21X1 U121 ( .A(n6), .B(n1034), .C(n1822), .Y(n1297) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1822) );
  OAI21X1 U123 ( .A(n6), .B(n1035), .C(n1821), .Y(n1296) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1821) );
  OAI21X1 U125 ( .A(n6), .B(n1036), .C(n1820), .Y(n1295) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1820) );
  OAI21X1 U127 ( .A(n6), .B(n1037), .C(n1819), .Y(n1294) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1819) );
  OAI21X1 U130 ( .A(n1038), .B(n1010), .C(n1815), .Y(n1293) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1815) );
  OAI21X1 U132 ( .A(n1039), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1814) );
  OAI21X1 U134 ( .A(n1040), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1813) );
  OAI21X1 U136 ( .A(n1041), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1812) );
  OAI21X1 U138 ( .A(n1042), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1811) );
  OAI21X1 U140 ( .A(n1043), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1810) );
  OAI21X1 U142 ( .A(n1044), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1809) );
  OAI21X1 U144 ( .A(n1045), .B(n1009), .C(n1808), .Y(n1286) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1808) );
  NAND3X1 U146 ( .A(n1807), .B(n1828), .C(n1806), .Y(n1816) );
  OAI21X1 U147 ( .A(n1030), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1804) );
  OAI21X1 U149 ( .A(n1031), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1803) );
  OAI21X1 U151 ( .A(n1032), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1802) );
  OAI21X1 U153 ( .A(n1033), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1801) );
  OAI21X1 U155 ( .A(n1034), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1800) );
  OAI21X1 U157 ( .A(n1035), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1799) );
  OAI21X1 U159 ( .A(n1036), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1798) );
  OAI21X1 U161 ( .A(n1037), .B(n1008), .C(n1797), .Y(n1278) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1797) );
  NAND3X1 U163 ( .A(n973), .B(n1828), .C(n1796), .Y(n1805) );
  OAI21X1 U164 ( .A(n1038), .B(n1007), .C(n1794), .Y(n1277) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1794) );
  OAI21X1 U166 ( .A(n1039), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1793) );
  OAI21X1 U168 ( .A(n1040), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1792) );
  OAI21X1 U170 ( .A(n1041), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1791) );
  OAI21X1 U172 ( .A(n1042), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1790) );
  OAI21X1 U174 ( .A(n1043), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1789) );
  OAI21X1 U176 ( .A(n1044), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1788) );
  OAI21X1 U178 ( .A(n1045), .B(n1006), .C(n1787), .Y(n1270) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1787) );
  NAND3X1 U180 ( .A(n1807), .B(n1828), .C(n1786), .Y(n1795) );
  OAI21X1 U181 ( .A(n1030), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1784) );
  OAI21X1 U183 ( .A(n1031), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1783) );
  OAI21X1 U185 ( .A(n1032), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1782) );
  OAI21X1 U187 ( .A(n1033), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1781) );
  OAI21X1 U189 ( .A(n1034), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1780) );
  OAI21X1 U191 ( .A(n1035), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1779) );
  OAI21X1 U193 ( .A(n1036), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1778) );
  OAI21X1 U195 ( .A(n1037), .B(n1005), .C(n1777), .Y(n1262) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1777) );
  NAND3X1 U197 ( .A(n973), .B(n1828), .C(n1776), .Y(n1785) );
  OAI21X1 U198 ( .A(n1038), .B(n1004), .C(n1774), .Y(n1261) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1774) );
  OAI21X1 U200 ( .A(n1039), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1773) );
  OAI21X1 U202 ( .A(n1040), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1772) );
  OAI21X1 U204 ( .A(n1041), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1771) );
  OAI21X1 U206 ( .A(n1042), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1770) );
  OAI21X1 U208 ( .A(n1043), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1769) );
  OAI21X1 U210 ( .A(n1044), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1768) );
  OAI21X1 U212 ( .A(n1045), .B(n1003), .C(n1767), .Y(n1254) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1767) );
  NAND3X1 U214 ( .A(n1806), .B(n1828), .C(n1766), .Y(n1775) );
  OAI21X1 U215 ( .A(n1030), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1764) );
  OAI21X1 U217 ( .A(n1031), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1763) );
  OAI21X1 U219 ( .A(n1032), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1762) );
  OAI21X1 U221 ( .A(n1033), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1761) );
  OAI21X1 U223 ( .A(n1034), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1760) );
  OAI21X1 U225 ( .A(n1035), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1759) );
  OAI21X1 U227 ( .A(n1036), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1758) );
  OAI21X1 U229 ( .A(n1037), .B(n1002), .C(n1757), .Y(n1246) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1757) );
  NAND3X1 U231 ( .A(n973), .B(n1828), .C(n1756), .Y(n1765) );
  OAI21X1 U232 ( .A(n1038), .B(n1001), .C(n1754), .Y(n1245) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1754) );
  OAI21X1 U234 ( .A(n1039), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1753) );
  OAI21X1 U236 ( .A(n1040), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1752) );
  OAI21X1 U238 ( .A(n1041), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1751) );
  OAI21X1 U240 ( .A(n1042), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1750) );
  OAI21X1 U242 ( .A(n1043), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1749) );
  OAI21X1 U244 ( .A(n1044), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1748) );
  OAI21X1 U246 ( .A(n1045), .B(n1000), .C(n1747), .Y(n1238) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1747) );
  NAND3X1 U248 ( .A(n1786), .B(n1828), .C(n1766), .Y(n1755) );
  OAI21X1 U249 ( .A(n1030), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1745) );
  OAI21X1 U251 ( .A(n1031), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1744) );
  OAI21X1 U253 ( .A(n1032), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1743) );
  OAI21X1 U255 ( .A(n1033), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1742) );
  OAI21X1 U257 ( .A(n1034), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1741) );
  OAI21X1 U259 ( .A(n1035), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1740) );
  OAI21X1 U261 ( .A(n1036), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1739) );
  OAI21X1 U263 ( .A(n1037), .B(n999), .C(n1738), .Y(n1230) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1738) );
  NAND3X1 U265 ( .A(n973), .B(n1828), .C(n1737), .Y(n1746) );
  OAI21X1 U266 ( .A(n1038), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1735) );
  OAI21X1 U268 ( .A(n1039), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1734) );
  OAI21X1 U270 ( .A(n1040), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1733) );
  OAI21X1 U272 ( .A(n1041), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1732) );
  OAI21X1 U274 ( .A(n1042), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1731) );
  OAI21X1 U276 ( .A(n1043), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1730) );
  OAI21X1 U278 ( .A(n1044), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1729) );
  OAI21X1 U280 ( .A(n1045), .B(n998), .C(n1728), .Y(n1222) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1728) );
  NAND3X1 U282 ( .A(n1806), .B(n1828), .C(n969), .Y(n1736) );
  OAI21X1 U283 ( .A(n1030), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1726) );
  OAI21X1 U285 ( .A(n1031), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1725) );
  OAI21X1 U287 ( .A(n1032), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1724) );
  OAI21X1 U289 ( .A(n1033), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1723) );
  OAI21X1 U291 ( .A(n1034), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1722) );
  OAI21X1 U293 ( .A(n1035), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1721) );
  OAI21X1 U295 ( .A(n1036), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1720) );
  OAI21X1 U297 ( .A(n1037), .B(n997), .C(n1719), .Y(n1214) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1719) );
  NAND3X1 U299 ( .A(n973), .B(n1828), .C(n1718), .Y(n1727) );
  OAI21X1 U300 ( .A(n1038), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1716) );
  OAI21X1 U302 ( .A(n1039), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1715) );
  OAI21X1 U304 ( .A(n1040), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1714) );
  OAI21X1 U306 ( .A(n1041), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1713) );
  OAI21X1 U308 ( .A(n1042), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1712) );
  OAI21X1 U310 ( .A(n1043), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1711) );
  OAI21X1 U312 ( .A(n1044), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1710) );
  OAI21X1 U314 ( .A(n1045), .B(n996), .C(n1709), .Y(n1206) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1709) );
  NAND3X1 U316 ( .A(n1786), .B(n1828), .C(n969), .Y(n1717) );
  OAI21X1 U317 ( .A(n1030), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1707) );
  OAI21X1 U319 ( .A(n1031), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1706) );
  OAI21X1 U321 ( .A(n1032), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1705) );
  OAI21X1 U323 ( .A(n1033), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1704) );
  OAI21X1 U325 ( .A(n1034), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1703) );
  OAI21X1 U327 ( .A(n1035), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1702) );
  OAI21X1 U329 ( .A(n1036), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1701) );
  OAI21X1 U331 ( .A(n1037), .B(n995), .C(n1700), .Y(n1198) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1700) );
  NAND3X1 U333 ( .A(n973), .B(n1828), .C(n1699), .Y(n1708) );
  OAI21X1 U334 ( .A(n1038), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1697) );
  OAI21X1 U336 ( .A(n1039), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1696) );
  OAI21X1 U338 ( .A(n1040), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1695) );
  OAI21X1 U340 ( .A(n1041), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1694) );
  OAI21X1 U342 ( .A(n1042), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1693) );
  OAI21X1 U344 ( .A(n1043), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1692) );
  OAI21X1 U346 ( .A(n1044), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1691) );
  OAI21X1 U348 ( .A(n1045), .B(n994), .C(n1690), .Y(n1190) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1690) );
  NAND3X1 U350 ( .A(n1806), .B(n1828), .C(n967), .Y(n1698) );
  OAI21X1 U351 ( .A(n1030), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1688) );
  OAI21X1 U353 ( .A(n1031), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1687) );
  OAI21X1 U355 ( .A(n1032), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1686) );
  OAI21X1 U357 ( .A(n1033), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1685) );
  OAI21X1 U359 ( .A(n1034), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1684) );
  OAI21X1 U361 ( .A(n1035), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1683) );
  OAI21X1 U363 ( .A(n1036), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1682) );
  OAI21X1 U365 ( .A(n1037), .B(n993), .C(n1681), .Y(n1182) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1681) );
  NAND3X1 U367 ( .A(n973), .B(n1828), .C(n1680), .Y(n1689) );
  OAI21X1 U368 ( .A(n1038), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1678) );
  OAI21X1 U370 ( .A(n1039), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1677) );
  OAI21X1 U372 ( .A(n1040), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1676) );
  OAI21X1 U374 ( .A(n1041), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1675) );
  OAI21X1 U376 ( .A(n1042), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1674) );
  OAI21X1 U378 ( .A(n1043), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1673) );
  OAI21X1 U380 ( .A(n1044), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1672) );
  OAI21X1 U382 ( .A(n1045), .B(n992), .C(n1671), .Y(n1174) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1671) );
  NAND3X1 U384 ( .A(n1786), .B(n1828), .C(n967), .Y(n1679) );
  OAI21X1 U385 ( .A(n1030), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1669) );
  OAI21X1 U387 ( .A(n1031), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1668) );
  OAI21X1 U389 ( .A(n1032), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1667) );
  OAI21X1 U391 ( .A(n1033), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1666) );
  OAI21X1 U393 ( .A(n1034), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1665) );
  OAI21X1 U395 ( .A(n1035), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1664) );
  OAI21X1 U397 ( .A(n1036), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1663) );
  OAI21X1 U399 ( .A(n1037), .B(n991), .C(n1662), .Y(n1166) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1662) );
  NAND3X1 U401 ( .A(n973), .B(n1828), .C(n1661), .Y(n1670) );
  OAI21X1 U402 ( .A(n1038), .B(n990), .C(n1659), .Y(n1165) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1659) );
  OAI21X1 U404 ( .A(n1039), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1658) );
  OAI21X1 U406 ( .A(n1040), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1657) );
  OAI21X1 U408 ( .A(n1041), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1656) );
  OAI21X1 U410 ( .A(n1042), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1655) );
  OAI21X1 U412 ( .A(n1043), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1654) );
  OAI21X1 U414 ( .A(n1044), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1653) );
  OAI21X1 U416 ( .A(n1045), .B(n989), .C(n1652), .Y(n1158) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1652) );
  NAND3X1 U418 ( .A(n1807), .B(n1828), .C(n1651), .Y(n1660) );
  OAI21X1 U419 ( .A(n1030), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1649) );
  OAI21X1 U421 ( .A(n1031), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1648) );
  OAI21X1 U423 ( .A(n1032), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1647) );
  OAI21X1 U425 ( .A(n1033), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1646) );
  OAI21X1 U427 ( .A(n1034), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1645) );
  OAI21X1 U429 ( .A(n1035), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1644) );
  OAI21X1 U431 ( .A(n1036), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1643) );
  OAI21X1 U433 ( .A(n1037), .B(n988), .C(n1642), .Y(n1150) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1642) );
  NAND3X1 U435 ( .A(n973), .B(n1828), .C(n1641), .Y(n1650) );
  OAI21X1 U436 ( .A(n1038), .B(n987), .C(n1639), .Y(n1149) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1639) );
  OAI21X1 U438 ( .A(n1039), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1638) );
  OAI21X1 U440 ( .A(n1040), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1637) );
  OAI21X1 U442 ( .A(n1041), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1636) );
  OAI21X1 U444 ( .A(n1042), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1635) );
  OAI21X1 U446 ( .A(n1043), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1634) );
  OAI21X1 U448 ( .A(n1044), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1633) );
  OAI21X1 U450 ( .A(n1045), .B(n986), .C(n1632), .Y(n1142) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1632) );
  NAND3X1 U452 ( .A(n1807), .B(n1828), .C(n1631), .Y(n1640) );
  OAI21X1 U453 ( .A(n1030), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1628) );
  OAI21X1 U455 ( .A(n1031), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1627) );
  OAI21X1 U457 ( .A(n1032), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1626) );
  OAI21X1 U459 ( .A(n1033), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1625) );
  OAI21X1 U461 ( .A(n1034), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1624) );
  OAI21X1 U463 ( .A(n1035), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1623) );
  OAI21X1 U465 ( .A(n1036), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1622) );
  OAI21X1 U467 ( .A(n1037), .B(n985), .C(n1621), .Y(n1134) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1621) );
  NAND3X1 U469 ( .A(n973), .B(n1828), .C(n1620), .Y(n1629) );
  OAI21X1 U470 ( .A(n1038), .B(n984), .C(n1618), .Y(n1133) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1618) );
  OAI21X1 U472 ( .A(n1039), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1617) );
  OAI21X1 U474 ( .A(n1040), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1616) );
  OAI21X1 U476 ( .A(n1041), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1615) );
  OAI21X1 U478 ( .A(n1042), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1614) );
  OAI21X1 U480 ( .A(n1043), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1613) );
  OAI21X1 U482 ( .A(n1044), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1612) );
  OAI21X1 U484 ( .A(n1045), .B(n983), .C(n1611), .Y(n1126) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1611) );
  NAND3X1 U486 ( .A(n1766), .B(n1828), .C(n1651), .Y(n1619) );
  OAI21X1 U487 ( .A(n1030), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1609) );
  OAI21X1 U489 ( .A(n1031), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1608) );
  OAI21X1 U491 ( .A(n1032), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1607) );
  OAI21X1 U493 ( .A(n1033), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1606) );
  OAI21X1 U495 ( .A(n1034), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1605) );
  OAI21X1 U497 ( .A(n1035), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1604) );
  OAI21X1 U499 ( .A(n1036), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1603) );
  OAI21X1 U501 ( .A(n1037), .B(n982), .C(n1602), .Y(n1118) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1602) );
  NAND3X1 U503 ( .A(n973), .B(n1828), .C(n1601), .Y(n1610) );
  OAI21X1 U504 ( .A(n1038), .B(n981), .C(n1599), .Y(n1117) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1599) );
  OAI21X1 U506 ( .A(n1039), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1598) );
  OAI21X1 U508 ( .A(n1040), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1597) );
  OAI21X1 U510 ( .A(n1041), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1596) );
  OAI21X1 U512 ( .A(n1042), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1595) );
  OAI21X1 U514 ( .A(n1043), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1594) );
  OAI21X1 U516 ( .A(n1044), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1593) );
  OAI21X1 U518 ( .A(n1045), .B(n980), .C(n1592), .Y(n1110) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1592) );
  NAND3X1 U520 ( .A(n1766), .B(n1828), .C(n1631), .Y(n1600) );
  OAI21X1 U521 ( .A(n1030), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1589) );
  OAI21X1 U523 ( .A(n1031), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1588) );
  OAI21X1 U525 ( .A(n1032), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1587) );
  OAI21X1 U527 ( .A(n1033), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1586) );
  OAI21X1 U529 ( .A(n1034), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1585) );
  OAI21X1 U531 ( .A(n1035), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1584) );
  OAI21X1 U533 ( .A(n1036), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1583) );
  OAI21X1 U535 ( .A(n1037), .B(n979), .C(n1582), .Y(n1102) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1582) );
  NAND3X1 U537 ( .A(n973), .B(n1828), .C(n1581), .Y(n1590) );
  OAI21X1 U538 ( .A(n1038), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1579) );
  OAI21X1 U540 ( .A(n1039), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1578) );
  OAI21X1 U542 ( .A(n1040), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1577) );
  OAI21X1 U544 ( .A(n1041), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1576) );
  OAI21X1 U546 ( .A(n1042), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1575) );
  OAI21X1 U548 ( .A(n1043), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1574) );
  OAI21X1 U550 ( .A(n1044), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1573) );
  OAI21X1 U552 ( .A(n1045), .B(n978), .C(n1572), .Y(n1094) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1572) );
  NAND3X1 U554 ( .A(n969), .B(n1828), .C(n1651), .Y(n1580) );
  OAI21X1 U555 ( .A(n1030), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1570) );
  OAI21X1 U557 ( .A(n1031), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1569) );
  OAI21X1 U559 ( .A(n1032), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1568) );
  OAI21X1 U561 ( .A(n1033), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1567) );
  OAI21X1 U563 ( .A(n1034), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1566) );
  OAI21X1 U565 ( .A(n1035), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1565) );
  OAI21X1 U567 ( .A(n1036), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1564) );
  OAI21X1 U569 ( .A(n1037), .B(n977), .C(n1563), .Y(n1086) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1563) );
  NAND3X1 U571 ( .A(n973), .B(n1828), .C(n1562), .Y(n1571) );
  OAI21X1 U572 ( .A(n1038), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1560) );
  OAI21X1 U574 ( .A(n1039), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1559) );
  OAI21X1 U576 ( .A(n1040), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1558) );
  OAI21X1 U578 ( .A(n1041), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1557) );
  OAI21X1 U580 ( .A(n1042), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1556) );
  OAI21X1 U582 ( .A(n1043), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1555) );
  OAI21X1 U584 ( .A(n1044), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1554) );
  OAI21X1 U586 ( .A(n1045), .B(n976), .C(n1553), .Y(n1078) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1553) );
  NAND3X1 U588 ( .A(n969), .B(n1828), .C(n1631), .Y(n1561) );
  OAI21X1 U590 ( .A(n1030), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1550) );
  OAI21X1 U592 ( .A(n1031), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1549) );
  OAI21X1 U594 ( .A(n1032), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1548) );
  OAI21X1 U596 ( .A(n1033), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1547) );
  OAI21X1 U598 ( .A(n1034), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1546) );
  OAI21X1 U600 ( .A(n1035), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1545) );
  OAI21X1 U602 ( .A(n1036), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1544) );
  OAI21X1 U604 ( .A(n1037), .B(n975), .C(n1543), .Y(n1070) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1543) );
  NAND3X1 U606 ( .A(n973), .B(n1828), .C(n1542), .Y(n1551) );
  OAI21X1 U607 ( .A(n1038), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1540) );
  OAI21X1 U609 ( .A(n1039), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1539) );
  OAI21X1 U611 ( .A(n1040), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1538) );
  OAI21X1 U613 ( .A(n1041), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1537) );
  OAI21X1 U615 ( .A(n1042), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1536) );
  OAI21X1 U617 ( .A(n1043), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1535) );
  OAI21X1 U619 ( .A(n1044), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1534) );
  OAI21X1 U621 ( .A(n1045), .B(n974), .C(n1533), .Y(n1062) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1533) );
  NAND3X1 U623 ( .A(n967), .B(n1828), .C(n1651), .Y(n1541) );
  OAI21X1 U624 ( .A(n1030), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1532) );
  OAI21X1 U626 ( .A(n1031), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1531) );
  OAI21X1 U628 ( .A(n1032), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1530) );
  OAI21X1 U630 ( .A(n1033), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1529) );
  OAI21X1 U632 ( .A(n1034), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1528) );
  OAI21X1 U634 ( .A(n1035), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1527) );
  OAI21X1 U636 ( .A(n1036), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1526) );
  OAI21X1 U638 ( .A(n1037), .B(n8), .C(n1525), .Y(n1054) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1525) );
  NOR2X1 U641 ( .A(n964), .B(\addr_1c<4> ), .Y(n1818) );
  OAI21X1 U642 ( .A(n1038), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1522) );
  OAI21X1 U644 ( .A(n1039), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1521) );
  OAI21X1 U646 ( .A(n1040), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1520) );
  OAI21X1 U648 ( .A(n1041), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1519) );
  OAI21X1 U650 ( .A(n1042), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1518) );
  OAI21X1 U652 ( .A(n1043), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1517) );
  OAI21X1 U654 ( .A(n1044), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1516) );
  OAI21X1 U656 ( .A(n1045), .B(n972), .C(n1515), .Y(n1046) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1515) );
  NAND3X1 U658 ( .A(n967), .B(n1828), .C(n1631), .Y(n1523) );
  NOR3X1 U661 ( .A(n1511), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1512) );
  NOR3X1 U662 ( .A(n1510), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1513) );
  AOI21X1 U663 ( .A(n461), .B(n1509), .C(n963), .Y(n1838) );
  OAI21X1 U665 ( .A(rd), .B(n1508), .C(wr), .Y(n1509) );
  NAND3X1 U667 ( .A(n1507), .B(n1025), .C(n1506), .Y(n1508) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1506) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1507) );
  AOI21X1 U670 ( .A(n448), .B(n1504), .C(n1024), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1503), .C(n4), .Y(n1504) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1786), .C(\mem<0><1> ), .D(n1631), .Y(
        n1501) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1806), .C(\mem<2><1> ), .D(n1651), .Y(
        n1502) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1786), .C(\mem<4><1> ), .D(n1631), .Y(
        n1499) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1806), .C(\mem<6><1> ), .D(n1651), .Y(
        n1500) );
  AOI22X1 U678 ( .A(n1591), .B(n892), .C(n1630), .D(n932), .Y(n1505) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1786), .C(\mem<12><1> ), .D(n1631), .Y(
        n1497) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1806), .C(\mem<14><1> ), .D(n1651), .Y(
        n1498) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1786), .C(\mem<8><1> ), .D(n1631), .Y(
        n1495) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1806), .C(\mem<10><1> ), .D(n1651), .Y(
        n1496) );
  AOI21X1 U685 ( .A(n447), .B(n1493), .C(n1024), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1491), .C(n950), .Y(n1493) );
  AOI21X1 U687 ( .A(n1489), .B(n1488), .C(n971), .Y(n1490) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1786), .C(\mem<0><0> ), .D(n1631), .Y(
        n1488) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1806), .C(\mem<2><0> ), .D(n1651), .Y(
        n1489) );
  AOI21X1 U690 ( .A(n1487), .B(n1486), .C(n970), .Y(n1492) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1786), .C(\mem<4><0> ), .D(n1631), .Y(
        n1486) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1806), .C(\mem<6><0> ), .D(n1651), .Y(
        n1487) );
  AOI22X1 U693 ( .A(n1591), .B(n890), .C(n1630), .D(n930), .Y(n1494) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1786), .C(\mem<12><0> ), .D(n1631), .Y(
        n1484) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1806), .C(\mem<14><0> ), .D(n1651), .Y(
        n1485) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1786), .C(\mem<8><0> ), .D(n1631), .Y(
        n1482) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1806), .C(\mem<10><0> ), .D(n1651), .Y(
        n1483) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1481) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1680), .C(\mem<19><7> ), .D(n1699), .Y(
        n1476) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1718), .C(\mem<23><7> ), .D(n1737), .Y(
        n1477) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1756), .C(\mem<27><7> ), .D(n1776), .Y(
        n1479) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1796), .C(\mem<31><7> ), .D(n1817), .Y(
        n1480) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1524), .C(\mem<3><7> ), .D(n1542), .Y(
        n1471) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1562), .C(\mem<7><7> ), .D(n1581), .Y(
        n1472) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1601), .C(\mem<11><7> ), .D(n1620), .Y(
        n1474) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1641), .C(\mem<15><7> ), .D(n1661), .Y(
        n1475) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1470) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1680), .C(\mem<19><6> ), .D(n1699), .Y(
        n1465) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1718), .C(\mem<23><6> ), .D(n1737), .Y(
        n1466) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1756), .C(\mem<27><6> ), .D(n1776), .Y(
        n1468) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1796), .C(\mem<31><6> ), .D(n1817), .Y(
        n1469) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1524), .C(\mem<3><6> ), .D(n1542), .Y(
        n1460) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1562), .C(\mem<7><6> ), .D(n1581), .Y(
        n1461) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1601), .C(\mem<11><6> ), .D(n1620), .Y(
        n1463) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1641), .C(\mem<15><6> ), .D(n1661), .Y(
        n1464) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1459) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1680), .C(\mem<19><5> ), .D(n1699), .Y(
        n1454) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1718), .C(\mem<23><5> ), .D(n1737), .Y(
        n1455) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1756), .C(\mem<27><5> ), .D(n1776), .Y(
        n1457) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1796), .C(\mem<31><5> ), .D(n1817), .Y(
        n1458) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1524), .C(\mem<3><5> ), .D(n1542), .Y(
        n1449) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1562), .C(\mem<7><5> ), .D(n1581), .Y(
        n1450) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1601), .C(\mem<11><5> ), .D(n1620), .Y(
        n1452) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1641), .C(\mem<15><5> ), .D(n1661), .Y(
        n1453) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1448) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1680), .C(\mem<19><4> ), .D(n1699), .Y(
        n1443) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1718), .C(\mem<23><4> ), .D(n1737), .Y(
        n1444) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1756), .C(\mem<27><4> ), .D(n1776), .Y(
        n1446) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1796), .C(\mem<31><4> ), .D(n1817), .Y(
        n1447) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1524), .C(\mem<3><4> ), .D(n1542), .Y(
        n1438) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1562), .C(\mem<7><4> ), .D(n1581), .Y(
        n1439) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1601), .C(\mem<11><4> ), .D(n1620), .Y(
        n1441) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1641), .C(\mem<15><4> ), .D(n1661), .Y(
        n1442) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1437) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1680), .C(\mem<19><3> ), .D(n1699), .Y(
        n1432) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1718), .C(\mem<23><3> ), .D(n1737), .Y(
        n1433) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1756), .C(\mem<27><3> ), .D(n1776), .Y(
        n1435) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1796), .C(\mem<31><3> ), .D(n1817), .Y(
        n1436) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1524), .C(\mem<3><3> ), .D(n1542), .Y(
        n1427) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1562), .C(\mem<7><3> ), .D(n1581), .Y(
        n1428) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1601), .C(\mem<11><3> ), .D(n1620), .Y(
        n1430) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1641), .C(\mem<15><3> ), .D(n1661), .Y(
        n1431) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1426) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1680), .C(\mem<19><2> ), .D(n1699), .Y(
        n1421) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1718), .C(\mem<23><2> ), .D(n1737), .Y(
        n1422) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1756), .C(\mem<27><2> ), .D(n1776), .Y(
        n1424) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1796), .C(\mem<31><2> ), .D(n1817), .Y(
        n1425) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1524), .C(\mem<3><2> ), .D(n1542), .Y(
        n1416) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1562), .C(\mem<7><2> ), .D(n1581), .Y(
        n1417) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1601), .C(\mem<11><2> ), .D(n1620), .Y(
        n1419) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1641), .C(\mem<15><2> ), .D(n1661), .Y(
        n1420) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1415) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1680), .C(\mem<19><1> ), .D(n1699), .Y(
        n1410) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1718), .C(\mem<23><1> ), .D(n1737), .Y(
        n1411) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1756), .C(\mem<27><1> ), .D(n1776), .Y(
        n1413) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1796), .C(\mem<31><1> ), .D(n1817), .Y(
        n1414) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1524), .C(\mem<3><1> ), .D(n1542), .Y(
        n1405) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1562), .C(\mem<7><1> ), .D(n1581), .Y(
        n1406) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1601), .C(\mem<11><1> ), .D(n1620), .Y(
        n1408) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1641), .C(\mem<15><1> ), .D(n1661), .Y(
        n1409) );
  AOI21X1 U777 ( .A(n435), .B(n1403), .C(n1024), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1401), .C(n949), .Y(n1403) );
  AOI21X1 U779 ( .A(n1399), .B(n1398), .C(n971), .Y(n1400) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1786), .C(\mem<0><7> ), .D(n1631), .Y(
        n1398) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1806), .C(\mem<2><7> ), .D(n1651), .Y(
        n1399) );
  AOI21X1 U782 ( .A(n1397), .B(n1396), .C(n970), .Y(n1402) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1786), .C(\mem<4><7> ), .D(n1631), .Y(
        n1396) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1806), .C(\mem<6><7> ), .D(n1651), .Y(
        n1397) );
  AOI22X1 U785 ( .A(n1591), .B(n888), .C(n1630), .D(n928), .Y(n1404) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1786), .C(\mem<12><7> ), .D(n1631), .Y(
        n1394) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1806), .C(\mem<14><7> ), .D(n1651), .Y(
        n1395) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1786), .C(\mem<8><7> ), .D(n1631), .Y(
        n1392) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1806), .C(\mem<10><7> ), .D(n1651), .Y(
        n1393) );
  AOI21X1 U792 ( .A(n434), .B(n1390), .C(n1024), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1388), .C(n948), .Y(n1390) );
  AOI21X1 U794 ( .A(n1386), .B(n1385), .C(n971), .Y(n1387) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1786), .C(\mem<0><6> ), .D(n1631), .Y(
        n1385) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1806), .C(\mem<2><6> ), .D(n1651), .Y(
        n1386) );
  AOI21X1 U797 ( .A(n1384), .B(n1383), .C(n970), .Y(n1389) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1786), .C(\mem<4><6> ), .D(n1631), .Y(
        n1383) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1806), .C(\mem<6><6> ), .D(n1651), .Y(
        n1384) );
  AOI22X1 U800 ( .A(n1591), .B(n886), .C(n1630), .D(n926), .Y(n1391) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1786), .C(\mem<12><6> ), .D(n1631), .Y(
        n1381) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1806), .C(\mem<14><6> ), .D(n1651), .Y(
        n1382) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1786), .C(\mem<8><6> ), .D(n1631), .Y(
        n1379) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1806), .C(\mem<10><6> ), .D(n1651), .Y(
        n1380) );
  AOI21X1 U807 ( .A(n422), .B(n1377), .C(n1024), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1375), .C(n947), .Y(n1377) );
  AOI21X1 U809 ( .A(n1373), .B(n1372), .C(n971), .Y(n1374) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1786), .C(\mem<0><5> ), .D(n1631), .Y(
        n1372) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1806), .C(\mem<2><5> ), .D(n1651), .Y(
        n1373) );
  AOI21X1 U812 ( .A(n1371), .B(n1370), .C(n970), .Y(n1376) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1786), .C(\mem<4><5> ), .D(n1631), .Y(
        n1370) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1806), .C(\mem<6><5> ), .D(n1651), .Y(
        n1371) );
  AOI22X1 U815 ( .A(n1591), .B(n884), .C(n1630), .D(n924), .Y(n1378) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1786), .C(\mem<12><5> ), .D(n1631), .Y(
        n1368) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1806), .C(\mem<14><5> ), .D(n1651), .Y(
        n1369) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1786), .C(\mem<8><5> ), .D(n1631), .Y(
        n1366) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1806), .C(\mem<10><5> ), .D(n1651), .Y(
        n1367) );
  AOI21X1 U822 ( .A(n421), .B(n1364), .C(n1024), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1362), .C(n946), .Y(n1364) );
  AOI21X1 U824 ( .A(n1360), .B(n1359), .C(n971), .Y(n1361) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1786), .C(\mem<0><4> ), .D(n1631), .Y(
        n1359) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1806), .C(\mem<2><4> ), .D(n1651), .Y(
        n1360) );
  AOI21X1 U827 ( .A(n1358), .B(n1357), .C(n970), .Y(n1363) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1786), .C(\mem<4><4> ), .D(n1631), .Y(
        n1357) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1806), .C(\mem<6><4> ), .D(n1651), .Y(
        n1358) );
  AOI22X1 U830 ( .A(n1591), .B(n882), .C(n1630), .D(n922), .Y(n1365) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1786), .C(\mem<12><4> ), .D(n1631), .Y(
        n1355) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1806), .C(\mem<14><4> ), .D(n1651), .Y(
        n1356) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1786), .C(\mem<8><4> ), .D(n1631), .Y(
        n1353) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1806), .C(\mem<10><4> ), .D(n1651), .Y(
        n1354) );
  AOI21X1 U837 ( .A(n409), .B(n1351), .C(n1024), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1349), .C(n945), .Y(n1351) );
  AOI21X1 U839 ( .A(n1347), .B(n1346), .C(n971), .Y(n1348) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1786), .C(\mem<0><3> ), .D(n1631), .Y(
        n1346) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1806), .C(\mem<2><3> ), .D(n1651), .Y(
        n1347) );
  AOI21X1 U842 ( .A(n1345), .B(n1344), .C(n970), .Y(n1350) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1786), .C(\mem<4><3> ), .D(n1631), .Y(
        n1344) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1806), .C(\mem<6><3> ), .D(n1651), .Y(
        n1345) );
  AOI22X1 U845 ( .A(n1591), .B(n880), .C(n1630), .D(n920), .Y(n1352) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1786), .C(\mem<12><3> ), .D(n1631), .Y(
        n1342) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1806), .C(\mem<14><3> ), .D(n1651), .Y(
        n1343) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1786), .C(\mem<8><3> ), .D(n1631), .Y(
        n1340) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1806), .C(\mem<10><3> ), .D(n1651), .Y(
        n1341) );
  AOI21X1 U852 ( .A(n408), .B(n1338), .C(n1024), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1336), .C(n944), .Y(n1338) );
  AOI21X1 U854 ( .A(n1334), .B(n1333), .C(n971), .Y(n1335) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1786), .C(\mem<0><2> ), .D(n1631), .Y(
        n1333) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1806), .C(\mem<2><2> ), .D(n1651), .Y(
        n1334) );
  AOI21X1 U857 ( .A(n1332), .B(n1331), .C(n970), .Y(n1337) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1786), .C(\mem<4><2> ), .D(n1631), .Y(
        n1331) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1806), .C(\mem<6><2> ), .D(n1651), .Y(
        n1332) );
  AOI22X1 U860 ( .A(n1591), .B(n878), .C(n1630), .D(n918), .Y(n1339) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1786), .C(\mem<12><2> ), .D(n1631), .Y(
        n1329) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1806), .C(\mem<14><2> ), .D(n1651), .Y(
        n1330) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1786), .C(\mem<8><2> ), .D(n1631), .Y(
        n1327) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1806), .C(\mem<10><2> ), .D(n1651), .Y(
        n1328) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1326) );
  NOR2X1 U868 ( .A(n1029), .B(\addr_1c<4> ), .Y(n1325) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1324) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1680), .C(\mem<19><0> ), .D(n1699), .Y(
        n1319) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1718), .C(\mem<23><0> ), .D(n1737), .Y(
        n1320) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1756), .C(\mem<27><0> ), .D(n1776), .Y(
        n1322) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1796), .C(\mem<31><0> ), .D(n1817), .Y(
        n1323) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1524), .C(\mem<3><0> ), .D(n1542), .Y(
        n1312) );
  NAND2X1 U877 ( .A(n1027), .B(n1028), .Y(n1514) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1562), .C(\mem<7><0> ), .D(n1581), .Y(
        n1313) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1028), .Y(n1552) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1601), .C(\mem<11><0> ), .D(n1620), .Y(
        n1315) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1641), .C(\mem<15><0> ), .D(n1661), .Y(
        n1316) );
  dff_152 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_151 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_150 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_149 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_148 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_147 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_146 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_145 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_144 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_143 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_142 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_141 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_140 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1012) );
  dff_139 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1012) );
  dff_138 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1012) );
  dff_137 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_136 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_135 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_134 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_133 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_132 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_131 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_130 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_129 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_128 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_127 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_126 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_125 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_124 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_123 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_122 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_121 \reg2[0]  ( .q(\data_out<0> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_120 \reg2[1]  ( .q(\data_out<1> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_119 \reg2[2]  ( .q(\data_out<2> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_118 \reg2[3]  ( .q(\data_out<3> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_117 \reg2[4]  ( .q(\data_out<4> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_116 \reg2[5]  ( .q(\data_out<5> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_115 \reg2[6]  ( .q(\data_out<6> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_114 \reg2[7]  ( .q(\data_out<7> ), .d(n1014), .clk(clk), .rst(n1012) );
  dff_113 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1012) );
  dff_112 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1012) );
  dff_111 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_110 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_109 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_108 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_107 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_106 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_105 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_104 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_103 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_102 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  INVX1 U2 ( .A(rd), .Y(n1023) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1510) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n1524), .Y(n1827) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1029) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1028) );
  OR2X1 U7 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1511) );
  AND2X1 U8 ( .A(n1630), .B(n965), .Y(n1807) );
  AND2X1 U23 ( .A(n1591), .B(n965), .Y(n1766) );
  INVX1 U24 ( .A(\addr_1c<0> ), .Y(n1026) );
  AND2X1 U25 ( .A(n1026), .B(n1029), .Y(n1310) );
  AND2X1 U26 ( .A(\addr_1c<0> ), .B(n1029), .Y(n1311) );
  AND2X1 U27 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1318) );
  AND2X1 U28 ( .A(\addr_1c<3> ), .B(n1026), .Y(n1317) );
  INVX1 U29 ( .A(\addr_1c<1> ), .Y(n1027) );
  INVX1 U35 ( .A(wr1), .Y(n1025) );
  AND2X1 U36 ( .A(n1591), .B(n1318), .Y(n1776) );
  AND2X1 U37 ( .A(n1591), .B(n1317), .Y(n1756) );
  AND2X1 U38 ( .A(n940), .B(n1318), .Y(n1737) );
  AND2X1 U39 ( .A(n940), .B(n1317), .Y(n1718) );
  AND2X1 U40 ( .A(n1318), .B(n951), .Y(n1699) );
  AND2X1 U41 ( .A(n1317), .B(n951), .Y(n1680) );
  AND2X1 U42 ( .A(n1311), .B(n1591), .Y(n1620) );
  AND2X1 U43 ( .A(n1591), .B(n1310), .Y(n1601) );
  AND2X1 U44 ( .A(n1311), .B(n940), .Y(n1581) );
  AND2X1 U46 ( .A(n940), .B(n1310), .Y(n1562) );
  OR2X1 U47 ( .A(n970), .B(n964), .Y(n968) );
  AND2X1 U48 ( .A(n1311), .B(n951), .Y(n1542) );
  OR2X1 U49 ( .A(n964), .B(n971), .Y(n966) );
  AND2X1 U50 ( .A(n1630), .B(n1310), .Y(n1641) );
  AND2X1 U51 ( .A(n1311), .B(n1630), .Y(n1661) );
  AND2X1 U52 ( .A(n1317), .B(n1630), .Y(n1796) );
  AND2X1 U53 ( .A(\addr_1c<2> ), .B(n1027), .Y(n1591) );
  AND2X1 U54 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1630) );
  BUFX2 U55 ( .A(n961), .Y(n1010) );
  BUFX2 U56 ( .A(n961), .Y(n1009) );
  BUFX2 U57 ( .A(n960), .Y(n1007) );
  BUFX2 U58 ( .A(n960), .Y(n1006) );
  BUFX2 U59 ( .A(n959), .Y(n1004) );
  BUFX2 U60 ( .A(n959), .Y(n1003) );
  BUFX2 U61 ( .A(n958), .Y(n1001) );
  BUFX2 U62 ( .A(n958), .Y(n1000) );
  BUFX2 U63 ( .A(n957), .Y(n990) );
  BUFX2 U64 ( .A(n957), .Y(n989) );
  BUFX2 U65 ( .A(n956), .Y(n987) );
  BUFX2 U66 ( .A(n956), .Y(n986) );
  BUFX2 U67 ( .A(n955), .Y(n984) );
  BUFX2 U68 ( .A(n955), .Y(n983) );
  BUFX2 U69 ( .A(n954), .Y(n981) );
  BUFX2 U70 ( .A(n954), .Y(n980) );
  INVX1 U71 ( .A(\data_in_1c<0> ), .Y(n1030) );
  INVX1 U72 ( .A(\data_in_1c<1> ), .Y(n1031) );
  INVX1 U73 ( .A(\data_in_1c<2> ), .Y(n1032) );
  INVX1 U74 ( .A(\data_in_1c<3> ), .Y(n1033) );
  INVX1 U75 ( .A(\data_in_1c<4> ), .Y(n1034) );
  INVX1 U76 ( .A(\data_in_1c<5> ), .Y(n1035) );
  INVX1 U77 ( .A(\data_in_1c<6> ), .Y(n1036) );
  INVX1 U78 ( .A(\data_in_1c<7> ), .Y(n1037) );
  INVX1 U79 ( .A(\data_in_1c<8> ), .Y(n1038) );
  INVX1 U80 ( .A(\data_in_1c<9> ), .Y(n1039) );
  INVX1 U81 ( .A(\data_in_1c<10> ), .Y(n1040) );
  INVX1 U82 ( .A(\data_in_1c<11> ), .Y(n1041) );
  INVX1 U83 ( .A(\data_in_1c<12> ), .Y(n1042) );
  INVX1 U84 ( .A(\data_in_1c<13> ), .Y(n1043) );
  INVX1 U85 ( .A(\data_in_1c<14> ), .Y(n1044) );
  INVX1 U86 ( .A(\data_in_1c<15> ), .Y(n1045) );
  AND2X1 U87 ( .A(n1827), .B(\mem<32><0> ), .Y(n1491) );
  AND2X1 U88 ( .A(n1827), .B(\mem<32><1> ), .Y(n1503) );
  AND2X1 U89 ( .A(n1827), .B(\mem<32><2> ), .Y(n1336) );
  AND2X1 U90 ( .A(n1827), .B(\mem<32><3> ), .Y(n1349) );
  AND2X1 U91 ( .A(n1827), .B(\mem<32><4> ), .Y(n1362) );
  AND2X1 U92 ( .A(n1827), .B(\mem<32><5> ), .Y(n1375) );
  AND2X1 U93 ( .A(n1827), .B(\mem<32><6> ), .Y(n1388) );
  AND2X1 U129 ( .A(n1827), .B(\mem<32><7> ), .Y(n1401) );
  INVX1 U589 ( .A(rd1), .Y(n1024) );
  INVX1 U640 ( .A(wr), .Y(n1022) );
  INVX1 U659 ( .A(n1324), .Y(n1021) );
  INVX1 U660 ( .A(n1415), .Y(n1020) );
  INVX1 U664 ( .A(n1426), .Y(n1019) );
  INVX1 U666 ( .A(n1437), .Y(n1018) );
  INVX1 U672 ( .A(n1448), .Y(n1017) );
  INVX1 U675 ( .A(n1459), .Y(n1016) );
  INVX1 U679 ( .A(n1470), .Y(n1015) );
  INVX1 U682 ( .A(n1481), .Y(n1014) );
  INVX1 U694 ( .A(rst), .Y(n1013) );
  INVX2 U697 ( .A(n1013), .Y(n1012) );
  AND2X1 U701 ( .A(wr1), .B(n1013), .Y(n1828) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n1817), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U761 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U772 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U789 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U804 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U819 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U834 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U849 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U864 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U875 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U883 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U885 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U887 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U889 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U891 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U893 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n1828), .Y(n189) );
  AND2X1 U896 ( .A(n1828), .B(n1524), .Y(n289) );
  AND2X1 U897 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1339), .Y(n408) );
  BUFX2 U906 ( .A(n1352), .Y(n409) );
  BUFX2 U907 ( .A(n1365), .Y(n421) );
  BUFX2 U908 ( .A(n1378), .Y(n422) );
  BUFX2 U909 ( .A(n1391), .Y(n434) );
  BUFX2 U910 ( .A(n1404), .Y(n435) );
  BUFX2 U911 ( .A(n1494), .Y(n447) );
  BUFX2 U912 ( .A(n1505), .Y(n448) );
  AND2X2 U913 ( .A(rd), .B(n1508), .Y(n460) );
  INVX1 U914 ( .A(n460), .Y(n461) );
  INVX1 U915 ( .A(n1314), .Y(n473) );
  INVX1 U916 ( .A(n1315), .Y(n474) );
  INVX1 U917 ( .A(n1316), .Y(n486) );
  INVX1 U918 ( .A(n1407), .Y(n487) );
  INVX1 U919 ( .A(n1408), .Y(n507) );
  INVX1 U920 ( .A(n1409), .Y(n508) );
  INVX1 U921 ( .A(n1418), .Y(n522) );
  INVX1 U922 ( .A(n1419), .Y(n523) );
  INVX1 U923 ( .A(n1420), .Y(n537) );
  INVX1 U924 ( .A(n1429), .Y(n538) );
  INVX1 U925 ( .A(n1430), .Y(n552) );
  INVX1 U926 ( .A(n1431), .Y(n553) );
  INVX1 U927 ( .A(n1440), .Y(n567) );
  INVX1 U928 ( .A(n1441), .Y(n568) );
  INVX1 U929 ( .A(n1442), .Y(n582) );
  INVX1 U930 ( .A(n1451), .Y(n583) );
  INVX1 U931 ( .A(n1452), .Y(n591) );
  INVX1 U932 ( .A(n1453), .Y(n592) );
  INVX1 U933 ( .A(n1462), .Y(n871) );
  INVX1 U934 ( .A(n1463), .Y(n872) );
  INVX1 U935 ( .A(n1464), .Y(n873) );
  INVX1 U936 ( .A(n1473), .Y(n874) );
  INVX1 U937 ( .A(n1474), .Y(n875) );
  INVX1 U938 ( .A(n1475), .Y(n876) );
  AND2X2 U939 ( .A(n1328), .B(n1327), .Y(n877) );
  INVX1 U940 ( .A(n877), .Y(n878) );
  AND2X2 U941 ( .A(n1341), .B(n1340), .Y(n879) );
  INVX1 U942 ( .A(n879), .Y(n880) );
  AND2X2 U943 ( .A(n1354), .B(n1353), .Y(n881) );
  INVX1 U944 ( .A(n881), .Y(n882) );
  AND2X2 U945 ( .A(n1367), .B(n1366), .Y(n883) );
  INVX1 U946 ( .A(n883), .Y(n884) );
  AND2X2 U947 ( .A(n1380), .B(n1379), .Y(n885) );
  INVX1 U948 ( .A(n885), .Y(n886) );
  AND2X2 U949 ( .A(n1393), .B(n1392), .Y(n887) );
  INVX1 U950 ( .A(n887), .Y(n888) );
  AND2X2 U951 ( .A(n1483), .B(n1482), .Y(n889) );
  INVX1 U952 ( .A(n889), .Y(n890) );
  AND2X2 U953 ( .A(n1496), .B(n1495), .Y(n891) );
  INVX1 U954 ( .A(n891), .Y(n892) );
  INVX1 U955 ( .A(n1321), .Y(n893) );
  INVX1 U956 ( .A(n1322), .Y(n894) );
  INVX1 U957 ( .A(n1323), .Y(n895) );
  INVX1 U958 ( .A(n1412), .Y(n896) );
  INVX1 U959 ( .A(n1413), .Y(n897) );
  INVX1 U960 ( .A(n1414), .Y(n898) );
  INVX1 U961 ( .A(n1423), .Y(n899) );
  INVX1 U962 ( .A(n1424), .Y(n900) );
  INVX1 U963 ( .A(n1425), .Y(n901) );
  INVX1 U964 ( .A(n1434), .Y(n902) );
  INVX1 U965 ( .A(n1435), .Y(n903) );
  INVX1 U966 ( .A(n1436), .Y(n904) );
  INVX1 U967 ( .A(n1445), .Y(n905) );
  INVX1 U968 ( .A(n1446), .Y(n906) );
  INVX1 U969 ( .A(n1447), .Y(n907) );
  INVX1 U970 ( .A(n1456), .Y(n908) );
  INVX1 U971 ( .A(n1457), .Y(n909) );
  INVX1 U972 ( .A(n1458), .Y(n910) );
  INVX1 U973 ( .A(n1467), .Y(n911) );
  INVX1 U974 ( .A(n1468), .Y(n912) );
  INVX1 U975 ( .A(n1469), .Y(n913) );
  INVX1 U976 ( .A(n1478), .Y(n914) );
  INVX1 U977 ( .A(n1479), .Y(n915) );
  INVX1 U978 ( .A(n1480), .Y(n916) );
  AND2X2 U979 ( .A(n1330), .B(n1329), .Y(n917) );
  INVX1 U980 ( .A(n917), .Y(n918) );
  AND2X2 U981 ( .A(n1343), .B(n1342), .Y(n919) );
  INVX1 U982 ( .A(n919), .Y(n920) );
  AND2X2 U983 ( .A(n1356), .B(n1355), .Y(n921) );
  INVX1 U984 ( .A(n921), .Y(n922) );
  AND2X2 U985 ( .A(n1369), .B(n1368), .Y(n923) );
  INVX1 U986 ( .A(n923), .Y(n924) );
  AND2X2 U987 ( .A(n1382), .B(n1381), .Y(n925) );
  INVX1 U988 ( .A(n925), .Y(n926) );
  AND2X2 U989 ( .A(n1395), .B(n1394), .Y(n927) );
  INVX1 U990 ( .A(n927), .Y(n928) );
  AND2X2 U991 ( .A(n1485), .B(n1484), .Y(n929) );
  INVX1 U992 ( .A(n929), .Y(n930) );
  AND2X2 U993 ( .A(n1498), .B(n1497), .Y(n931) );
  INVX1 U994 ( .A(n931), .Y(n932) );
  BUFX2 U995 ( .A(n1337), .Y(n933) );
  BUFX2 U996 ( .A(n1350), .Y(n934) );
  BUFX2 U997 ( .A(n1363), .Y(n935) );
  BUFX2 U998 ( .A(n1376), .Y(n936) );
  BUFX2 U999 ( .A(n1389), .Y(n937) );
  BUFX2 U1000 ( .A(n1402), .Y(n938) );
  BUFX2 U1001 ( .A(n1492), .Y(n939) );
  INVX1 U1002 ( .A(n970), .Y(n940) );
  INVX1 U1003 ( .A(n1499), .Y(n941) );
  INVX1 U1004 ( .A(n1500), .Y(n942) );
  BUFX2 U1005 ( .A(n1552), .Y(n970) );
  BUFX2 U1006 ( .A(n1838), .Y(err) );
  BUFX2 U1007 ( .A(n1335), .Y(n944) );
  BUFX2 U1008 ( .A(n1348), .Y(n945) );
  BUFX2 U1009 ( .A(n1361), .Y(n946) );
  BUFX2 U1010 ( .A(n1374), .Y(n947) );
  BUFX2 U1011 ( .A(n1387), .Y(n948) );
  BUFX2 U1012 ( .A(n1400), .Y(n949) );
  BUFX2 U1013 ( .A(n1490), .Y(n950) );
  INVX1 U1014 ( .A(n971), .Y(n951) );
  INVX1 U1015 ( .A(n1501), .Y(n952) );
  INVX1 U1016 ( .A(n1502), .Y(n953) );
  BUFX2 U1017 ( .A(n1514), .Y(n971) );
  BUFX2 U1018 ( .A(n1523), .Y(n972) );
  BUFX2 U1019 ( .A(n1541), .Y(n974) );
  BUFX2 U1020 ( .A(n1551), .Y(n975) );
  BUFX2 U1021 ( .A(n1561), .Y(n976) );
  BUFX2 U1022 ( .A(n1571), .Y(n977) );
  BUFX2 U1023 ( .A(n1580), .Y(n978) );
  BUFX2 U1024 ( .A(n1590), .Y(n979) );
  BUFX2 U1025 ( .A(n1610), .Y(n982) );
  BUFX2 U1026 ( .A(n1629), .Y(n985) );
  BUFX2 U1027 ( .A(n1650), .Y(n988) );
  BUFX2 U1028 ( .A(n1670), .Y(n991) );
  BUFX2 U1029 ( .A(n1679), .Y(n992) );
  BUFX2 U1030 ( .A(n1689), .Y(n993) );
  BUFX2 U1031 ( .A(n1698), .Y(n994) );
  BUFX2 U1032 ( .A(n1708), .Y(n995) );
  BUFX2 U1033 ( .A(n1717), .Y(n996) );
  BUFX2 U1034 ( .A(n1727), .Y(n997) );
  BUFX2 U1035 ( .A(n1736), .Y(n998) );
  BUFX2 U1036 ( .A(n1746), .Y(n999) );
  BUFX2 U1037 ( .A(n1765), .Y(n1002) );
  BUFX2 U1038 ( .A(n1785), .Y(n1005) );
  BUFX2 U1039 ( .A(n1805), .Y(n1008) );
  BUFX2 U1040 ( .A(n1818), .Y(n973) );
  AND2X1 U1041 ( .A(n1630), .B(n1318), .Y(n1817) );
  BUFX2 U1042 ( .A(n1837), .Y(n1011) );
  BUFX2 U1043 ( .A(n1600), .Y(n954) );
  BUFX2 U1044 ( .A(n1619), .Y(n955) );
  BUFX2 U1045 ( .A(n1640), .Y(n956) );
  BUFX2 U1046 ( .A(n1660), .Y(n957) );
  BUFX2 U1047 ( .A(n1755), .Y(n958) );
  BUFX2 U1048 ( .A(n1775), .Y(n959) );
  BUFX2 U1049 ( .A(n1795), .Y(n960) );
  BUFX2 U1050 ( .A(n1816), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  INVX1 U1053 ( .A(n965), .Y(n964) );
  AND2X1 U1054 ( .A(n1513), .B(n1512), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n951), .B(n1310), .Y(n1524) );
endmodule


module final_memory_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1838, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1046), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1047), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1048), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1049), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1050), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1051), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1052), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1053), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1054), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1055), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1056), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1057), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1058), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1059), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1060), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1061), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1062), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1063), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1064), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1065), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1066), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1067), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1068), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1069), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1070), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1071), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1072), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1073), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1074), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1075), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1076), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1077), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1078), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1079), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1080), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1081), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1082), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1083), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1085), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1086), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1087), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1088), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1089), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1090), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1091), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1092), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1093), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1094), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1095), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1096), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1097), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1098), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1099), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1100), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1101), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1102), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1103), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1104), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1105), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1106), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1107), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1108), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1109), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1110), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1111), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1112), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1113), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1114), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1115), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1116), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1117), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1118), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1119), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1120), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1121), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1122), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1123), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1124), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1125), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1126), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1127), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1128), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1129), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1130), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1131), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1132), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1133), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1134), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1135), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1136), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1137), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1138), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1139), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1140), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1141), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1142), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1143), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1144), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1145), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1146), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1147), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1148), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1149), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1150), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1151), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1152), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1153), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1154), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1155), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1156), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1157), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1166), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1167), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1168), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1169), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1170), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1171), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1172), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1173), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1174), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1175), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1176), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1177), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1178), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1179), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1180), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1181), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1182), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1183), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1184), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1185), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1186), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1187), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1188), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1189), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1190), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1191), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1192), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1193), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1194), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1195), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1196), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1197), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1198), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1199), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1200), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1201), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1202), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1203), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1204), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1205), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1214), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1215), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1216), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1217), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1218), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1219), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1220), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1221), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1222), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1223), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1224), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1225), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1226), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1227), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1228), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1229), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1230), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1231), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1232), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1233), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1234), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1235), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1236), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1238), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1239), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1240), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1241), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1242), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1243), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1244), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1245), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1246), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1247), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1248), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1249), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1250), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1251), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1252), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1253), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1254), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1255), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1256), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1257), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1258), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1259), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1260), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1261), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1262), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1263), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1264), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1265), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1266), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1267), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1268), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1269), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1270), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1271), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1272), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1273), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1274), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1275), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1276), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1277), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1278), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1279), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1280), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1281), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1282), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1283), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1284), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1285), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1286), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1287), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1288), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1289), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1290), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1291), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1292), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1294), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1295), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1296), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1297), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1298), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1299), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1300), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1301), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1302), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1303), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1304), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1305), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1306), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1307), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1308), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1309), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1477), .B(n1476), .Y(n1478) );
  AND2X2 U10 ( .A(n1472), .B(n1471), .Y(n1473) );
  AND2X2 U11 ( .A(n1466), .B(n1465), .Y(n1467) );
  AND2X2 U12 ( .A(n1461), .B(n1460), .Y(n1462) );
  AND2X2 U13 ( .A(n1455), .B(n1454), .Y(n1456) );
  AND2X2 U14 ( .A(n1450), .B(n1449), .Y(n1451) );
  AND2X2 U15 ( .A(n1444), .B(n1443), .Y(n1445) );
  AND2X2 U16 ( .A(n1439), .B(n1438), .Y(n1440) );
  AND2X2 U17 ( .A(n1433), .B(n1432), .Y(n1434) );
  AND2X2 U18 ( .A(n1428), .B(n1427), .Y(n1429) );
  AND2X2 U19 ( .A(n1422), .B(n1421), .Y(n1423) );
  AND2X2 U20 ( .A(n1417), .B(n1416), .Y(n1418) );
  AND2X2 U21 ( .A(n1411), .B(n1410), .Y(n1412) );
  AND2X2 U22 ( .A(n1406), .B(n1405), .Y(n1407) );
  AND2X2 U30 ( .A(n1326), .B(n1026), .Y(n1631) );
  AND2X2 U31 ( .A(n1325), .B(n1026), .Y(n1786) );
  AND2X2 U32 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1651) );
  AND2X2 U33 ( .A(n1325), .B(\addr_1c<0> ), .Y(n1806) );
  AND2X2 U34 ( .A(n1320), .B(n1319), .Y(n1321) );
  AND2X2 U45 ( .A(n1313), .B(n1312), .Y(n1314) );
  NOR3X1 U94 ( .A(n1022), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1023), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1038), .C(n1836), .Y(n1309) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1836) );
  OAI21X1 U98 ( .A(n1011), .B(n1039), .C(n1835), .Y(n1308) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1835) );
  OAI21X1 U100 ( .A(n1011), .B(n1040), .C(n1834), .Y(n1307) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1834) );
  OAI21X1 U102 ( .A(n1011), .B(n1041), .C(n1833), .Y(n1306) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1833) );
  OAI21X1 U104 ( .A(n1011), .B(n1042), .C(n1832), .Y(n1305) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1832) );
  OAI21X1 U106 ( .A(n1011), .B(n1043), .C(n1831), .Y(n1304) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1831) );
  OAI21X1 U108 ( .A(n1011), .B(n1044), .C(n1830), .Y(n1303) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1830) );
  OAI21X1 U110 ( .A(n1011), .B(n1045), .C(n1829), .Y(n1302) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1829) );
  NAND3X1 U112 ( .A(n1828), .B(n1827), .C(n965), .Y(n1837) );
  OAI21X1 U113 ( .A(n6), .B(n1030), .C(n1826), .Y(n1301) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1826) );
  OAI21X1 U115 ( .A(n6), .B(n1031), .C(n1825), .Y(n1300) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1825) );
  OAI21X1 U117 ( .A(n6), .B(n1032), .C(n1824), .Y(n1299) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1824) );
  OAI21X1 U119 ( .A(n6), .B(n1033), .C(n1823), .Y(n1298) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1823) );
  OAI21X1 U121 ( .A(n6), .B(n1034), .C(n1822), .Y(n1297) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1822) );
  OAI21X1 U123 ( .A(n6), .B(n1035), .C(n1821), .Y(n1296) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1821) );
  OAI21X1 U125 ( .A(n6), .B(n1036), .C(n1820), .Y(n1295) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1820) );
  OAI21X1 U127 ( .A(n6), .B(n1037), .C(n1819), .Y(n1294) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1819) );
  OAI21X1 U130 ( .A(n1038), .B(n1010), .C(n1815), .Y(n1293) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1815) );
  OAI21X1 U132 ( .A(n1039), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1814) );
  OAI21X1 U134 ( .A(n1040), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1813) );
  OAI21X1 U136 ( .A(n1041), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1812) );
  OAI21X1 U138 ( .A(n1042), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1811) );
  OAI21X1 U140 ( .A(n1043), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1810) );
  OAI21X1 U142 ( .A(n1044), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1809) );
  OAI21X1 U144 ( .A(n1045), .B(n1009), .C(n1808), .Y(n1286) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1808) );
  NAND3X1 U146 ( .A(n1807), .B(n1828), .C(n1806), .Y(n1816) );
  OAI21X1 U147 ( .A(n1030), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1804) );
  OAI21X1 U149 ( .A(n1031), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1803) );
  OAI21X1 U151 ( .A(n1032), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1802) );
  OAI21X1 U153 ( .A(n1033), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1801) );
  OAI21X1 U155 ( .A(n1034), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1800) );
  OAI21X1 U157 ( .A(n1035), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1799) );
  OAI21X1 U159 ( .A(n1036), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1798) );
  OAI21X1 U161 ( .A(n1037), .B(n1008), .C(n1797), .Y(n1278) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1797) );
  NAND3X1 U163 ( .A(n973), .B(n1828), .C(n1796), .Y(n1805) );
  OAI21X1 U164 ( .A(n1038), .B(n1007), .C(n1794), .Y(n1277) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1794) );
  OAI21X1 U166 ( .A(n1039), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1793) );
  OAI21X1 U168 ( .A(n1040), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1792) );
  OAI21X1 U170 ( .A(n1041), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1791) );
  OAI21X1 U172 ( .A(n1042), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1790) );
  OAI21X1 U174 ( .A(n1043), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1789) );
  OAI21X1 U176 ( .A(n1044), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1788) );
  OAI21X1 U178 ( .A(n1045), .B(n1006), .C(n1787), .Y(n1270) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1787) );
  NAND3X1 U180 ( .A(n1807), .B(n1828), .C(n1786), .Y(n1795) );
  OAI21X1 U181 ( .A(n1030), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1784) );
  OAI21X1 U183 ( .A(n1031), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1783) );
  OAI21X1 U185 ( .A(n1032), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1782) );
  OAI21X1 U187 ( .A(n1033), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1781) );
  OAI21X1 U189 ( .A(n1034), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1780) );
  OAI21X1 U191 ( .A(n1035), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1779) );
  OAI21X1 U193 ( .A(n1036), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1778) );
  OAI21X1 U195 ( .A(n1037), .B(n1005), .C(n1777), .Y(n1262) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1777) );
  NAND3X1 U197 ( .A(n973), .B(n1828), .C(n1776), .Y(n1785) );
  OAI21X1 U198 ( .A(n1038), .B(n1004), .C(n1774), .Y(n1261) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1774) );
  OAI21X1 U200 ( .A(n1039), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1773) );
  OAI21X1 U202 ( .A(n1040), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1772) );
  OAI21X1 U204 ( .A(n1041), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1771) );
  OAI21X1 U206 ( .A(n1042), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1770) );
  OAI21X1 U208 ( .A(n1043), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1769) );
  OAI21X1 U210 ( .A(n1044), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1768) );
  OAI21X1 U212 ( .A(n1045), .B(n1003), .C(n1767), .Y(n1254) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1767) );
  NAND3X1 U214 ( .A(n1806), .B(n1828), .C(n1766), .Y(n1775) );
  OAI21X1 U215 ( .A(n1030), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1764) );
  OAI21X1 U217 ( .A(n1031), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1763) );
  OAI21X1 U219 ( .A(n1032), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1762) );
  OAI21X1 U221 ( .A(n1033), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1761) );
  OAI21X1 U223 ( .A(n1034), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1760) );
  OAI21X1 U225 ( .A(n1035), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1759) );
  OAI21X1 U227 ( .A(n1036), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1758) );
  OAI21X1 U229 ( .A(n1037), .B(n1002), .C(n1757), .Y(n1246) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1757) );
  NAND3X1 U231 ( .A(n973), .B(n1828), .C(n1756), .Y(n1765) );
  OAI21X1 U232 ( .A(n1038), .B(n1001), .C(n1754), .Y(n1245) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1754) );
  OAI21X1 U234 ( .A(n1039), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1753) );
  OAI21X1 U236 ( .A(n1040), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1752) );
  OAI21X1 U238 ( .A(n1041), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1751) );
  OAI21X1 U240 ( .A(n1042), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1750) );
  OAI21X1 U242 ( .A(n1043), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1749) );
  OAI21X1 U244 ( .A(n1044), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1748) );
  OAI21X1 U246 ( .A(n1045), .B(n1000), .C(n1747), .Y(n1238) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1747) );
  NAND3X1 U248 ( .A(n1786), .B(n1828), .C(n1766), .Y(n1755) );
  OAI21X1 U249 ( .A(n1030), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1745) );
  OAI21X1 U251 ( .A(n1031), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1744) );
  OAI21X1 U253 ( .A(n1032), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1743) );
  OAI21X1 U255 ( .A(n1033), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1742) );
  OAI21X1 U257 ( .A(n1034), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1741) );
  OAI21X1 U259 ( .A(n1035), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1740) );
  OAI21X1 U261 ( .A(n1036), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1739) );
  OAI21X1 U263 ( .A(n1037), .B(n999), .C(n1738), .Y(n1230) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1738) );
  NAND3X1 U265 ( .A(n973), .B(n1828), .C(n1737), .Y(n1746) );
  OAI21X1 U266 ( .A(n1038), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1735) );
  OAI21X1 U268 ( .A(n1039), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1734) );
  OAI21X1 U270 ( .A(n1040), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1733) );
  OAI21X1 U272 ( .A(n1041), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1732) );
  OAI21X1 U274 ( .A(n1042), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1731) );
  OAI21X1 U276 ( .A(n1043), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1730) );
  OAI21X1 U278 ( .A(n1044), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1729) );
  OAI21X1 U280 ( .A(n1045), .B(n998), .C(n1728), .Y(n1222) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1728) );
  NAND3X1 U282 ( .A(n1806), .B(n1828), .C(n969), .Y(n1736) );
  OAI21X1 U283 ( .A(n1030), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1726) );
  OAI21X1 U285 ( .A(n1031), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1725) );
  OAI21X1 U287 ( .A(n1032), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1724) );
  OAI21X1 U289 ( .A(n1033), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1723) );
  OAI21X1 U291 ( .A(n1034), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1722) );
  OAI21X1 U293 ( .A(n1035), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1721) );
  OAI21X1 U295 ( .A(n1036), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1720) );
  OAI21X1 U297 ( .A(n1037), .B(n997), .C(n1719), .Y(n1214) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1719) );
  NAND3X1 U299 ( .A(n973), .B(n1828), .C(n1718), .Y(n1727) );
  OAI21X1 U300 ( .A(n1038), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1716) );
  OAI21X1 U302 ( .A(n1039), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1715) );
  OAI21X1 U304 ( .A(n1040), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1714) );
  OAI21X1 U306 ( .A(n1041), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1713) );
  OAI21X1 U308 ( .A(n1042), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1712) );
  OAI21X1 U310 ( .A(n1043), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1711) );
  OAI21X1 U312 ( .A(n1044), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1710) );
  OAI21X1 U314 ( .A(n1045), .B(n996), .C(n1709), .Y(n1206) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1709) );
  NAND3X1 U316 ( .A(n1786), .B(n1828), .C(n969), .Y(n1717) );
  OAI21X1 U317 ( .A(n1030), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1707) );
  OAI21X1 U319 ( .A(n1031), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1706) );
  OAI21X1 U321 ( .A(n1032), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1705) );
  OAI21X1 U323 ( .A(n1033), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1704) );
  OAI21X1 U325 ( .A(n1034), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1703) );
  OAI21X1 U327 ( .A(n1035), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1702) );
  OAI21X1 U329 ( .A(n1036), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1701) );
  OAI21X1 U331 ( .A(n1037), .B(n995), .C(n1700), .Y(n1198) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1700) );
  NAND3X1 U333 ( .A(n973), .B(n1828), .C(n1699), .Y(n1708) );
  OAI21X1 U334 ( .A(n1038), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1697) );
  OAI21X1 U336 ( .A(n1039), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1696) );
  OAI21X1 U338 ( .A(n1040), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1695) );
  OAI21X1 U340 ( .A(n1041), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1694) );
  OAI21X1 U342 ( .A(n1042), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1693) );
  OAI21X1 U344 ( .A(n1043), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1692) );
  OAI21X1 U346 ( .A(n1044), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1691) );
  OAI21X1 U348 ( .A(n1045), .B(n994), .C(n1690), .Y(n1190) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1690) );
  NAND3X1 U350 ( .A(n1806), .B(n1828), .C(n967), .Y(n1698) );
  OAI21X1 U351 ( .A(n1030), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1688) );
  OAI21X1 U353 ( .A(n1031), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1687) );
  OAI21X1 U355 ( .A(n1032), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1686) );
  OAI21X1 U357 ( .A(n1033), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1685) );
  OAI21X1 U359 ( .A(n1034), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1684) );
  OAI21X1 U361 ( .A(n1035), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1683) );
  OAI21X1 U363 ( .A(n1036), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1682) );
  OAI21X1 U365 ( .A(n1037), .B(n993), .C(n1681), .Y(n1182) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1681) );
  NAND3X1 U367 ( .A(n973), .B(n1828), .C(n1680), .Y(n1689) );
  OAI21X1 U368 ( .A(n1038), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1678) );
  OAI21X1 U370 ( .A(n1039), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1677) );
  OAI21X1 U372 ( .A(n1040), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1676) );
  OAI21X1 U374 ( .A(n1041), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1675) );
  OAI21X1 U376 ( .A(n1042), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1674) );
  OAI21X1 U378 ( .A(n1043), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1673) );
  OAI21X1 U380 ( .A(n1044), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1672) );
  OAI21X1 U382 ( .A(n1045), .B(n992), .C(n1671), .Y(n1174) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1671) );
  NAND3X1 U384 ( .A(n1786), .B(n1828), .C(n967), .Y(n1679) );
  OAI21X1 U385 ( .A(n1030), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1669) );
  OAI21X1 U387 ( .A(n1031), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1668) );
  OAI21X1 U389 ( .A(n1032), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1667) );
  OAI21X1 U391 ( .A(n1033), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1666) );
  OAI21X1 U393 ( .A(n1034), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1665) );
  OAI21X1 U395 ( .A(n1035), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1664) );
  OAI21X1 U397 ( .A(n1036), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1663) );
  OAI21X1 U399 ( .A(n1037), .B(n991), .C(n1662), .Y(n1166) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1662) );
  NAND3X1 U401 ( .A(n973), .B(n1828), .C(n1661), .Y(n1670) );
  OAI21X1 U402 ( .A(n1038), .B(n990), .C(n1659), .Y(n1165) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1659) );
  OAI21X1 U404 ( .A(n1039), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1658) );
  OAI21X1 U406 ( .A(n1040), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1657) );
  OAI21X1 U408 ( .A(n1041), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1656) );
  OAI21X1 U410 ( .A(n1042), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1655) );
  OAI21X1 U412 ( .A(n1043), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1654) );
  OAI21X1 U414 ( .A(n1044), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1653) );
  OAI21X1 U416 ( .A(n1045), .B(n989), .C(n1652), .Y(n1158) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1652) );
  NAND3X1 U418 ( .A(n1807), .B(n1828), .C(n1651), .Y(n1660) );
  OAI21X1 U419 ( .A(n1030), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1649) );
  OAI21X1 U421 ( .A(n1031), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1648) );
  OAI21X1 U423 ( .A(n1032), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1647) );
  OAI21X1 U425 ( .A(n1033), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1646) );
  OAI21X1 U427 ( .A(n1034), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1645) );
  OAI21X1 U429 ( .A(n1035), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1644) );
  OAI21X1 U431 ( .A(n1036), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1643) );
  OAI21X1 U433 ( .A(n1037), .B(n988), .C(n1642), .Y(n1150) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1642) );
  NAND3X1 U435 ( .A(n973), .B(n1828), .C(n1641), .Y(n1650) );
  OAI21X1 U436 ( .A(n1038), .B(n987), .C(n1639), .Y(n1149) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1639) );
  OAI21X1 U438 ( .A(n1039), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1638) );
  OAI21X1 U440 ( .A(n1040), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1637) );
  OAI21X1 U442 ( .A(n1041), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1636) );
  OAI21X1 U444 ( .A(n1042), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1635) );
  OAI21X1 U446 ( .A(n1043), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1634) );
  OAI21X1 U448 ( .A(n1044), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1633) );
  OAI21X1 U450 ( .A(n1045), .B(n986), .C(n1632), .Y(n1142) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1632) );
  NAND3X1 U452 ( .A(n1807), .B(n1828), .C(n1631), .Y(n1640) );
  OAI21X1 U453 ( .A(n1030), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1628) );
  OAI21X1 U455 ( .A(n1031), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1627) );
  OAI21X1 U457 ( .A(n1032), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1626) );
  OAI21X1 U459 ( .A(n1033), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1625) );
  OAI21X1 U461 ( .A(n1034), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1624) );
  OAI21X1 U463 ( .A(n1035), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1623) );
  OAI21X1 U465 ( .A(n1036), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1622) );
  OAI21X1 U467 ( .A(n1037), .B(n985), .C(n1621), .Y(n1134) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1621) );
  NAND3X1 U469 ( .A(n973), .B(n1828), .C(n1620), .Y(n1629) );
  OAI21X1 U470 ( .A(n1038), .B(n984), .C(n1618), .Y(n1133) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1618) );
  OAI21X1 U472 ( .A(n1039), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1617) );
  OAI21X1 U474 ( .A(n1040), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1616) );
  OAI21X1 U476 ( .A(n1041), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1615) );
  OAI21X1 U478 ( .A(n1042), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1614) );
  OAI21X1 U480 ( .A(n1043), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1613) );
  OAI21X1 U482 ( .A(n1044), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1612) );
  OAI21X1 U484 ( .A(n1045), .B(n983), .C(n1611), .Y(n1126) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1611) );
  NAND3X1 U486 ( .A(n1766), .B(n1828), .C(n1651), .Y(n1619) );
  OAI21X1 U487 ( .A(n1030), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1609) );
  OAI21X1 U489 ( .A(n1031), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1608) );
  OAI21X1 U491 ( .A(n1032), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1607) );
  OAI21X1 U493 ( .A(n1033), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1606) );
  OAI21X1 U495 ( .A(n1034), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1605) );
  OAI21X1 U497 ( .A(n1035), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1604) );
  OAI21X1 U499 ( .A(n1036), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1603) );
  OAI21X1 U501 ( .A(n1037), .B(n982), .C(n1602), .Y(n1118) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1602) );
  NAND3X1 U503 ( .A(n973), .B(n1828), .C(n1601), .Y(n1610) );
  OAI21X1 U504 ( .A(n1038), .B(n981), .C(n1599), .Y(n1117) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1599) );
  OAI21X1 U506 ( .A(n1039), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1598) );
  OAI21X1 U508 ( .A(n1040), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1597) );
  OAI21X1 U510 ( .A(n1041), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1596) );
  OAI21X1 U512 ( .A(n1042), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1595) );
  OAI21X1 U514 ( .A(n1043), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1594) );
  OAI21X1 U516 ( .A(n1044), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1593) );
  OAI21X1 U518 ( .A(n1045), .B(n980), .C(n1592), .Y(n1110) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1592) );
  NAND3X1 U520 ( .A(n1766), .B(n1828), .C(n1631), .Y(n1600) );
  OAI21X1 U521 ( .A(n1030), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1589) );
  OAI21X1 U523 ( .A(n1031), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1588) );
  OAI21X1 U525 ( .A(n1032), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1587) );
  OAI21X1 U527 ( .A(n1033), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1586) );
  OAI21X1 U529 ( .A(n1034), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1585) );
  OAI21X1 U531 ( .A(n1035), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1584) );
  OAI21X1 U533 ( .A(n1036), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1583) );
  OAI21X1 U535 ( .A(n1037), .B(n979), .C(n1582), .Y(n1102) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1582) );
  NAND3X1 U537 ( .A(n973), .B(n1828), .C(n1581), .Y(n1590) );
  OAI21X1 U538 ( .A(n1038), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1579) );
  OAI21X1 U540 ( .A(n1039), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1578) );
  OAI21X1 U542 ( .A(n1040), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1577) );
  OAI21X1 U544 ( .A(n1041), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1576) );
  OAI21X1 U546 ( .A(n1042), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1575) );
  OAI21X1 U548 ( .A(n1043), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1574) );
  OAI21X1 U550 ( .A(n1044), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1573) );
  OAI21X1 U552 ( .A(n1045), .B(n978), .C(n1572), .Y(n1094) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1572) );
  NAND3X1 U554 ( .A(n969), .B(n1828), .C(n1651), .Y(n1580) );
  OAI21X1 U555 ( .A(n1030), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1570) );
  OAI21X1 U557 ( .A(n1031), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1569) );
  OAI21X1 U559 ( .A(n1032), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1568) );
  OAI21X1 U561 ( .A(n1033), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1567) );
  OAI21X1 U563 ( .A(n1034), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1566) );
  OAI21X1 U565 ( .A(n1035), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1565) );
  OAI21X1 U567 ( .A(n1036), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1564) );
  OAI21X1 U569 ( .A(n1037), .B(n977), .C(n1563), .Y(n1086) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1563) );
  NAND3X1 U571 ( .A(n973), .B(n1828), .C(n1562), .Y(n1571) );
  OAI21X1 U572 ( .A(n1038), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1560) );
  OAI21X1 U574 ( .A(n1039), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1559) );
  OAI21X1 U576 ( .A(n1040), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1558) );
  OAI21X1 U578 ( .A(n1041), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1557) );
  OAI21X1 U580 ( .A(n1042), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1556) );
  OAI21X1 U582 ( .A(n1043), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1555) );
  OAI21X1 U584 ( .A(n1044), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1554) );
  OAI21X1 U586 ( .A(n1045), .B(n976), .C(n1553), .Y(n1078) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1553) );
  NAND3X1 U588 ( .A(n969), .B(n1828), .C(n1631), .Y(n1561) );
  OAI21X1 U590 ( .A(n1030), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1550) );
  OAI21X1 U592 ( .A(n1031), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1549) );
  OAI21X1 U594 ( .A(n1032), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1548) );
  OAI21X1 U596 ( .A(n1033), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1547) );
  OAI21X1 U598 ( .A(n1034), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1546) );
  OAI21X1 U600 ( .A(n1035), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1545) );
  OAI21X1 U602 ( .A(n1036), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1544) );
  OAI21X1 U604 ( .A(n1037), .B(n975), .C(n1543), .Y(n1070) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1543) );
  NAND3X1 U606 ( .A(n973), .B(n1828), .C(n1542), .Y(n1551) );
  OAI21X1 U607 ( .A(n1038), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1540) );
  OAI21X1 U609 ( .A(n1039), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1539) );
  OAI21X1 U611 ( .A(n1040), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1538) );
  OAI21X1 U613 ( .A(n1041), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1537) );
  OAI21X1 U615 ( .A(n1042), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1536) );
  OAI21X1 U617 ( .A(n1043), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1535) );
  OAI21X1 U619 ( .A(n1044), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1534) );
  OAI21X1 U621 ( .A(n1045), .B(n974), .C(n1533), .Y(n1062) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1533) );
  NAND3X1 U623 ( .A(n967), .B(n1828), .C(n1651), .Y(n1541) );
  OAI21X1 U624 ( .A(n1030), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1532) );
  OAI21X1 U626 ( .A(n1031), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1531) );
  OAI21X1 U628 ( .A(n1032), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1530) );
  OAI21X1 U630 ( .A(n1033), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1529) );
  OAI21X1 U632 ( .A(n1034), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1528) );
  OAI21X1 U634 ( .A(n1035), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1527) );
  OAI21X1 U636 ( .A(n1036), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1526) );
  OAI21X1 U638 ( .A(n1037), .B(n8), .C(n1525), .Y(n1054) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1525) );
  NOR2X1 U641 ( .A(n964), .B(\addr_1c<4> ), .Y(n1818) );
  OAI21X1 U642 ( .A(n1038), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1522) );
  OAI21X1 U644 ( .A(n1039), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1521) );
  OAI21X1 U646 ( .A(n1040), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1520) );
  OAI21X1 U648 ( .A(n1041), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1519) );
  OAI21X1 U650 ( .A(n1042), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1518) );
  OAI21X1 U652 ( .A(n1043), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1517) );
  OAI21X1 U654 ( .A(n1044), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1516) );
  OAI21X1 U656 ( .A(n1045), .B(n972), .C(n1515), .Y(n1046) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1515) );
  NAND3X1 U658 ( .A(n967), .B(n1828), .C(n1631), .Y(n1523) );
  NOR3X1 U661 ( .A(n1511), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1512) );
  NOR3X1 U662 ( .A(n1510), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1513) );
  AOI21X1 U663 ( .A(n461), .B(n1509), .C(n963), .Y(n1838) );
  OAI21X1 U665 ( .A(rd), .B(n1508), .C(wr), .Y(n1509) );
  NAND3X1 U667 ( .A(n1507), .B(n1025), .C(n1506), .Y(n1508) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1506) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1507) );
  AOI21X1 U670 ( .A(n448), .B(n1504), .C(n1024), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1503), .C(n4), .Y(n1504) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1786), .C(\mem<0><1> ), .D(n1631), .Y(
        n1501) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1806), .C(\mem<2><1> ), .D(n1651), .Y(
        n1502) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1786), .C(\mem<4><1> ), .D(n1631), .Y(
        n1499) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1806), .C(\mem<6><1> ), .D(n1651), .Y(
        n1500) );
  AOI22X1 U678 ( .A(n1591), .B(n892), .C(n1630), .D(n932), .Y(n1505) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1786), .C(\mem<12><1> ), .D(n1631), .Y(
        n1497) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1806), .C(\mem<14><1> ), .D(n1651), .Y(
        n1498) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1786), .C(\mem<8><1> ), .D(n1631), .Y(
        n1495) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1806), .C(\mem<10><1> ), .D(n1651), .Y(
        n1496) );
  AOI21X1 U685 ( .A(n447), .B(n1493), .C(n1024), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1491), .C(n949), .Y(n1493) );
  AOI21X1 U687 ( .A(n1489), .B(n1488), .C(n971), .Y(n1490) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1786), .C(\mem<0><0> ), .D(n1631), .Y(
        n1488) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1806), .C(\mem<2><0> ), .D(n1651), .Y(
        n1489) );
  AOI21X1 U690 ( .A(n1487), .B(n1486), .C(n970), .Y(n1492) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1786), .C(\mem<4><0> ), .D(n1631), .Y(
        n1486) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1806), .C(\mem<6><0> ), .D(n1651), .Y(
        n1487) );
  AOI22X1 U693 ( .A(n1591), .B(n890), .C(n1630), .D(n930), .Y(n1494) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1786), .C(\mem<12><0> ), .D(n1631), .Y(
        n1484) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1806), .C(\mem<14><0> ), .D(n1651), .Y(
        n1485) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1786), .C(\mem<8><0> ), .D(n1631), .Y(
        n1482) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1806), .C(\mem<10><0> ), .D(n1651), .Y(
        n1483) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1481) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1680), .C(\mem<19><7> ), .D(n1699), .Y(
        n1476) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1718), .C(\mem<23><7> ), .D(n1737), .Y(
        n1477) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1756), .C(\mem<27><7> ), .D(n1776), .Y(
        n1479) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1796), .C(\mem<31><7> ), .D(n1817), .Y(
        n1480) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1524), .C(\mem<3><7> ), .D(n1542), .Y(
        n1471) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1562), .C(\mem<7><7> ), .D(n1581), .Y(
        n1472) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1601), .C(\mem<11><7> ), .D(n1620), .Y(
        n1474) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1641), .C(\mem<15><7> ), .D(n1661), .Y(
        n1475) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1470) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1680), .C(\mem<19><6> ), .D(n1699), .Y(
        n1465) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1718), .C(\mem<23><6> ), .D(n1737), .Y(
        n1466) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1756), .C(\mem<27><6> ), .D(n1776), .Y(
        n1468) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1796), .C(\mem<31><6> ), .D(n1817), .Y(
        n1469) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1524), .C(\mem<3><6> ), .D(n1542), .Y(
        n1460) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1562), .C(\mem<7><6> ), .D(n1581), .Y(
        n1461) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1601), .C(\mem<11><6> ), .D(n1620), .Y(
        n1463) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1641), .C(\mem<15><6> ), .D(n1661), .Y(
        n1464) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1459) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1680), .C(\mem<19><5> ), .D(n1699), .Y(
        n1454) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1718), .C(\mem<23><5> ), .D(n1737), .Y(
        n1455) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1756), .C(\mem<27><5> ), .D(n1776), .Y(
        n1457) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1796), .C(\mem<31><5> ), .D(n1817), .Y(
        n1458) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1524), .C(\mem<3><5> ), .D(n1542), .Y(
        n1449) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1562), .C(\mem<7><5> ), .D(n1581), .Y(
        n1450) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1601), .C(\mem<11><5> ), .D(n1620), .Y(
        n1452) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1641), .C(\mem<15><5> ), .D(n1661), .Y(
        n1453) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1448) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1680), .C(\mem<19><4> ), .D(n1699), .Y(
        n1443) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1718), .C(\mem<23><4> ), .D(n1737), .Y(
        n1444) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1756), .C(\mem<27><4> ), .D(n1776), .Y(
        n1446) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1796), .C(\mem<31><4> ), .D(n1817), .Y(
        n1447) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1524), .C(\mem<3><4> ), .D(n1542), .Y(
        n1438) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1562), .C(\mem<7><4> ), .D(n1581), .Y(
        n1439) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1601), .C(\mem<11><4> ), .D(n1620), .Y(
        n1441) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1641), .C(\mem<15><4> ), .D(n1661), .Y(
        n1442) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1437) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1680), .C(\mem<19><3> ), .D(n1699), .Y(
        n1432) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1718), .C(\mem<23><3> ), .D(n1737), .Y(
        n1433) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1756), .C(\mem<27><3> ), .D(n1776), .Y(
        n1435) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1796), .C(\mem<31><3> ), .D(n1817), .Y(
        n1436) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1524), .C(\mem<3><3> ), .D(n1542), .Y(
        n1427) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1562), .C(\mem<7><3> ), .D(n1581), .Y(
        n1428) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1601), .C(\mem<11><3> ), .D(n1620), .Y(
        n1430) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1641), .C(\mem<15><3> ), .D(n1661), .Y(
        n1431) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1426) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1680), .C(\mem<19><2> ), .D(n1699), .Y(
        n1421) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1718), .C(\mem<23><2> ), .D(n1737), .Y(
        n1422) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1756), .C(\mem<27><2> ), .D(n1776), .Y(
        n1424) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1796), .C(\mem<31><2> ), .D(n1817), .Y(
        n1425) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1524), .C(\mem<3><2> ), .D(n1542), .Y(
        n1416) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1562), .C(\mem<7><2> ), .D(n1581), .Y(
        n1417) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1601), .C(\mem<11><2> ), .D(n1620), .Y(
        n1419) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1641), .C(\mem<15><2> ), .D(n1661), .Y(
        n1420) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1415) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1680), .C(\mem<19><1> ), .D(n1699), .Y(
        n1410) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1718), .C(\mem<23><1> ), .D(n1737), .Y(
        n1411) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1756), .C(\mem<27><1> ), .D(n1776), .Y(
        n1413) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1796), .C(\mem<31><1> ), .D(n1817), .Y(
        n1414) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1524), .C(\mem<3><1> ), .D(n1542), .Y(
        n1405) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1562), .C(\mem<7><1> ), .D(n1581), .Y(
        n1406) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1601), .C(\mem<11><1> ), .D(n1620), .Y(
        n1408) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1641), .C(\mem<15><1> ), .D(n1661), .Y(
        n1409) );
  AOI21X1 U777 ( .A(n435), .B(n1403), .C(n1024), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1401), .C(n948), .Y(n1403) );
  AOI21X1 U779 ( .A(n1399), .B(n1398), .C(n971), .Y(n1400) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1786), .C(\mem<0><7> ), .D(n1631), .Y(
        n1398) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1806), .C(\mem<2><7> ), .D(n1651), .Y(
        n1399) );
  AOI21X1 U782 ( .A(n1397), .B(n1396), .C(n970), .Y(n1402) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1786), .C(\mem<4><7> ), .D(n1631), .Y(
        n1396) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1806), .C(\mem<6><7> ), .D(n1651), .Y(
        n1397) );
  AOI22X1 U785 ( .A(n1591), .B(n888), .C(n1630), .D(n928), .Y(n1404) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1786), .C(\mem<12><7> ), .D(n1631), .Y(
        n1394) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1806), .C(\mem<14><7> ), .D(n1651), .Y(
        n1395) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1786), .C(\mem<8><7> ), .D(n1631), .Y(
        n1392) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1806), .C(\mem<10><7> ), .D(n1651), .Y(
        n1393) );
  AOI21X1 U792 ( .A(n434), .B(n1390), .C(n1024), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1388), .C(n947), .Y(n1390) );
  AOI21X1 U794 ( .A(n1386), .B(n1385), .C(n971), .Y(n1387) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1786), .C(\mem<0><6> ), .D(n1631), .Y(
        n1385) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1806), .C(\mem<2><6> ), .D(n1651), .Y(
        n1386) );
  AOI21X1 U797 ( .A(n1384), .B(n1383), .C(n970), .Y(n1389) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1786), .C(\mem<4><6> ), .D(n1631), .Y(
        n1383) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1806), .C(\mem<6><6> ), .D(n1651), .Y(
        n1384) );
  AOI22X1 U800 ( .A(n1591), .B(n886), .C(n1630), .D(n926), .Y(n1391) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1786), .C(\mem<12><6> ), .D(n1631), .Y(
        n1381) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1806), .C(\mem<14><6> ), .D(n1651), .Y(
        n1382) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1786), .C(\mem<8><6> ), .D(n1631), .Y(
        n1379) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1806), .C(\mem<10><6> ), .D(n1651), .Y(
        n1380) );
  AOI21X1 U807 ( .A(n422), .B(n1377), .C(n1024), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1375), .C(n946), .Y(n1377) );
  AOI21X1 U809 ( .A(n1373), .B(n1372), .C(n971), .Y(n1374) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1786), .C(\mem<0><5> ), .D(n1631), .Y(
        n1372) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1806), .C(\mem<2><5> ), .D(n1651), .Y(
        n1373) );
  AOI21X1 U812 ( .A(n1371), .B(n1370), .C(n970), .Y(n1376) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1786), .C(\mem<4><5> ), .D(n1631), .Y(
        n1370) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1806), .C(\mem<6><5> ), .D(n1651), .Y(
        n1371) );
  AOI22X1 U815 ( .A(n1591), .B(n884), .C(n1630), .D(n924), .Y(n1378) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1786), .C(\mem<12><5> ), .D(n1631), .Y(
        n1368) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1806), .C(\mem<14><5> ), .D(n1651), .Y(
        n1369) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1786), .C(\mem<8><5> ), .D(n1631), .Y(
        n1366) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1806), .C(\mem<10><5> ), .D(n1651), .Y(
        n1367) );
  AOI21X1 U822 ( .A(n421), .B(n1364), .C(n1024), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1362), .C(n945), .Y(n1364) );
  AOI21X1 U824 ( .A(n1360), .B(n1359), .C(n971), .Y(n1361) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1786), .C(\mem<0><4> ), .D(n1631), .Y(
        n1359) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1806), .C(\mem<2><4> ), .D(n1651), .Y(
        n1360) );
  AOI21X1 U827 ( .A(n1358), .B(n1357), .C(n970), .Y(n1363) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1786), .C(\mem<4><4> ), .D(n1631), .Y(
        n1357) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1806), .C(\mem<6><4> ), .D(n1651), .Y(
        n1358) );
  AOI22X1 U830 ( .A(n1591), .B(n882), .C(n1630), .D(n922), .Y(n1365) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1786), .C(\mem<12><4> ), .D(n1631), .Y(
        n1355) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1806), .C(\mem<14><4> ), .D(n1651), .Y(
        n1356) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1786), .C(\mem<8><4> ), .D(n1631), .Y(
        n1353) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1806), .C(\mem<10><4> ), .D(n1651), .Y(
        n1354) );
  AOI21X1 U837 ( .A(n409), .B(n1351), .C(n1024), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1349), .C(n944), .Y(n1351) );
  AOI21X1 U839 ( .A(n1347), .B(n1346), .C(n971), .Y(n1348) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1786), .C(\mem<0><3> ), .D(n1631), .Y(
        n1346) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1806), .C(\mem<2><3> ), .D(n1651), .Y(
        n1347) );
  AOI21X1 U842 ( .A(n1345), .B(n1344), .C(n970), .Y(n1350) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1786), .C(\mem<4><3> ), .D(n1631), .Y(
        n1344) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1806), .C(\mem<6><3> ), .D(n1651), .Y(
        n1345) );
  AOI22X1 U845 ( .A(n1591), .B(n880), .C(n1630), .D(n920), .Y(n1352) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1786), .C(\mem<12><3> ), .D(n1631), .Y(
        n1342) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1806), .C(\mem<14><3> ), .D(n1651), .Y(
        n1343) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1786), .C(\mem<8><3> ), .D(n1631), .Y(
        n1340) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1806), .C(\mem<10><3> ), .D(n1651), .Y(
        n1341) );
  AOI21X1 U852 ( .A(n408), .B(n1338), .C(n1024), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1336), .C(n943), .Y(n1338) );
  AOI21X1 U854 ( .A(n1334), .B(n1333), .C(n971), .Y(n1335) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1786), .C(\mem<0><2> ), .D(n1631), .Y(
        n1333) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1806), .C(\mem<2><2> ), .D(n1651), .Y(
        n1334) );
  AOI21X1 U857 ( .A(n1332), .B(n1331), .C(n970), .Y(n1337) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1786), .C(\mem<4><2> ), .D(n1631), .Y(
        n1331) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1806), .C(\mem<6><2> ), .D(n1651), .Y(
        n1332) );
  AOI22X1 U860 ( .A(n1591), .B(n878), .C(n1630), .D(n918), .Y(n1339) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1786), .C(\mem<12><2> ), .D(n1631), .Y(
        n1329) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1806), .C(\mem<14><2> ), .D(n1651), .Y(
        n1330) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1786), .C(\mem<8><2> ), .D(n1631), .Y(
        n1327) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1806), .C(\mem<10><2> ), .D(n1651), .Y(
        n1328) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1326) );
  NOR2X1 U868 ( .A(n1029), .B(\addr_1c<4> ), .Y(n1325) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1324) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1680), .C(\mem<19><0> ), .D(n1699), .Y(
        n1319) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1718), .C(\mem<23><0> ), .D(n1737), .Y(
        n1320) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1756), .C(\mem<27><0> ), .D(n1776), .Y(
        n1322) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1796), .C(\mem<31><0> ), .D(n1817), .Y(
        n1323) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1524), .C(\mem<3><0> ), .D(n1542), .Y(
        n1312) );
  NAND2X1 U877 ( .A(n1027), .B(n1028), .Y(n1514) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1562), .C(\mem<7><0> ), .D(n1581), .Y(
        n1313) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1028), .Y(n1552) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1601), .C(\mem<11><0> ), .D(n1620), .Y(
        n1315) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1641), .C(\mem<15><0> ), .D(n1661), .Y(
        n1316) );
  dff_101 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(rst) );
  dff_100 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(rst) );
  dff_99 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(rst) );
  dff_98 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(rst) );
  dff_97 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(rst) );
  dff_96 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(rst) );
  dff_95 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(rst) );
  dff_94 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(rst) );
  dff_93 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(rst) );
  dff_92 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(rst) );
  dff_91 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(rst) );
  dff_90 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(rst) );
  dff_89 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(rst)
         );
  dff_88 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(rst)
         );
  dff_87 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(rst)
         );
  dff_86 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_85 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_84 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_83 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_82 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_81 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_80 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_79 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_78 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_77 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_76 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_75 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_74 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_73 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_72 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_71 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_70 \reg2[0]  ( .q(\data_out<0> ), .d(n1021), .clk(clk), .rst(rst) );
  dff_69 \reg2[1]  ( .q(\data_out<1> ), .d(n1020), .clk(clk), .rst(rst) );
  dff_68 \reg2[2]  ( .q(\data_out<2> ), .d(n1019), .clk(clk), .rst(rst) );
  dff_67 \reg2[3]  ( .q(\data_out<3> ), .d(n1018), .clk(clk), .rst(rst) );
  dff_66 \reg2[4]  ( .q(\data_out<4> ), .d(n1017), .clk(clk), .rst(rst) );
  dff_65 \reg2[5]  ( .q(\data_out<5> ), .d(n1016), .clk(clk), .rst(rst) );
  dff_64 \reg2[6]  ( .q(\data_out<6> ), .d(n1015), .clk(clk), .rst(rst) );
  dff_63 \reg2[7]  ( .q(\data_out<7> ), .d(n1014), .clk(clk), .rst(rst) );
  dff_62 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        rst) );
  dff_61 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        rst) );
  dff_60 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(rst) );
  dff_59 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(rst) );
  dff_58 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(rst) );
  dff_57 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(rst) );
  dff_56 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(rst) );
  dff_55 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(rst) );
  dff_54 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(rst) );
  dff_53 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(rst) );
  dff_52 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(rst) );
  dff_51 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(rst) );
  INVX1 U2 ( .A(rd), .Y(n1023) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1510) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n1524), .Y(n1827) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1029) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1028) );
  OR2X1 U7 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1511) );
  AND2X1 U8 ( .A(n1630), .B(n965), .Y(n1807) );
  AND2X1 U23 ( .A(n1591), .B(n965), .Y(n1766) );
  INVX1 U24 ( .A(\addr_1c<0> ), .Y(n1026) );
  AND2X1 U25 ( .A(n1026), .B(n1029), .Y(n1310) );
  AND2X1 U26 ( .A(\addr_1c<0> ), .B(n1029), .Y(n1311) );
  AND2X1 U27 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1318) );
  AND2X1 U28 ( .A(\addr_1c<3> ), .B(n1026), .Y(n1317) );
  INVX1 U29 ( .A(\addr_1c<1> ), .Y(n1027) );
  INVX1 U35 ( .A(wr1), .Y(n1025) );
  AND2X1 U36 ( .A(n1591), .B(n1318), .Y(n1776) );
  AND2X1 U37 ( .A(n1591), .B(n1317), .Y(n1756) );
  AND2X1 U38 ( .A(n940), .B(n1318), .Y(n1737) );
  AND2X1 U39 ( .A(n940), .B(n1317), .Y(n1718) );
  AND2X1 U40 ( .A(n1318), .B(n950), .Y(n1699) );
  AND2X1 U41 ( .A(n1317), .B(n950), .Y(n1680) );
  AND2X1 U42 ( .A(n1311), .B(n1591), .Y(n1620) );
  AND2X1 U43 ( .A(n1591), .B(n1310), .Y(n1601) );
  AND2X1 U44 ( .A(n1311), .B(n940), .Y(n1581) );
  AND2X1 U46 ( .A(n940), .B(n1310), .Y(n1562) );
  OR2X1 U47 ( .A(n970), .B(n964), .Y(n968) );
  AND2X1 U48 ( .A(n1311), .B(n950), .Y(n1542) );
  OR2X1 U49 ( .A(n964), .B(n971), .Y(n966) );
  AND2X1 U50 ( .A(n1630), .B(n1310), .Y(n1641) );
  AND2X1 U51 ( .A(n1311), .B(n1630), .Y(n1661) );
  AND2X1 U52 ( .A(n1317), .B(n1630), .Y(n1796) );
  AND2X1 U53 ( .A(\addr_1c<2> ), .B(n1027), .Y(n1591) );
  AND2X1 U54 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1630) );
  BUFX2 U55 ( .A(n961), .Y(n1010) );
  BUFX2 U56 ( .A(n961), .Y(n1009) );
  BUFX2 U57 ( .A(n960), .Y(n1007) );
  BUFX2 U58 ( .A(n960), .Y(n1006) );
  BUFX2 U59 ( .A(n959), .Y(n1004) );
  BUFX2 U60 ( .A(n959), .Y(n1003) );
  BUFX2 U61 ( .A(n958), .Y(n1001) );
  BUFX2 U62 ( .A(n958), .Y(n1000) );
  BUFX2 U63 ( .A(n957), .Y(n990) );
  BUFX2 U64 ( .A(n957), .Y(n989) );
  BUFX2 U65 ( .A(n956), .Y(n987) );
  BUFX2 U66 ( .A(n956), .Y(n986) );
  BUFX2 U67 ( .A(n955), .Y(n984) );
  BUFX2 U68 ( .A(n955), .Y(n983) );
  BUFX2 U69 ( .A(n954), .Y(n981) );
  BUFX2 U70 ( .A(n954), .Y(n980) );
  INVX1 U71 ( .A(\data_in_1c<0> ), .Y(n1030) );
  INVX1 U72 ( .A(\data_in_1c<1> ), .Y(n1031) );
  INVX1 U73 ( .A(\data_in_1c<2> ), .Y(n1032) );
  INVX1 U74 ( .A(\data_in_1c<3> ), .Y(n1033) );
  INVX1 U75 ( .A(\data_in_1c<4> ), .Y(n1034) );
  INVX1 U76 ( .A(\data_in_1c<5> ), .Y(n1035) );
  INVX1 U77 ( .A(\data_in_1c<6> ), .Y(n1036) );
  INVX1 U78 ( .A(\data_in_1c<7> ), .Y(n1037) );
  INVX1 U79 ( .A(\data_in_1c<8> ), .Y(n1038) );
  INVX1 U80 ( .A(\data_in_1c<9> ), .Y(n1039) );
  INVX1 U81 ( .A(\data_in_1c<10> ), .Y(n1040) );
  INVX1 U82 ( .A(\data_in_1c<11> ), .Y(n1041) );
  INVX1 U83 ( .A(\data_in_1c<12> ), .Y(n1042) );
  INVX1 U84 ( .A(\data_in_1c<13> ), .Y(n1043) );
  INVX1 U85 ( .A(\data_in_1c<14> ), .Y(n1044) );
  INVX1 U86 ( .A(\data_in_1c<15> ), .Y(n1045) );
  AND2X1 U87 ( .A(n1827), .B(\mem<32><0> ), .Y(n1491) );
  AND2X1 U88 ( .A(n1827), .B(\mem<32><1> ), .Y(n1503) );
  AND2X1 U89 ( .A(n1827), .B(\mem<32><2> ), .Y(n1336) );
  AND2X1 U90 ( .A(n1827), .B(\mem<32><3> ), .Y(n1349) );
  AND2X1 U91 ( .A(n1827), .B(\mem<32><4> ), .Y(n1362) );
  AND2X1 U92 ( .A(n1827), .B(\mem<32><5> ), .Y(n1375) );
  AND2X1 U93 ( .A(n1827), .B(\mem<32><6> ), .Y(n1388) );
  AND2X1 U129 ( .A(n1827), .B(\mem<32><7> ), .Y(n1401) );
  INVX1 U589 ( .A(rd1), .Y(n1024) );
  INVX1 U640 ( .A(wr), .Y(n1022) );
  INVX1 U659 ( .A(n1324), .Y(n1021) );
  INVX1 U660 ( .A(n1415), .Y(n1020) );
  INVX1 U664 ( .A(n1426), .Y(n1019) );
  INVX1 U666 ( .A(n1437), .Y(n1018) );
  INVX1 U672 ( .A(n1448), .Y(n1017) );
  INVX1 U675 ( .A(n1459), .Y(n1016) );
  INVX1 U679 ( .A(n1470), .Y(n1015) );
  INVX1 U682 ( .A(n1481), .Y(n1014) );
  INVX1 U694 ( .A(rst), .Y(n1013) );
  INVX1 U697 ( .A(n1013), .Y(n1012) );
  AND2X1 U701 ( .A(wr1), .B(n1013), .Y(n1828) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n1817), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U761 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U772 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U789 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U804 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U819 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U834 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U849 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U864 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U875 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U883 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U885 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U887 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U889 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U891 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U893 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n1828), .Y(n189) );
  AND2X1 U896 ( .A(n1828), .B(n1524), .Y(n289) );
  AND2X1 U897 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n950), .B(n952), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n950), .B(n951), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1339), .Y(n408) );
  BUFX2 U906 ( .A(n1352), .Y(n409) );
  BUFX2 U907 ( .A(n1365), .Y(n421) );
  BUFX2 U908 ( .A(n1378), .Y(n422) );
  BUFX2 U909 ( .A(n1391), .Y(n434) );
  BUFX2 U910 ( .A(n1404), .Y(n435) );
  BUFX2 U911 ( .A(n1494), .Y(n447) );
  BUFX2 U912 ( .A(n1505), .Y(n448) );
  AND2X2 U913 ( .A(rd), .B(n1508), .Y(n460) );
  INVX1 U914 ( .A(n460), .Y(n461) );
  INVX1 U915 ( .A(n1314), .Y(n473) );
  INVX1 U916 ( .A(n1315), .Y(n474) );
  INVX1 U917 ( .A(n1316), .Y(n486) );
  INVX1 U918 ( .A(n1407), .Y(n487) );
  INVX1 U919 ( .A(n1408), .Y(n507) );
  INVX1 U920 ( .A(n1409), .Y(n508) );
  INVX1 U921 ( .A(n1418), .Y(n522) );
  INVX1 U922 ( .A(n1419), .Y(n523) );
  INVX1 U923 ( .A(n1420), .Y(n537) );
  INVX1 U924 ( .A(n1429), .Y(n538) );
  INVX1 U925 ( .A(n1430), .Y(n552) );
  INVX1 U926 ( .A(n1431), .Y(n553) );
  INVX1 U927 ( .A(n1440), .Y(n567) );
  INVX1 U928 ( .A(n1441), .Y(n568) );
  INVX1 U929 ( .A(n1442), .Y(n582) );
  INVX1 U930 ( .A(n1451), .Y(n583) );
  INVX1 U931 ( .A(n1452), .Y(n591) );
  INVX1 U932 ( .A(n1453), .Y(n592) );
  INVX1 U933 ( .A(n1462), .Y(n871) );
  INVX1 U934 ( .A(n1463), .Y(n872) );
  INVX1 U935 ( .A(n1464), .Y(n873) );
  INVX1 U936 ( .A(n1473), .Y(n874) );
  INVX1 U937 ( .A(n1474), .Y(n875) );
  INVX1 U938 ( .A(n1475), .Y(n876) );
  AND2X2 U939 ( .A(n1328), .B(n1327), .Y(n877) );
  INVX1 U940 ( .A(n877), .Y(n878) );
  AND2X2 U941 ( .A(n1341), .B(n1340), .Y(n879) );
  INVX1 U942 ( .A(n879), .Y(n880) );
  AND2X2 U943 ( .A(n1354), .B(n1353), .Y(n881) );
  INVX1 U944 ( .A(n881), .Y(n882) );
  AND2X2 U945 ( .A(n1367), .B(n1366), .Y(n883) );
  INVX1 U946 ( .A(n883), .Y(n884) );
  AND2X2 U947 ( .A(n1380), .B(n1379), .Y(n885) );
  INVX1 U948 ( .A(n885), .Y(n886) );
  AND2X2 U949 ( .A(n1393), .B(n1392), .Y(n887) );
  INVX1 U950 ( .A(n887), .Y(n888) );
  AND2X2 U951 ( .A(n1483), .B(n1482), .Y(n889) );
  INVX1 U952 ( .A(n889), .Y(n890) );
  AND2X2 U953 ( .A(n1496), .B(n1495), .Y(n891) );
  INVX1 U954 ( .A(n891), .Y(n892) );
  INVX1 U955 ( .A(n1321), .Y(n893) );
  INVX1 U956 ( .A(n1322), .Y(n894) );
  INVX1 U957 ( .A(n1323), .Y(n895) );
  INVX1 U958 ( .A(n1412), .Y(n896) );
  INVX1 U959 ( .A(n1413), .Y(n897) );
  INVX1 U960 ( .A(n1414), .Y(n898) );
  INVX1 U961 ( .A(n1423), .Y(n899) );
  INVX1 U962 ( .A(n1424), .Y(n900) );
  INVX1 U963 ( .A(n1425), .Y(n901) );
  INVX1 U964 ( .A(n1434), .Y(n902) );
  INVX1 U965 ( .A(n1435), .Y(n903) );
  INVX1 U966 ( .A(n1436), .Y(n904) );
  INVX1 U967 ( .A(n1445), .Y(n905) );
  INVX1 U968 ( .A(n1446), .Y(n906) );
  INVX1 U969 ( .A(n1447), .Y(n907) );
  INVX1 U970 ( .A(n1456), .Y(n908) );
  INVX1 U971 ( .A(n1457), .Y(n909) );
  INVX1 U972 ( .A(n1458), .Y(n910) );
  INVX1 U973 ( .A(n1467), .Y(n911) );
  INVX1 U974 ( .A(n1468), .Y(n912) );
  INVX1 U975 ( .A(n1469), .Y(n913) );
  INVX1 U976 ( .A(n1478), .Y(n914) );
  INVX1 U977 ( .A(n1479), .Y(n915) );
  INVX1 U978 ( .A(n1480), .Y(n916) );
  AND2X2 U979 ( .A(n1330), .B(n1329), .Y(n917) );
  INVX1 U980 ( .A(n917), .Y(n918) );
  AND2X2 U981 ( .A(n1343), .B(n1342), .Y(n919) );
  INVX1 U982 ( .A(n919), .Y(n920) );
  AND2X2 U983 ( .A(n1356), .B(n1355), .Y(n921) );
  INVX1 U984 ( .A(n921), .Y(n922) );
  AND2X2 U985 ( .A(n1369), .B(n1368), .Y(n923) );
  INVX1 U986 ( .A(n923), .Y(n924) );
  AND2X2 U987 ( .A(n1382), .B(n1381), .Y(n925) );
  INVX1 U988 ( .A(n925), .Y(n926) );
  AND2X2 U989 ( .A(n1395), .B(n1394), .Y(n927) );
  INVX1 U990 ( .A(n927), .Y(n928) );
  AND2X2 U991 ( .A(n1485), .B(n1484), .Y(n929) );
  INVX1 U992 ( .A(n929), .Y(n930) );
  AND2X2 U993 ( .A(n1498), .B(n1497), .Y(n931) );
  INVX1 U994 ( .A(n931), .Y(n932) );
  BUFX2 U995 ( .A(n1337), .Y(n933) );
  BUFX2 U996 ( .A(n1350), .Y(n934) );
  BUFX2 U997 ( .A(n1363), .Y(n935) );
  BUFX2 U998 ( .A(n1376), .Y(n936) );
  BUFX2 U999 ( .A(n1389), .Y(n937) );
  BUFX2 U1000 ( .A(n1402), .Y(n938) );
  BUFX2 U1001 ( .A(n1492), .Y(n939) );
  INVX1 U1002 ( .A(n970), .Y(n940) );
  INVX1 U1003 ( .A(n1499), .Y(n941) );
  INVX1 U1004 ( .A(n1500), .Y(n942) );
  BUFX2 U1005 ( .A(n1552), .Y(n970) );
  BUFX2 U1006 ( .A(n1335), .Y(n943) );
  BUFX2 U1007 ( .A(n1348), .Y(n944) );
  BUFX2 U1008 ( .A(n1361), .Y(n945) );
  BUFX2 U1009 ( .A(n1374), .Y(n946) );
  BUFX2 U1010 ( .A(n1387), .Y(n947) );
  BUFX2 U1011 ( .A(n1400), .Y(n948) );
  BUFX2 U1012 ( .A(n1490), .Y(n949) );
  INVX1 U1013 ( .A(n971), .Y(n950) );
  INVX1 U1014 ( .A(n1501), .Y(n951) );
  INVX1 U1015 ( .A(n1502), .Y(n952) );
  BUFX2 U1016 ( .A(n1514), .Y(n971) );
  BUFX2 U1017 ( .A(n1838), .Y(err) );
  BUFX2 U1018 ( .A(n1523), .Y(n972) );
  BUFX2 U1019 ( .A(n1541), .Y(n974) );
  BUFX2 U1020 ( .A(n1551), .Y(n975) );
  BUFX2 U1021 ( .A(n1561), .Y(n976) );
  BUFX2 U1022 ( .A(n1571), .Y(n977) );
  BUFX2 U1023 ( .A(n1580), .Y(n978) );
  BUFX2 U1024 ( .A(n1590), .Y(n979) );
  BUFX2 U1025 ( .A(n1610), .Y(n982) );
  BUFX2 U1026 ( .A(n1629), .Y(n985) );
  BUFX2 U1027 ( .A(n1650), .Y(n988) );
  BUFX2 U1028 ( .A(n1670), .Y(n991) );
  BUFX2 U1029 ( .A(n1679), .Y(n992) );
  BUFX2 U1030 ( .A(n1689), .Y(n993) );
  BUFX2 U1031 ( .A(n1698), .Y(n994) );
  BUFX2 U1032 ( .A(n1708), .Y(n995) );
  BUFX2 U1033 ( .A(n1717), .Y(n996) );
  BUFX2 U1034 ( .A(n1727), .Y(n997) );
  BUFX2 U1035 ( .A(n1736), .Y(n998) );
  BUFX2 U1036 ( .A(n1746), .Y(n999) );
  BUFX2 U1037 ( .A(n1765), .Y(n1002) );
  BUFX2 U1038 ( .A(n1785), .Y(n1005) );
  BUFX2 U1039 ( .A(n1805), .Y(n1008) );
  BUFX2 U1040 ( .A(n1818), .Y(n973) );
  AND2X1 U1041 ( .A(n1630), .B(n1318), .Y(n1817) );
  BUFX2 U1042 ( .A(n1837), .Y(n1011) );
  BUFX2 U1043 ( .A(n1600), .Y(n954) );
  BUFX2 U1044 ( .A(n1619), .Y(n955) );
  BUFX2 U1045 ( .A(n1640), .Y(n956) );
  BUFX2 U1046 ( .A(n1660), .Y(n957) );
  BUFX2 U1047 ( .A(n1755), .Y(n958) );
  BUFX2 U1048 ( .A(n1775), .Y(n959) );
  BUFX2 U1049 ( .A(n1795), .Y(n960) );
  BUFX2 U1050 ( .A(n1816), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  INVX1 U1053 ( .A(n965), .Y(n964) );
  AND2X1 U1054 ( .A(n1513), .B(n1512), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n950), .B(n1310), .Y(n1524) );
endmodule


module final_memory_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1838, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1046), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1047), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1048), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1049), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1050), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1051), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1052), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1053), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1054), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1055), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1056), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1057), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1058), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1059), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1060), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1061), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1062), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1063), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1064), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1065), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1066), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1067), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1068), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1069), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1070), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1071), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1072), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1073), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1074), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1075), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1076), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1077), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1078), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1079), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1080), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1081), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1082), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1083), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1085), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1086), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1087), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1088), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1089), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1090), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1091), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1092), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1093), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1094), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1095), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1096), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1097), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1098), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1099), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1100), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1101), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1102), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1103), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1104), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1105), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1106), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1107), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1108), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1109), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1110), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1111), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1112), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1113), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1114), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1115), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1116), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1117), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1118), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1119), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1120), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1121), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1122), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1123), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1124), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1125), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1126), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1127), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1128), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1129), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1130), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1131), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1132), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1133), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1134), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1135), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1136), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1137), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1138), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1139), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1140), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1141), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1142), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1143), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1144), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1145), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1146), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1147), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1148), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1149), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1150), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1151), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1152), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1153), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1154), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1155), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1156), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1157), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1158), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1159), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1160), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1161), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1162), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1163), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1164), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1165), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1166), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1167), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1168), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1169), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1170), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1171), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1172), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1173), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1174), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1175), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1176), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1177), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1178), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1179), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1180), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1181), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1182), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1183), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1184), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1185), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1186), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1187), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1188), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1189), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1190), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1191), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1192), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1193), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1194), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1195), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1196), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1197), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1198), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1199), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1200), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1201), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1202), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1203), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1204), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1205), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1206), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1207), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1208), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1209), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1210), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1211), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1212), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1213), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1214), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1215), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1216), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1217), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1218), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1219), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1220), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1221), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1222), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1223), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1224), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1225), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1226), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1227), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1228), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1229), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1230), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1231), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1232), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1233), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1234), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1235), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1236), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1237), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1238), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1239), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1240), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1241), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1242), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1243), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1244), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1245), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1246), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1247), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1248), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1249), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1250), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1251), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1252), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1253), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1254), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1255), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1256), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1257), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1258), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1259), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1260), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1261), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1262), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1263), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1264), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1265), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1266), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1267), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1268), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1269), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1270), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1271), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1272), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1273), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1274), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1275), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1276), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1277), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1278), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1279), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1280), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1281), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1282), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1283), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1284), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1285), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1286), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1287), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1288), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1289), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1290), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1291), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1292), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1294), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1295), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1296), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1297), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1298), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1299), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1300), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1301), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1302), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1303), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1304), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1305), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1306), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1307), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1308), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1309), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1477), .B(n1476), .Y(n1478) );
  AND2X2 U10 ( .A(n1472), .B(n1471), .Y(n1473) );
  AND2X2 U11 ( .A(n1466), .B(n1465), .Y(n1467) );
  AND2X2 U12 ( .A(n1461), .B(n1460), .Y(n1462) );
  AND2X2 U13 ( .A(n1455), .B(n1454), .Y(n1456) );
  AND2X2 U14 ( .A(n1450), .B(n1449), .Y(n1451) );
  AND2X2 U15 ( .A(n1444), .B(n1443), .Y(n1445) );
  AND2X2 U16 ( .A(n1439), .B(n1438), .Y(n1440) );
  AND2X2 U17 ( .A(n1433), .B(n1432), .Y(n1434) );
  AND2X2 U18 ( .A(n1428), .B(n1427), .Y(n1429) );
  AND2X2 U19 ( .A(n1422), .B(n1421), .Y(n1423) );
  AND2X2 U20 ( .A(n1417), .B(n1416), .Y(n1418) );
  AND2X2 U21 ( .A(n1411), .B(n1410), .Y(n1412) );
  AND2X2 U22 ( .A(n1406), .B(n1405), .Y(n1407) );
  AND2X2 U30 ( .A(n1326), .B(n1026), .Y(n1631) );
  AND2X2 U31 ( .A(n1325), .B(n1026), .Y(n1786) );
  AND2X2 U32 ( .A(n1326), .B(\addr_1c<0> ), .Y(n1651) );
  AND2X2 U33 ( .A(n1325), .B(\addr_1c<0> ), .Y(n1806) );
  AND2X2 U34 ( .A(n1320), .B(n1319), .Y(n1321) );
  AND2X2 U45 ( .A(n1313), .B(n1312), .Y(n1314) );
  NOR3X1 U94 ( .A(n1022), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1023), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1038), .C(n1836), .Y(n1309) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1836) );
  OAI21X1 U98 ( .A(n1011), .B(n1039), .C(n1835), .Y(n1308) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1835) );
  OAI21X1 U100 ( .A(n1011), .B(n1040), .C(n1834), .Y(n1307) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1834) );
  OAI21X1 U102 ( .A(n1011), .B(n1041), .C(n1833), .Y(n1306) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1833) );
  OAI21X1 U104 ( .A(n1011), .B(n1042), .C(n1832), .Y(n1305) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1832) );
  OAI21X1 U106 ( .A(n1011), .B(n1043), .C(n1831), .Y(n1304) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1831) );
  OAI21X1 U108 ( .A(n1011), .B(n1044), .C(n1830), .Y(n1303) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1830) );
  OAI21X1 U110 ( .A(n1011), .B(n1045), .C(n1829), .Y(n1302) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1829) );
  NAND3X1 U112 ( .A(n1828), .B(n1827), .C(n965), .Y(n1837) );
  OAI21X1 U113 ( .A(n6), .B(n1030), .C(n1826), .Y(n1301) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1826) );
  OAI21X1 U115 ( .A(n6), .B(n1031), .C(n1825), .Y(n1300) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1825) );
  OAI21X1 U117 ( .A(n6), .B(n1032), .C(n1824), .Y(n1299) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1824) );
  OAI21X1 U119 ( .A(n6), .B(n1033), .C(n1823), .Y(n1298) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1823) );
  OAI21X1 U121 ( .A(n6), .B(n1034), .C(n1822), .Y(n1297) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1822) );
  OAI21X1 U123 ( .A(n6), .B(n1035), .C(n1821), .Y(n1296) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1821) );
  OAI21X1 U125 ( .A(n6), .B(n1036), .C(n1820), .Y(n1295) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1820) );
  OAI21X1 U127 ( .A(n6), .B(n1037), .C(n1819), .Y(n1294) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1819) );
  OAI21X1 U130 ( .A(n1038), .B(n1010), .C(n1815), .Y(n1293) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1815) );
  OAI21X1 U132 ( .A(n1039), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1814) );
  OAI21X1 U134 ( .A(n1040), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1813) );
  OAI21X1 U136 ( .A(n1041), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1812) );
  OAI21X1 U138 ( .A(n1042), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1811) );
  OAI21X1 U140 ( .A(n1043), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1810) );
  OAI21X1 U142 ( .A(n1044), .B(n1009), .C(n1809), .Y(n1287) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1809) );
  OAI21X1 U144 ( .A(n1045), .B(n1009), .C(n1808), .Y(n1286) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1808) );
  NAND3X1 U146 ( .A(n1807), .B(n1828), .C(n1806), .Y(n1816) );
  OAI21X1 U147 ( .A(n1030), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1804) );
  OAI21X1 U149 ( .A(n1031), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1803) );
  OAI21X1 U151 ( .A(n1032), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1802) );
  OAI21X1 U153 ( .A(n1033), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1801) );
  OAI21X1 U155 ( .A(n1034), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1800) );
  OAI21X1 U157 ( .A(n1035), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1799) );
  OAI21X1 U159 ( .A(n1036), .B(n1008), .C(n1798), .Y(n1279) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1798) );
  OAI21X1 U161 ( .A(n1037), .B(n1008), .C(n1797), .Y(n1278) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1797) );
  NAND3X1 U163 ( .A(n973), .B(n1828), .C(n1796), .Y(n1805) );
  OAI21X1 U164 ( .A(n1038), .B(n1007), .C(n1794), .Y(n1277) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1794) );
  OAI21X1 U166 ( .A(n1039), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1793) );
  OAI21X1 U168 ( .A(n1040), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1792) );
  OAI21X1 U170 ( .A(n1041), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1791) );
  OAI21X1 U172 ( .A(n1042), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1790) );
  OAI21X1 U174 ( .A(n1043), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1789) );
  OAI21X1 U176 ( .A(n1044), .B(n1006), .C(n1788), .Y(n1271) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1788) );
  OAI21X1 U178 ( .A(n1045), .B(n1006), .C(n1787), .Y(n1270) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1787) );
  NAND3X1 U180 ( .A(n1807), .B(n1828), .C(n1786), .Y(n1795) );
  OAI21X1 U181 ( .A(n1030), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1784) );
  OAI21X1 U183 ( .A(n1031), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1783) );
  OAI21X1 U185 ( .A(n1032), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1782) );
  OAI21X1 U187 ( .A(n1033), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1781) );
  OAI21X1 U189 ( .A(n1034), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1780) );
  OAI21X1 U191 ( .A(n1035), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1779) );
  OAI21X1 U193 ( .A(n1036), .B(n1005), .C(n1778), .Y(n1263) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1778) );
  OAI21X1 U195 ( .A(n1037), .B(n1005), .C(n1777), .Y(n1262) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1777) );
  NAND3X1 U197 ( .A(n973), .B(n1828), .C(n1776), .Y(n1785) );
  OAI21X1 U198 ( .A(n1038), .B(n1004), .C(n1774), .Y(n1261) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1774) );
  OAI21X1 U200 ( .A(n1039), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1773) );
  OAI21X1 U202 ( .A(n1040), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1772) );
  OAI21X1 U204 ( .A(n1041), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1771) );
  OAI21X1 U206 ( .A(n1042), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1770) );
  OAI21X1 U208 ( .A(n1043), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1769) );
  OAI21X1 U210 ( .A(n1044), .B(n1003), .C(n1768), .Y(n1255) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1768) );
  OAI21X1 U212 ( .A(n1045), .B(n1003), .C(n1767), .Y(n1254) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1767) );
  NAND3X1 U214 ( .A(n1806), .B(n1828), .C(n1766), .Y(n1775) );
  OAI21X1 U215 ( .A(n1030), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1764) );
  OAI21X1 U217 ( .A(n1031), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1763) );
  OAI21X1 U219 ( .A(n1032), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1762) );
  OAI21X1 U221 ( .A(n1033), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1761) );
  OAI21X1 U223 ( .A(n1034), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1760) );
  OAI21X1 U225 ( .A(n1035), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1759) );
  OAI21X1 U227 ( .A(n1036), .B(n1002), .C(n1758), .Y(n1247) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1758) );
  OAI21X1 U229 ( .A(n1037), .B(n1002), .C(n1757), .Y(n1246) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1757) );
  NAND3X1 U231 ( .A(n973), .B(n1828), .C(n1756), .Y(n1765) );
  OAI21X1 U232 ( .A(n1038), .B(n1001), .C(n1754), .Y(n1245) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1754) );
  OAI21X1 U234 ( .A(n1039), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1753) );
  OAI21X1 U236 ( .A(n1040), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1752) );
  OAI21X1 U238 ( .A(n1041), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1751) );
  OAI21X1 U240 ( .A(n1042), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1750) );
  OAI21X1 U242 ( .A(n1043), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1749) );
  OAI21X1 U244 ( .A(n1044), .B(n1000), .C(n1748), .Y(n1239) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1748) );
  OAI21X1 U246 ( .A(n1045), .B(n1000), .C(n1747), .Y(n1238) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1747) );
  NAND3X1 U248 ( .A(n1786), .B(n1828), .C(n1766), .Y(n1755) );
  OAI21X1 U249 ( .A(n1030), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1745) );
  OAI21X1 U251 ( .A(n1031), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1744) );
  OAI21X1 U253 ( .A(n1032), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1743) );
  OAI21X1 U255 ( .A(n1033), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1742) );
  OAI21X1 U257 ( .A(n1034), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1741) );
  OAI21X1 U259 ( .A(n1035), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1740) );
  OAI21X1 U261 ( .A(n1036), .B(n999), .C(n1739), .Y(n1231) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1739) );
  OAI21X1 U263 ( .A(n1037), .B(n999), .C(n1738), .Y(n1230) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1738) );
  NAND3X1 U265 ( .A(n973), .B(n1828), .C(n1737), .Y(n1746) );
  OAI21X1 U266 ( .A(n1038), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1735) );
  OAI21X1 U268 ( .A(n1039), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1734) );
  OAI21X1 U270 ( .A(n1040), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1733) );
  OAI21X1 U272 ( .A(n1041), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1732) );
  OAI21X1 U274 ( .A(n1042), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1731) );
  OAI21X1 U276 ( .A(n1043), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1730) );
  OAI21X1 U278 ( .A(n1044), .B(n998), .C(n1729), .Y(n1223) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1729) );
  OAI21X1 U280 ( .A(n1045), .B(n998), .C(n1728), .Y(n1222) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1728) );
  NAND3X1 U282 ( .A(n1806), .B(n1828), .C(n969), .Y(n1736) );
  OAI21X1 U283 ( .A(n1030), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1726) );
  OAI21X1 U285 ( .A(n1031), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1725) );
  OAI21X1 U287 ( .A(n1032), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1724) );
  OAI21X1 U289 ( .A(n1033), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1723) );
  OAI21X1 U291 ( .A(n1034), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1722) );
  OAI21X1 U293 ( .A(n1035), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1721) );
  OAI21X1 U295 ( .A(n1036), .B(n997), .C(n1720), .Y(n1215) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1720) );
  OAI21X1 U297 ( .A(n1037), .B(n997), .C(n1719), .Y(n1214) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1719) );
  NAND3X1 U299 ( .A(n973), .B(n1828), .C(n1718), .Y(n1727) );
  OAI21X1 U300 ( .A(n1038), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1716) );
  OAI21X1 U302 ( .A(n1039), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1715) );
  OAI21X1 U304 ( .A(n1040), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1714) );
  OAI21X1 U306 ( .A(n1041), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1713) );
  OAI21X1 U308 ( .A(n1042), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1712) );
  OAI21X1 U310 ( .A(n1043), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1711) );
  OAI21X1 U312 ( .A(n1044), .B(n996), .C(n1710), .Y(n1207) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1710) );
  OAI21X1 U314 ( .A(n1045), .B(n996), .C(n1709), .Y(n1206) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1709) );
  NAND3X1 U316 ( .A(n1786), .B(n1828), .C(n969), .Y(n1717) );
  OAI21X1 U317 ( .A(n1030), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1707) );
  OAI21X1 U319 ( .A(n1031), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1706) );
  OAI21X1 U321 ( .A(n1032), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1705) );
  OAI21X1 U323 ( .A(n1033), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1704) );
  OAI21X1 U325 ( .A(n1034), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1703) );
  OAI21X1 U327 ( .A(n1035), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1702) );
  OAI21X1 U329 ( .A(n1036), .B(n995), .C(n1701), .Y(n1199) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1701) );
  OAI21X1 U331 ( .A(n1037), .B(n995), .C(n1700), .Y(n1198) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1700) );
  NAND3X1 U333 ( .A(n973), .B(n1828), .C(n1699), .Y(n1708) );
  OAI21X1 U334 ( .A(n1038), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1697) );
  OAI21X1 U336 ( .A(n1039), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1696) );
  OAI21X1 U338 ( .A(n1040), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1695) );
  OAI21X1 U340 ( .A(n1041), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1694) );
  OAI21X1 U342 ( .A(n1042), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1693) );
  OAI21X1 U344 ( .A(n1043), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1692) );
  OAI21X1 U346 ( .A(n1044), .B(n994), .C(n1691), .Y(n1191) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1691) );
  OAI21X1 U348 ( .A(n1045), .B(n994), .C(n1690), .Y(n1190) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1690) );
  NAND3X1 U350 ( .A(n1806), .B(n1828), .C(n967), .Y(n1698) );
  OAI21X1 U351 ( .A(n1030), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1688) );
  OAI21X1 U353 ( .A(n1031), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1687) );
  OAI21X1 U355 ( .A(n1032), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1686) );
  OAI21X1 U357 ( .A(n1033), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1685) );
  OAI21X1 U359 ( .A(n1034), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1684) );
  OAI21X1 U361 ( .A(n1035), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1683) );
  OAI21X1 U363 ( .A(n1036), .B(n993), .C(n1682), .Y(n1183) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1682) );
  OAI21X1 U365 ( .A(n1037), .B(n993), .C(n1681), .Y(n1182) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1681) );
  NAND3X1 U367 ( .A(n973), .B(n1828), .C(n1680), .Y(n1689) );
  OAI21X1 U368 ( .A(n1038), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1678) );
  OAI21X1 U370 ( .A(n1039), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1677) );
  OAI21X1 U372 ( .A(n1040), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1676) );
  OAI21X1 U374 ( .A(n1041), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1675) );
  OAI21X1 U376 ( .A(n1042), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1674) );
  OAI21X1 U378 ( .A(n1043), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1673) );
  OAI21X1 U380 ( .A(n1044), .B(n992), .C(n1672), .Y(n1175) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1672) );
  OAI21X1 U382 ( .A(n1045), .B(n992), .C(n1671), .Y(n1174) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1671) );
  NAND3X1 U384 ( .A(n1786), .B(n1828), .C(n967), .Y(n1679) );
  OAI21X1 U385 ( .A(n1030), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1669) );
  OAI21X1 U387 ( .A(n1031), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1668) );
  OAI21X1 U389 ( .A(n1032), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1667) );
  OAI21X1 U391 ( .A(n1033), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1666) );
  OAI21X1 U393 ( .A(n1034), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1665) );
  OAI21X1 U395 ( .A(n1035), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1664) );
  OAI21X1 U397 ( .A(n1036), .B(n991), .C(n1663), .Y(n1167) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1663) );
  OAI21X1 U399 ( .A(n1037), .B(n991), .C(n1662), .Y(n1166) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1662) );
  NAND3X1 U401 ( .A(n973), .B(n1828), .C(n1661), .Y(n1670) );
  OAI21X1 U402 ( .A(n1038), .B(n990), .C(n1659), .Y(n1165) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1659) );
  OAI21X1 U404 ( .A(n1039), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1658) );
  OAI21X1 U406 ( .A(n1040), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1657) );
  OAI21X1 U408 ( .A(n1041), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1656) );
  OAI21X1 U410 ( .A(n1042), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1655) );
  OAI21X1 U412 ( .A(n1043), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1654) );
  OAI21X1 U414 ( .A(n1044), .B(n989), .C(n1653), .Y(n1159) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1653) );
  OAI21X1 U416 ( .A(n1045), .B(n989), .C(n1652), .Y(n1158) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1652) );
  NAND3X1 U418 ( .A(n1807), .B(n1828), .C(n1651), .Y(n1660) );
  OAI21X1 U419 ( .A(n1030), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1649) );
  OAI21X1 U421 ( .A(n1031), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1648) );
  OAI21X1 U423 ( .A(n1032), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1647) );
  OAI21X1 U425 ( .A(n1033), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1646) );
  OAI21X1 U427 ( .A(n1034), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1645) );
  OAI21X1 U429 ( .A(n1035), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1644) );
  OAI21X1 U431 ( .A(n1036), .B(n988), .C(n1643), .Y(n1151) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1643) );
  OAI21X1 U433 ( .A(n1037), .B(n988), .C(n1642), .Y(n1150) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1642) );
  NAND3X1 U435 ( .A(n973), .B(n1828), .C(n1641), .Y(n1650) );
  OAI21X1 U436 ( .A(n1038), .B(n987), .C(n1639), .Y(n1149) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1639) );
  OAI21X1 U438 ( .A(n1039), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1638) );
  OAI21X1 U440 ( .A(n1040), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1637) );
  OAI21X1 U442 ( .A(n1041), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1636) );
  OAI21X1 U444 ( .A(n1042), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1635) );
  OAI21X1 U446 ( .A(n1043), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1634) );
  OAI21X1 U448 ( .A(n1044), .B(n986), .C(n1633), .Y(n1143) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1633) );
  OAI21X1 U450 ( .A(n1045), .B(n986), .C(n1632), .Y(n1142) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1632) );
  NAND3X1 U452 ( .A(n1807), .B(n1828), .C(n1631), .Y(n1640) );
  OAI21X1 U453 ( .A(n1030), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1628) );
  OAI21X1 U455 ( .A(n1031), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1627) );
  OAI21X1 U457 ( .A(n1032), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1626) );
  OAI21X1 U459 ( .A(n1033), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1625) );
  OAI21X1 U461 ( .A(n1034), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1624) );
  OAI21X1 U463 ( .A(n1035), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1623) );
  OAI21X1 U465 ( .A(n1036), .B(n985), .C(n1622), .Y(n1135) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1622) );
  OAI21X1 U467 ( .A(n1037), .B(n985), .C(n1621), .Y(n1134) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1621) );
  NAND3X1 U469 ( .A(n973), .B(n1828), .C(n1620), .Y(n1629) );
  OAI21X1 U470 ( .A(n1038), .B(n984), .C(n1618), .Y(n1133) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1618) );
  OAI21X1 U472 ( .A(n1039), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1617) );
  OAI21X1 U474 ( .A(n1040), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1616) );
  OAI21X1 U476 ( .A(n1041), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1615) );
  OAI21X1 U478 ( .A(n1042), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1614) );
  OAI21X1 U480 ( .A(n1043), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1613) );
  OAI21X1 U482 ( .A(n1044), .B(n983), .C(n1612), .Y(n1127) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1612) );
  OAI21X1 U484 ( .A(n1045), .B(n983), .C(n1611), .Y(n1126) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1611) );
  NAND3X1 U486 ( .A(n1766), .B(n1828), .C(n1651), .Y(n1619) );
  OAI21X1 U487 ( .A(n1030), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1609) );
  OAI21X1 U489 ( .A(n1031), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1608) );
  OAI21X1 U491 ( .A(n1032), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1607) );
  OAI21X1 U493 ( .A(n1033), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1606) );
  OAI21X1 U495 ( .A(n1034), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1605) );
  OAI21X1 U497 ( .A(n1035), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1604) );
  OAI21X1 U499 ( .A(n1036), .B(n982), .C(n1603), .Y(n1119) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1603) );
  OAI21X1 U501 ( .A(n1037), .B(n982), .C(n1602), .Y(n1118) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1602) );
  NAND3X1 U503 ( .A(n973), .B(n1828), .C(n1601), .Y(n1610) );
  OAI21X1 U504 ( .A(n1038), .B(n981), .C(n1599), .Y(n1117) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1599) );
  OAI21X1 U506 ( .A(n1039), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1598) );
  OAI21X1 U508 ( .A(n1040), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1597) );
  OAI21X1 U510 ( .A(n1041), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1596) );
  OAI21X1 U512 ( .A(n1042), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1595) );
  OAI21X1 U514 ( .A(n1043), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1594) );
  OAI21X1 U516 ( .A(n1044), .B(n980), .C(n1593), .Y(n1111) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1593) );
  OAI21X1 U518 ( .A(n1045), .B(n980), .C(n1592), .Y(n1110) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1592) );
  NAND3X1 U520 ( .A(n1766), .B(n1828), .C(n1631), .Y(n1600) );
  OAI21X1 U521 ( .A(n1030), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1589) );
  OAI21X1 U523 ( .A(n1031), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1588) );
  OAI21X1 U525 ( .A(n1032), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1587) );
  OAI21X1 U527 ( .A(n1033), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1586) );
  OAI21X1 U529 ( .A(n1034), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1585) );
  OAI21X1 U531 ( .A(n1035), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1584) );
  OAI21X1 U533 ( .A(n1036), .B(n979), .C(n1583), .Y(n1103) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1583) );
  OAI21X1 U535 ( .A(n1037), .B(n979), .C(n1582), .Y(n1102) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1582) );
  NAND3X1 U537 ( .A(n973), .B(n1828), .C(n1581), .Y(n1590) );
  OAI21X1 U538 ( .A(n1038), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1579) );
  OAI21X1 U540 ( .A(n1039), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1578) );
  OAI21X1 U542 ( .A(n1040), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1577) );
  OAI21X1 U544 ( .A(n1041), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1576) );
  OAI21X1 U546 ( .A(n1042), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1575) );
  OAI21X1 U548 ( .A(n1043), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1574) );
  OAI21X1 U550 ( .A(n1044), .B(n978), .C(n1573), .Y(n1095) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1573) );
  OAI21X1 U552 ( .A(n1045), .B(n978), .C(n1572), .Y(n1094) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1572) );
  NAND3X1 U554 ( .A(n969), .B(n1828), .C(n1651), .Y(n1580) );
  OAI21X1 U555 ( .A(n1030), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1570) );
  OAI21X1 U557 ( .A(n1031), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1569) );
  OAI21X1 U559 ( .A(n1032), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1568) );
  OAI21X1 U561 ( .A(n1033), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1567) );
  OAI21X1 U563 ( .A(n1034), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1566) );
  OAI21X1 U565 ( .A(n1035), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1565) );
  OAI21X1 U567 ( .A(n1036), .B(n977), .C(n1564), .Y(n1087) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1564) );
  OAI21X1 U569 ( .A(n1037), .B(n977), .C(n1563), .Y(n1086) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1563) );
  NAND3X1 U571 ( .A(n973), .B(n1828), .C(n1562), .Y(n1571) );
  OAI21X1 U572 ( .A(n1038), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1560) );
  OAI21X1 U574 ( .A(n1039), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1559) );
  OAI21X1 U576 ( .A(n1040), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1558) );
  OAI21X1 U578 ( .A(n1041), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1557) );
  OAI21X1 U580 ( .A(n1042), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1556) );
  OAI21X1 U582 ( .A(n1043), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1555) );
  OAI21X1 U584 ( .A(n1044), .B(n976), .C(n1554), .Y(n1079) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1554) );
  OAI21X1 U586 ( .A(n1045), .B(n976), .C(n1553), .Y(n1078) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1553) );
  NAND3X1 U588 ( .A(n969), .B(n1828), .C(n1631), .Y(n1561) );
  OAI21X1 U590 ( .A(n1030), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1550) );
  OAI21X1 U592 ( .A(n1031), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1549) );
  OAI21X1 U594 ( .A(n1032), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1548) );
  OAI21X1 U596 ( .A(n1033), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1547) );
  OAI21X1 U598 ( .A(n1034), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1546) );
  OAI21X1 U600 ( .A(n1035), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1545) );
  OAI21X1 U602 ( .A(n1036), .B(n975), .C(n1544), .Y(n1071) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1544) );
  OAI21X1 U604 ( .A(n1037), .B(n975), .C(n1543), .Y(n1070) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1543) );
  NAND3X1 U606 ( .A(n973), .B(n1828), .C(n1542), .Y(n1551) );
  OAI21X1 U607 ( .A(n1038), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1540) );
  OAI21X1 U609 ( .A(n1039), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1539) );
  OAI21X1 U611 ( .A(n1040), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1538) );
  OAI21X1 U613 ( .A(n1041), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1537) );
  OAI21X1 U615 ( .A(n1042), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1536) );
  OAI21X1 U617 ( .A(n1043), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1535) );
  OAI21X1 U619 ( .A(n1044), .B(n974), .C(n1534), .Y(n1063) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1534) );
  OAI21X1 U621 ( .A(n1045), .B(n974), .C(n1533), .Y(n1062) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1533) );
  NAND3X1 U623 ( .A(n967), .B(n1828), .C(n1651), .Y(n1541) );
  OAI21X1 U624 ( .A(n1030), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1532) );
  OAI21X1 U626 ( .A(n1031), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1531) );
  OAI21X1 U628 ( .A(n1032), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1530) );
  OAI21X1 U630 ( .A(n1033), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1529) );
  OAI21X1 U632 ( .A(n1034), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1528) );
  OAI21X1 U634 ( .A(n1035), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1527) );
  OAI21X1 U636 ( .A(n1036), .B(n8), .C(n1526), .Y(n1055) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1526) );
  OAI21X1 U638 ( .A(n1037), .B(n8), .C(n1525), .Y(n1054) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1525) );
  NOR2X1 U641 ( .A(n964), .B(\addr_1c<4> ), .Y(n1818) );
  OAI21X1 U642 ( .A(n1038), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1522) );
  OAI21X1 U644 ( .A(n1039), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1521) );
  OAI21X1 U646 ( .A(n1040), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1520) );
  OAI21X1 U648 ( .A(n1041), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1519) );
  OAI21X1 U650 ( .A(n1042), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1518) );
  OAI21X1 U652 ( .A(n1043), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1517) );
  OAI21X1 U654 ( .A(n1044), .B(n972), .C(n1516), .Y(n1047) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1516) );
  OAI21X1 U656 ( .A(n1045), .B(n972), .C(n1515), .Y(n1046) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1515) );
  NAND3X1 U658 ( .A(n967), .B(n1828), .C(n1631), .Y(n1523) );
  NOR3X1 U661 ( .A(n1511), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1512) );
  NOR3X1 U662 ( .A(n1510), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1513) );
  AOI21X1 U663 ( .A(n461), .B(n1509), .C(n963), .Y(n1838) );
  OAI21X1 U665 ( .A(rd), .B(n1508), .C(wr), .Y(n1509) );
  NAND3X1 U667 ( .A(n1507), .B(n1025), .C(n1506), .Y(n1508) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1506) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1507) );
  AOI21X1 U670 ( .A(n448), .B(n1504), .C(n1024), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1503), .C(n4), .Y(n1504) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1786), .C(\mem<0><1> ), .D(n1631), .Y(
        n1501) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1806), .C(\mem<2><1> ), .D(n1651), .Y(
        n1502) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1786), .C(\mem<4><1> ), .D(n1631), .Y(
        n1499) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1806), .C(\mem<6><1> ), .D(n1651), .Y(
        n1500) );
  AOI22X1 U678 ( .A(n1591), .B(n892), .C(n1630), .D(n932), .Y(n1505) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1786), .C(\mem<12><1> ), .D(n1631), .Y(
        n1497) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1806), .C(\mem<14><1> ), .D(n1651), .Y(
        n1498) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1786), .C(\mem<8><1> ), .D(n1631), .Y(
        n1495) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1806), .C(\mem<10><1> ), .D(n1651), .Y(
        n1496) );
  AOI21X1 U685 ( .A(n447), .B(n1493), .C(n1024), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1491), .C(n950), .Y(n1493) );
  AOI21X1 U687 ( .A(n1489), .B(n1488), .C(n971), .Y(n1490) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1786), .C(\mem<0><0> ), .D(n1631), .Y(
        n1488) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1806), .C(\mem<2><0> ), .D(n1651), .Y(
        n1489) );
  AOI21X1 U690 ( .A(n1487), .B(n1486), .C(n970), .Y(n1492) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1786), .C(\mem<4><0> ), .D(n1631), .Y(
        n1486) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1806), .C(\mem<6><0> ), .D(n1651), .Y(
        n1487) );
  AOI22X1 U693 ( .A(n1591), .B(n890), .C(n1630), .D(n930), .Y(n1494) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1786), .C(\mem<12><0> ), .D(n1631), .Y(
        n1484) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1806), .C(\mem<14><0> ), .D(n1651), .Y(
        n1485) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1786), .C(\mem<8><0> ), .D(n1631), .Y(
        n1482) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1806), .C(\mem<10><0> ), .D(n1651), .Y(
        n1483) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1481) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1680), .C(\mem<19><7> ), .D(n1699), .Y(
        n1476) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1718), .C(\mem<23><7> ), .D(n1737), .Y(
        n1477) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1756), .C(\mem<27><7> ), .D(n1776), .Y(
        n1479) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1796), .C(\mem<31><7> ), .D(n1817), .Y(
        n1480) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1524), .C(\mem<3><7> ), .D(n1542), .Y(
        n1471) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1562), .C(\mem<7><7> ), .D(n1581), .Y(
        n1472) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1601), .C(\mem<11><7> ), .D(n1620), .Y(
        n1474) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1641), .C(\mem<15><7> ), .D(n1661), .Y(
        n1475) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1470) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1680), .C(\mem<19><6> ), .D(n1699), .Y(
        n1465) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1718), .C(\mem<23><6> ), .D(n1737), .Y(
        n1466) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1756), .C(\mem<27><6> ), .D(n1776), .Y(
        n1468) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1796), .C(\mem<31><6> ), .D(n1817), .Y(
        n1469) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1524), .C(\mem<3><6> ), .D(n1542), .Y(
        n1460) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1562), .C(\mem<7><6> ), .D(n1581), .Y(
        n1461) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1601), .C(\mem<11><6> ), .D(n1620), .Y(
        n1463) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1641), .C(\mem<15><6> ), .D(n1661), .Y(
        n1464) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1459) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1680), .C(\mem<19><5> ), .D(n1699), .Y(
        n1454) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1718), .C(\mem<23><5> ), .D(n1737), .Y(
        n1455) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1756), .C(\mem<27><5> ), .D(n1776), .Y(
        n1457) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1796), .C(\mem<31><5> ), .D(n1817), .Y(
        n1458) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1524), .C(\mem<3><5> ), .D(n1542), .Y(
        n1449) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1562), .C(\mem<7><5> ), .D(n1581), .Y(
        n1450) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1601), .C(\mem<11><5> ), .D(n1620), .Y(
        n1452) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1641), .C(\mem<15><5> ), .D(n1661), .Y(
        n1453) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1448) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1680), .C(\mem<19><4> ), .D(n1699), .Y(
        n1443) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1718), .C(\mem<23><4> ), .D(n1737), .Y(
        n1444) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1756), .C(\mem<27><4> ), .D(n1776), .Y(
        n1446) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1796), .C(\mem<31><4> ), .D(n1817), .Y(
        n1447) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1524), .C(\mem<3><4> ), .D(n1542), .Y(
        n1438) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1562), .C(\mem<7><4> ), .D(n1581), .Y(
        n1439) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1601), .C(\mem<11><4> ), .D(n1620), .Y(
        n1441) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1641), .C(\mem<15><4> ), .D(n1661), .Y(
        n1442) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1437) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1680), .C(\mem<19><3> ), .D(n1699), .Y(
        n1432) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1718), .C(\mem<23><3> ), .D(n1737), .Y(
        n1433) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1756), .C(\mem<27><3> ), .D(n1776), .Y(
        n1435) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1796), .C(\mem<31><3> ), .D(n1817), .Y(
        n1436) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1524), .C(\mem<3><3> ), .D(n1542), .Y(
        n1427) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1562), .C(\mem<7><3> ), .D(n1581), .Y(
        n1428) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1601), .C(\mem<11><3> ), .D(n1620), .Y(
        n1430) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1641), .C(\mem<15><3> ), .D(n1661), .Y(
        n1431) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1426) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1680), .C(\mem<19><2> ), .D(n1699), .Y(
        n1421) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1718), .C(\mem<23><2> ), .D(n1737), .Y(
        n1422) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1756), .C(\mem<27><2> ), .D(n1776), .Y(
        n1424) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1796), .C(\mem<31><2> ), .D(n1817), .Y(
        n1425) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1524), .C(\mem<3><2> ), .D(n1542), .Y(
        n1416) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1562), .C(\mem<7><2> ), .D(n1581), .Y(
        n1417) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1601), .C(\mem<11><2> ), .D(n1620), .Y(
        n1419) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1641), .C(\mem<15><2> ), .D(n1661), .Y(
        n1420) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1415) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1680), .C(\mem<19><1> ), .D(n1699), .Y(
        n1410) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1718), .C(\mem<23><1> ), .D(n1737), .Y(
        n1411) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1756), .C(\mem<27><1> ), .D(n1776), .Y(
        n1413) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1796), .C(\mem<31><1> ), .D(n1817), .Y(
        n1414) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1524), .C(\mem<3><1> ), .D(n1542), .Y(
        n1405) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1562), .C(\mem<7><1> ), .D(n1581), .Y(
        n1406) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1601), .C(\mem<11><1> ), .D(n1620), .Y(
        n1408) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1641), .C(\mem<15><1> ), .D(n1661), .Y(
        n1409) );
  AOI21X1 U777 ( .A(n435), .B(n1403), .C(n1024), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1401), .C(n949), .Y(n1403) );
  AOI21X1 U779 ( .A(n1399), .B(n1398), .C(n971), .Y(n1400) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1786), .C(\mem<0><7> ), .D(n1631), .Y(
        n1398) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1806), .C(\mem<2><7> ), .D(n1651), .Y(
        n1399) );
  AOI21X1 U782 ( .A(n1397), .B(n1396), .C(n970), .Y(n1402) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1786), .C(\mem<4><7> ), .D(n1631), .Y(
        n1396) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1806), .C(\mem<6><7> ), .D(n1651), .Y(
        n1397) );
  AOI22X1 U785 ( .A(n1591), .B(n888), .C(n1630), .D(n928), .Y(n1404) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1786), .C(\mem<12><7> ), .D(n1631), .Y(
        n1394) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1806), .C(\mem<14><7> ), .D(n1651), .Y(
        n1395) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1786), .C(\mem<8><7> ), .D(n1631), .Y(
        n1392) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1806), .C(\mem<10><7> ), .D(n1651), .Y(
        n1393) );
  AOI21X1 U792 ( .A(n434), .B(n1390), .C(n1024), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1388), .C(n948), .Y(n1390) );
  AOI21X1 U794 ( .A(n1386), .B(n1385), .C(n971), .Y(n1387) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1786), .C(\mem<0><6> ), .D(n1631), .Y(
        n1385) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1806), .C(\mem<2><6> ), .D(n1651), .Y(
        n1386) );
  AOI21X1 U797 ( .A(n1384), .B(n1383), .C(n970), .Y(n1389) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1786), .C(\mem<4><6> ), .D(n1631), .Y(
        n1383) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1806), .C(\mem<6><6> ), .D(n1651), .Y(
        n1384) );
  AOI22X1 U800 ( .A(n1591), .B(n886), .C(n1630), .D(n926), .Y(n1391) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1786), .C(\mem<12><6> ), .D(n1631), .Y(
        n1381) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1806), .C(\mem<14><6> ), .D(n1651), .Y(
        n1382) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1786), .C(\mem<8><6> ), .D(n1631), .Y(
        n1379) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1806), .C(\mem<10><6> ), .D(n1651), .Y(
        n1380) );
  AOI21X1 U807 ( .A(n422), .B(n1377), .C(n1024), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1375), .C(n947), .Y(n1377) );
  AOI21X1 U809 ( .A(n1373), .B(n1372), .C(n971), .Y(n1374) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1786), .C(\mem<0><5> ), .D(n1631), .Y(
        n1372) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1806), .C(\mem<2><5> ), .D(n1651), .Y(
        n1373) );
  AOI21X1 U812 ( .A(n1371), .B(n1370), .C(n970), .Y(n1376) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1786), .C(\mem<4><5> ), .D(n1631), .Y(
        n1370) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1806), .C(\mem<6><5> ), .D(n1651), .Y(
        n1371) );
  AOI22X1 U815 ( .A(n1591), .B(n884), .C(n1630), .D(n924), .Y(n1378) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1786), .C(\mem<12><5> ), .D(n1631), .Y(
        n1368) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1806), .C(\mem<14><5> ), .D(n1651), .Y(
        n1369) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1786), .C(\mem<8><5> ), .D(n1631), .Y(
        n1366) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1806), .C(\mem<10><5> ), .D(n1651), .Y(
        n1367) );
  AOI21X1 U822 ( .A(n421), .B(n1364), .C(n1024), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1362), .C(n946), .Y(n1364) );
  AOI21X1 U824 ( .A(n1360), .B(n1359), .C(n971), .Y(n1361) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1786), .C(\mem<0><4> ), .D(n1631), .Y(
        n1359) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1806), .C(\mem<2><4> ), .D(n1651), .Y(
        n1360) );
  AOI21X1 U827 ( .A(n1358), .B(n1357), .C(n970), .Y(n1363) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1786), .C(\mem<4><4> ), .D(n1631), .Y(
        n1357) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1806), .C(\mem<6><4> ), .D(n1651), .Y(
        n1358) );
  AOI22X1 U830 ( .A(n1591), .B(n882), .C(n1630), .D(n922), .Y(n1365) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1786), .C(\mem<12><4> ), .D(n1631), .Y(
        n1355) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1806), .C(\mem<14><4> ), .D(n1651), .Y(
        n1356) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1786), .C(\mem<8><4> ), .D(n1631), .Y(
        n1353) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1806), .C(\mem<10><4> ), .D(n1651), .Y(
        n1354) );
  AOI21X1 U837 ( .A(n409), .B(n1351), .C(n1024), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1349), .C(n945), .Y(n1351) );
  AOI21X1 U839 ( .A(n1347), .B(n1346), .C(n971), .Y(n1348) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1786), .C(\mem<0><3> ), .D(n1631), .Y(
        n1346) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1806), .C(\mem<2><3> ), .D(n1651), .Y(
        n1347) );
  AOI21X1 U842 ( .A(n1345), .B(n1344), .C(n970), .Y(n1350) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1786), .C(\mem<4><3> ), .D(n1631), .Y(
        n1344) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1806), .C(\mem<6><3> ), .D(n1651), .Y(
        n1345) );
  AOI22X1 U845 ( .A(n1591), .B(n880), .C(n1630), .D(n920), .Y(n1352) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1786), .C(\mem<12><3> ), .D(n1631), .Y(
        n1342) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1806), .C(\mem<14><3> ), .D(n1651), .Y(
        n1343) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1786), .C(\mem<8><3> ), .D(n1631), .Y(
        n1340) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1806), .C(\mem<10><3> ), .D(n1651), .Y(
        n1341) );
  AOI21X1 U852 ( .A(n408), .B(n1338), .C(n1024), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1336), .C(n944), .Y(n1338) );
  AOI21X1 U854 ( .A(n1334), .B(n1333), .C(n971), .Y(n1335) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1786), .C(\mem<0><2> ), .D(n1631), .Y(
        n1333) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1806), .C(\mem<2><2> ), .D(n1651), .Y(
        n1334) );
  AOI21X1 U857 ( .A(n1332), .B(n1331), .C(n970), .Y(n1337) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1786), .C(\mem<4><2> ), .D(n1631), .Y(
        n1331) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1806), .C(\mem<6><2> ), .D(n1651), .Y(
        n1332) );
  AOI22X1 U860 ( .A(n1591), .B(n878), .C(n1630), .D(n918), .Y(n1339) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1786), .C(\mem<12><2> ), .D(n1631), .Y(
        n1329) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1806), .C(\mem<14><2> ), .D(n1651), .Y(
        n1330) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1786), .C(\mem<8><2> ), .D(n1631), .Y(
        n1327) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1806), .C(\mem<10><2> ), .D(n1651), .Y(
        n1328) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1326) );
  NOR2X1 U868 ( .A(n1029), .B(\addr_1c<4> ), .Y(n1325) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1324) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1680), .C(\mem<19><0> ), .D(n1699), .Y(
        n1319) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1718), .C(\mem<23><0> ), .D(n1737), .Y(
        n1320) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1756), .C(\mem<27><0> ), .D(n1776), .Y(
        n1322) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1796), .C(\mem<31><0> ), .D(n1817), .Y(
        n1323) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1524), .C(\mem<3><0> ), .D(n1542), .Y(
        n1312) );
  NAND2X1 U877 ( .A(n1027), .B(n1028), .Y(n1514) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1562), .C(\mem<7><0> ), .D(n1581), .Y(
        n1313) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1028), .Y(n1552) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1601), .C(\mem<11><0> ), .D(n1620), .Y(
        n1315) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1641), .C(\mem<15><0> ), .D(n1661), .Y(
        n1316) );
  dff_50 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1012) );
  dff_49 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1012) );
  dff_48 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1012)
         );
  dff_47 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1012)
         );
  dff_46 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1012)
         );
  dff_45 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1012)
         );
  dff_44 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1012)
         );
  dff_43 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1012)
         );
  dff_42 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1012)
         );
  dff_41 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1012)
         );
  dff_40 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1012)
         );
  dff_39 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1012)
         );
  dff_38 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(n1012) );
  dff_37 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(n1012) );
  dff_36 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(n1012) );
  dff_35 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1012) );
  dff_34 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1012) );
  dff_33 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1012) );
  dff_32 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1012) );
  dff_31 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1012) );
  dff_30 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1012) );
  dff_29 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1012) );
  dff_28 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1012) );
  dff_27 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1012) );
  dff_26 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1012) );
  dff_25 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1012) );
  dff_24 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1012) );
  dff_23 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1012) );
  dff_22 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1012) );
  dff_21 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1012) );
  dff_20 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1012) );
  dff_19 \reg2[0]  ( .q(\data_out<0> ), .d(n1021), .clk(clk), .rst(n1012) );
  dff_18 \reg2[1]  ( .q(\data_out<1> ), .d(n1020), .clk(clk), .rst(n1012) );
  dff_17 \reg2[2]  ( .q(\data_out<2> ), .d(n1019), .clk(clk), .rst(n1012) );
  dff_16 \reg2[3]  ( .q(\data_out<3> ), .d(n1018), .clk(clk), .rst(n1012) );
  dff_15 \reg2[4]  ( .q(\data_out<4> ), .d(n1017), .clk(clk), .rst(n1012) );
  dff_14 \reg2[5]  ( .q(\data_out<5> ), .d(n1016), .clk(clk), .rst(n1012) );
  dff_13 \reg2[6]  ( .q(\data_out<6> ), .d(n1015), .clk(clk), .rst(n1012) );
  dff_12 \reg2[7]  ( .q(\data_out<7> ), .d(n1014), .clk(clk), .rst(n1012) );
  dff_11 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        n1012) );
  dff_10 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        n1012) );
  dff_9 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1012) );
  dff_8 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1012) );
  dff_7 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1012) );
  dff_6 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1012) );
  dff_5 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1012) );
  dff_4 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1012) );
  dff_3 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1012) );
  dff_2 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1012) );
  dff_1 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1012) );
  dff_0 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1012) );
  INVX1 U2 ( .A(rd), .Y(n1023) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1510) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n1524), .Y(n1827) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1029) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1028) );
  OR2X1 U7 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1511) );
  AND2X1 U8 ( .A(n1630), .B(n965), .Y(n1807) );
  AND2X1 U23 ( .A(n1591), .B(n965), .Y(n1766) );
  INVX1 U24 ( .A(\addr_1c<0> ), .Y(n1026) );
  AND2X1 U25 ( .A(n1026), .B(n1029), .Y(n1310) );
  AND2X1 U26 ( .A(\addr_1c<0> ), .B(n1029), .Y(n1311) );
  AND2X1 U27 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1318) );
  AND2X1 U28 ( .A(\addr_1c<3> ), .B(n1026), .Y(n1317) );
  INVX1 U29 ( .A(\addr_1c<1> ), .Y(n1027) );
  INVX1 U35 ( .A(wr1), .Y(n1025) );
  AND2X1 U36 ( .A(n1591), .B(n1318), .Y(n1776) );
  AND2X1 U37 ( .A(n1591), .B(n1317), .Y(n1756) );
  AND2X1 U38 ( .A(n940), .B(n1318), .Y(n1737) );
  AND2X1 U39 ( .A(n940), .B(n1317), .Y(n1718) );
  AND2X1 U40 ( .A(n1318), .B(n951), .Y(n1699) );
  AND2X1 U41 ( .A(n1317), .B(n951), .Y(n1680) );
  AND2X1 U42 ( .A(n1311), .B(n1591), .Y(n1620) );
  AND2X1 U43 ( .A(n1591), .B(n1310), .Y(n1601) );
  AND2X1 U44 ( .A(n1311), .B(n940), .Y(n1581) );
  AND2X1 U46 ( .A(n940), .B(n1310), .Y(n1562) );
  OR2X1 U47 ( .A(n970), .B(n964), .Y(n968) );
  AND2X1 U48 ( .A(n1311), .B(n951), .Y(n1542) );
  OR2X1 U49 ( .A(n964), .B(n971), .Y(n966) );
  AND2X1 U50 ( .A(n1630), .B(n1310), .Y(n1641) );
  AND2X1 U51 ( .A(n1311), .B(n1630), .Y(n1661) );
  AND2X1 U52 ( .A(n1317), .B(n1630), .Y(n1796) );
  AND2X1 U53 ( .A(\addr_1c<2> ), .B(n1027), .Y(n1591) );
  AND2X1 U54 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1630) );
  BUFX2 U55 ( .A(n961), .Y(n1010) );
  BUFX2 U56 ( .A(n961), .Y(n1009) );
  BUFX2 U57 ( .A(n960), .Y(n1007) );
  BUFX2 U58 ( .A(n960), .Y(n1006) );
  BUFX2 U59 ( .A(n959), .Y(n1004) );
  BUFX2 U60 ( .A(n959), .Y(n1003) );
  BUFX2 U61 ( .A(n958), .Y(n1001) );
  BUFX2 U62 ( .A(n958), .Y(n1000) );
  BUFX2 U63 ( .A(n957), .Y(n990) );
  BUFX2 U64 ( .A(n957), .Y(n989) );
  BUFX2 U65 ( .A(n956), .Y(n987) );
  BUFX2 U66 ( .A(n956), .Y(n986) );
  BUFX2 U67 ( .A(n955), .Y(n984) );
  BUFX2 U68 ( .A(n955), .Y(n983) );
  BUFX2 U69 ( .A(n954), .Y(n981) );
  BUFX2 U70 ( .A(n954), .Y(n980) );
  INVX1 U71 ( .A(\data_in_1c<0> ), .Y(n1030) );
  INVX1 U72 ( .A(\data_in_1c<1> ), .Y(n1031) );
  INVX1 U73 ( .A(\data_in_1c<2> ), .Y(n1032) );
  INVX1 U74 ( .A(\data_in_1c<3> ), .Y(n1033) );
  INVX1 U75 ( .A(\data_in_1c<4> ), .Y(n1034) );
  INVX1 U76 ( .A(\data_in_1c<5> ), .Y(n1035) );
  INVX1 U77 ( .A(\data_in_1c<6> ), .Y(n1036) );
  INVX1 U78 ( .A(\data_in_1c<7> ), .Y(n1037) );
  INVX1 U79 ( .A(\data_in_1c<8> ), .Y(n1038) );
  INVX1 U80 ( .A(\data_in_1c<9> ), .Y(n1039) );
  INVX1 U81 ( .A(\data_in_1c<10> ), .Y(n1040) );
  INVX1 U82 ( .A(\data_in_1c<11> ), .Y(n1041) );
  INVX1 U83 ( .A(\data_in_1c<12> ), .Y(n1042) );
  INVX1 U84 ( .A(\data_in_1c<13> ), .Y(n1043) );
  INVX1 U85 ( .A(\data_in_1c<14> ), .Y(n1044) );
  INVX1 U86 ( .A(\data_in_1c<15> ), .Y(n1045) );
  AND2X1 U87 ( .A(n1827), .B(\mem<32><0> ), .Y(n1491) );
  AND2X1 U88 ( .A(n1827), .B(\mem<32><1> ), .Y(n1503) );
  AND2X1 U89 ( .A(n1827), .B(\mem<32><2> ), .Y(n1336) );
  AND2X1 U90 ( .A(n1827), .B(\mem<32><3> ), .Y(n1349) );
  AND2X1 U91 ( .A(n1827), .B(\mem<32><4> ), .Y(n1362) );
  AND2X1 U92 ( .A(n1827), .B(\mem<32><5> ), .Y(n1375) );
  AND2X1 U93 ( .A(n1827), .B(\mem<32><6> ), .Y(n1388) );
  AND2X1 U129 ( .A(n1827), .B(\mem<32><7> ), .Y(n1401) );
  INVX1 U589 ( .A(rd1), .Y(n1024) );
  INVX1 U640 ( .A(wr), .Y(n1022) );
  INVX1 U659 ( .A(n1324), .Y(n1021) );
  INVX1 U660 ( .A(n1415), .Y(n1020) );
  INVX1 U664 ( .A(n1426), .Y(n1019) );
  INVX1 U666 ( .A(n1437), .Y(n1018) );
  INVX1 U672 ( .A(n1448), .Y(n1017) );
  INVX1 U675 ( .A(n1459), .Y(n1016) );
  INVX1 U679 ( .A(n1470), .Y(n1015) );
  INVX1 U682 ( .A(n1481), .Y(n1014) );
  AND2X1 U694 ( .A(wr1), .B(n1013), .Y(n1828) );
  INVX1 U697 ( .A(rst), .Y(n1013) );
  INVX2 U701 ( .A(n1013), .Y(n1012) );
  AND2X1 U706 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U712 ( .A(n1), .Y(n2) );
  AND2X1 U717 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U723 ( .A(n3), .Y(n4) );
  AND2X1 U728 ( .A(n1817), .B(n189), .Y(n5) );
  INVX1 U734 ( .A(n5), .Y(n6) );
  AND2X1 U739 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U745 ( .A(n7), .Y(n8) );
  OR2X1 U750 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U756 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U761 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U767 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U772 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U786 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U789 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U801 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U804 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U816 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U819 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U831 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U834 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U846 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U849 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U861 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U864 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U870 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U875 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U882 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U883 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U884 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U885 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U886 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U887 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U888 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U889 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U890 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U891 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U892 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U893 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U894 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U895 ( .A(n973), .B(n1828), .Y(n189) );
  AND2X1 U896 ( .A(n1828), .B(n1524), .Y(n289) );
  AND2X1 U897 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U898 ( .A(n348), .Y(n372) );
  AND2X1 U899 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U900 ( .A(n379), .Y(n381) );
  AND2X1 U901 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U902 ( .A(n386), .Y(n387) );
  AND2X1 U903 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U904 ( .A(n401), .Y(n402) );
  BUFX2 U905 ( .A(n1339), .Y(n408) );
  BUFX2 U906 ( .A(n1352), .Y(n409) );
  BUFX2 U907 ( .A(n1365), .Y(n421) );
  BUFX2 U908 ( .A(n1378), .Y(n422) );
  BUFX2 U909 ( .A(n1391), .Y(n434) );
  BUFX2 U910 ( .A(n1404), .Y(n435) );
  BUFX2 U911 ( .A(n1494), .Y(n447) );
  BUFX2 U912 ( .A(n1505), .Y(n448) );
  AND2X2 U913 ( .A(rd), .B(n1508), .Y(n460) );
  INVX1 U914 ( .A(n460), .Y(n461) );
  INVX1 U915 ( .A(n1314), .Y(n473) );
  INVX1 U916 ( .A(n1315), .Y(n474) );
  INVX1 U917 ( .A(n1316), .Y(n486) );
  INVX1 U918 ( .A(n1407), .Y(n487) );
  INVX1 U919 ( .A(n1408), .Y(n507) );
  INVX1 U920 ( .A(n1409), .Y(n508) );
  INVX1 U921 ( .A(n1418), .Y(n522) );
  INVX1 U922 ( .A(n1419), .Y(n523) );
  INVX1 U923 ( .A(n1420), .Y(n537) );
  INVX1 U924 ( .A(n1429), .Y(n538) );
  INVX1 U925 ( .A(n1430), .Y(n552) );
  INVX1 U926 ( .A(n1431), .Y(n553) );
  INVX1 U927 ( .A(n1440), .Y(n567) );
  INVX1 U928 ( .A(n1441), .Y(n568) );
  INVX1 U929 ( .A(n1442), .Y(n582) );
  INVX1 U930 ( .A(n1451), .Y(n583) );
  INVX1 U931 ( .A(n1452), .Y(n591) );
  INVX1 U932 ( .A(n1453), .Y(n592) );
  INVX1 U933 ( .A(n1462), .Y(n871) );
  INVX1 U934 ( .A(n1463), .Y(n872) );
  INVX1 U935 ( .A(n1464), .Y(n873) );
  INVX1 U936 ( .A(n1473), .Y(n874) );
  INVX1 U937 ( .A(n1474), .Y(n875) );
  INVX1 U938 ( .A(n1475), .Y(n876) );
  AND2X2 U939 ( .A(n1328), .B(n1327), .Y(n877) );
  INVX1 U940 ( .A(n877), .Y(n878) );
  AND2X2 U941 ( .A(n1341), .B(n1340), .Y(n879) );
  INVX1 U942 ( .A(n879), .Y(n880) );
  AND2X2 U943 ( .A(n1354), .B(n1353), .Y(n881) );
  INVX1 U944 ( .A(n881), .Y(n882) );
  AND2X2 U945 ( .A(n1367), .B(n1366), .Y(n883) );
  INVX1 U946 ( .A(n883), .Y(n884) );
  AND2X2 U947 ( .A(n1380), .B(n1379), .Y(n885) );
  INVX1 U948 ( .A(n885), .Y(n886) );
  AND2X2 U949 ( .A(n1393), .B(n1392), .Y(n887) );
  INVX1 U950 ( .A(n887), .Y(n888) );
  AND2X2 U951 ( .A(n1483), .B(n1482), .Y(n889) );
  INVX1 U952 ( .A(n889), .Y(n890) );
  AND2X2 U953 ( .A(n1496), .B(n1495), .Y(n891) );
  INVX1 U954 ( .A(n891), .Y(n892) );
  INVX1 U955 ( .A(n1321), .Y(n893) );
  INVX1 U956 ( .A(n1322), .Y(n894) );
  INVX1 U957 ( .A(n1323), .Y(n895) );
  INVX1 U958 ( .A(n1412), .Y(n896) );
  INVX1 U959 ( .A(n1413), .Y(n897) );
  INVX1 U960 ( .A(n1414), .Y(n898) );
  INVX1 U961 ( .A(n1423), .Y(n899) );
  INVX1 U962 ( .A(n1424), .Y(n900) );
  INVX1 U963 ( .A(n1425), .Y(n901) );
  INVX1 U964 ( .A(n1434), .Y(n902) );
  INVX1 U965 ( .A(n1435), .Y(n903) );
  INVX1 U966 ( .A(n1436), .Y(n904) );
  INVX1 U967 ( .A(n1445), .Y(n905) );
  INVX1 U968 ( .A(n1446), .Y(n906) );
  INVX1 U969 ( .A(n1447), .Y(n907) );
  INVX1 U970 ( .A(n1456), .Y(n908) );
  INVX1 U971 ( .A(n1457), .Y(n909) );
  INVX1 U972 ( .A(n1458), .Y(n910) );
  INVX1 U973 ( .A(n1467), .Y(n911) );
  INVX1 U974 ( .A(n1468), .Y(n912) );
  INVX1 U975 ( .A(n1469), .Y(n913) );
  INVX1 U976 ( .A(n1478), .Y(n914) );
  INVX1 U977 ( .A(n1479), .Y(n915) );
  INVX1 U978 ( .A(n1480), .Y(n916) );
  AND2X2 U979 ( .A(n1330), .B(n1329), .Y(n917) );
  INVX1 U980 ( .A(n917), .Y(n918) );
  AND2X2 U981 ( .A(n1343), .B(n1342), .Y(n919) );
  INVX1 U982 ( .A(n919), .Y(n920) );
  AND2X2 U983 ( .A(n1356), .B(n1355), .Y(n921) );
  INVX1 U984 ( .A(n921), .Y(n922) );
  AND2X2 U985 ( .A(n1369), .B(n1368), .Y(n923) );
  INVX1 U986 ( .A(n923), .Y(n924) );
  AND2X2 U987 ( .A(n1382), .B(n1381), .Y(n925) );
  INVX1 U988 ( .A(n925), .Y(n926) );
  AND2X2 U989 ( .A(n1395), .B(n1394), .Y(n927) );
  INVX1 U990 ( .A(n927), .Y(n928) );
  AND2X2 U991 ( .A(n1485), .B(n1484), .Y(n929) );
  INVX1 U992 ( .A(n929), .Y(n930) );
  AND2X2 U993 ( .A(n1498), .B(n1497), .Y(n931) );
  INVX1 U994 ( .A(n931), .Y(n932) );
  BUFX2 U995 ( .A(n1337), .Y(n933) );
  BUFX2 U996 ( .A(n1350), .Y(n934) );
  BUFX2 U997 ( .A(n1363), .Y(n935) );
  BUFX2 U998 ( .A(n1376), .Y(n936) );
  BUFX2 U999 ( .A(n1389), .Y(n937) );
  BUFX2 U1000 ( .A(n1402), .Y(n938) );
  BUFX2 U1001 ( .A(n1492), .Y(n939) );
  INVX1 U1002 ( .A(n970), .Y(n940) );
  INVX1 U1003 ( .A(n1499), .Y(n941) );
  INVX1 U1004 ( .A(n1500), .Y(n942) );
  BUFX2 U1005 ( .A(n1552), .Y(n970) );
  BUFX2 U1006 ( .A(n1838), .Y(err) );
  BUFX2 U1007 ( .A(n1335), .Y(n944) );
  BUFX2 U1008 ( .A(n1348), .Y(n945) );
  BUFX2 U1009 ( .A(n1361), .Y(n946) );
  BUFX2 U1010 ( .A(n1374), .Y(n947) );
  BUFX2 U1011 ( .A(n1387), .Y(n948) );
  BUFX2 U1012 ( .A(n1400), .Y(n949) );
  BUFX2 U1013 ( .A(n1490), .Y(n950) );
  INVX1 U1014 ( .A(n971), .Y(n951) );
  INVX1 U1015 ( .A(n1501), .Y(n952) );
  INVX1 U1016 ( .A(n1502), .Y(n953) );
  BUFX2 U1017 ( .A(n1514), .Y(n971) );
  BUFX2 U1018 ( .A(n1523), .Y(n972) );
  BUFX2 U1019 ( .A(n1541), .Y(n974) );
  BUFX2 U1020 ( .A(n1551), .Y(n975) );
  BUFX2 U1021 ( .A(n1561), .Y(n976) );
  BUFX2 U1022 ( .A(n1571), .Y(n977) );
  BUFX2 U1023 ( .A(n1580), .Y(n978) );
  BUFX2 U1024 ( .A(n1590), .Y(n979) );
  BUFX2 U1025 ( .A(n1610), .Y(n982) );
  BUFX2 U1026 ( .A(n1629), .Y(n985) );
  BUFX2 U1027 ( .A(n1650), .Y(n988) );
  BUFX2 U1028 ( .A(n1670), .Y(n991) );
  BUFX2 U1029 ( .A(n1679), .Y(n992) );
  BUFX2 U1030 ( .A(n1689), .Y(n993) );
  BUFX2 U1031 ( .A(n1698), .Y(n994) );
  BUFX2 U1032 ( .A(n1708), .Y(n995) );
  BUFX2 U1033 ( .A(n1717), .Y(n996) );
  BUFX2 U1034 ( .A(n1727), .Y(n997) );
  BUFX2 U1035 ( .A(n1736), .Y(n998) );
  BUFX2 U1036 ( .A(n1746), .Y(n999) );
  BUFX2 U1037 ( .A(n1765), .Y(n1002) );
  BUFX2 U1038 ( .A(n1785), .Y(n1005) );
  BUFX2 U1039 ( .A(n1805), .Y(n1008) );
  BUFX2 U1040 ( .A(n1818), .Y(n973) );
  AND2X1 U1041 ( .A(n1630), .B(n1318), .Y(n1817) );
  BUFX2 U1042 ( .A(n1837), .Y(n1011) );
  BUFX2 U1043 ( .A(n1600), .Y(n954) );
  BUFX2 U1044 ( .A(n1619), .Y(n955) );
  BUFX2 U1045 ( .A(n1640), .Y(n956) );
  BUFX2 U1046 ( .A(n1660), .Y(n957) );
  BUFX2 U1047 ( .A(n1755), .Y(n958) );
  BUFX2 U1048 ( .A(n1775), .Y(n959) );
  BUFX2 U1049 ( .A(n1795), .Y(n960) );
  BUFX2 U1050 ( .A(n1816), .Y(n961) );
  AND2X1 U1051 ( .A(enable), .B(n1013), .Y(n962) );
  INVX1 U1052 ( .A(n962), .Y(n963) );
  INVX1 U1053 ( .A(n965), .Y(n964) );
  AND2X1 U1054 ( .A(n1513), .B(n1512), .Y(n965) );
  INVX1 U1055 ( .A(n966), .Y(n967) );
  INVX1 U1056 ( .A(n968), .Y(n969) );
  AND2X1 U1057 ( .A(n951), .B(n1310), .Y(n1524) );
endmodule


module dff_212 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_213 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_214 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_215 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_208 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_209 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_210 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_211 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_204 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_205 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_206 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_207 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module cache_cache_id0 ( enable, clk, rst, createdump, .tag_in({\tag_in<4> , 
        \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), .index({
        \index<7> , \index<6> , \index<5> , \index<4> , \index<3> , \index<2> , 
        \index<1> , \index<0> }), .offset({\offset<2> , \offset<1> , 
        \offset<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), comp, write, 
        valid_in, .tag_out({\tag_out<4> , \tag_out<3> , \tag_out<2> , 
        \tag_out<1> , \tag_out<0> }), .data_out({\data_out<15> , 
        \data_out<14> , \data_out<13> , \data_out<12> , \data_out<11> , 
        \data_out<10> , \data_out<9> , \data_out<8> , \data_out<7> , 
        \data_out<6> , \data_out<5> , \data_out<4> , \data_out<3> , 
        \data_out<2> , \data_out<1> , \data_out<0> }), hit, dirty, valid, err
 );
  input enable, clk, rst, createdump, \tag_in<4> , \tag_in<3> , \tag_in<2> ,
         \tag_in<1> , \tag_in<0> , \index<7> , \index<6> , \index<5> ,
         \index<4> , \index<3> , \index<2> , \index<1> , \index<0> ,
         \offset<2> , \offset<1> , \offset<0> , \data_in<15> , \data_in<14> ,
         \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> ,
         \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> ,
         \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> ,
         comp, write, valid_in;
  output \tag_out<4> , \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , hit,
         dirty, valid, err;
  wire   n195, n196, n197, n198, wr_word0, \w0<15> , \w0<14> , \w0<13> ,
         \w0<12> , \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> ,
         \w0<5> , \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> , \w1<15> ,
         \w1<14> , \w1<13> , \w1<12> , \w1<11> , \w1<10> , \w1<9> , \w1<8> ,
         \w1<7> , \w1<6> , \w1<5> , \w1<4> , \w1<3> , \w1<2> , \w1<1> ,
         \w1<0> , \w2<15> , \w2<14> , \w2<13> , \w2<12> , \w2<11> , \w2<10> ,
         \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , \w2<4> , \w2<3> ,
         \w2<2> , \w2<1> , \w2<0> , \w3<15> , \w3<14> , \w3<13> , \w3<12> ,
         \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> ,
         \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> , dirtybit, validbit, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n23, n25, n27, n29, n31, n33, n35, n37, n39,
         n41, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n84, n86,
         n88, n90, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n117, n118, n119, n120, n121, n122, n124, n125, n126, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193;

  memc_Size16_7 mem_w0 ( .data_out({\w0<15> , \w0<14> , \w0<13> , \w0<12> , 
        \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> , 
        \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> }), .addr({n146, n144, n142, 
        n140, n138, n136, n134, n126}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(wr_word0), .clk(clk), .rst(n130), .createdump(createdump), 
        .file_id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  memc_Size16_6 mem_w1 ( .data_out({\w1<15> , \w1<14> , \w1<13> , \w1<12> , 
        \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , 
        \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> }), .addr({n146, n144, n142, 
        n140, n138, n136, n134, n126}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(n18), .clk(clk), .rst(n130), .createdump(createdump), .file_id(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b1}) );
  memc_Size16_5 mem_w2 ( .data_out({\w2<15> , \w2<14> , \w2<13> , \w2<12> , 
        \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , 
        \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> }), .addr({n146, n144, n142, 
        n140, n138, n136, n134, n126}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(n10), .clk(clk), .rst(n130), .createdump(createdump), .file_id(
        {1'b0, 1'b0, 1'b0, 1'b1, 1'b0}) );
  memc_Size16_4 mem_w3 ( .data_out({\w3<15> , \w3<14> , \w3<13> , \w3<12> , 
        \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , 
        \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> }), .addr({n146, n144, n142, 
        n140, n138, n136, n134, n126}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(n8), .clk(clk), .rst(n130), .createdump(createdump), .file_id({
        1'b0, 1'b0, 1'b0, 1'b1, 1'b1}) );
  memc_Size5_1 mem_tg ( .data_out({\tag_out<4> , n195, n196, n197, n198}), 
        .addr({n146, n144, n142, n140, n138, n136, n134, n124}), .data_in({
        \tag_in<4> , \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), 
        .write(n6), .clk(clk), .rst(n130), .createdump(createdump), .file_id({
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}) );
  memc_Size1_1 mem_dr ( .data_out(dirtybit), .addr({n146, n144, n142, n140, 
        n138, n136, n134, n126}), .data_in(comp), .write(n129), .clk(clk), 
        .rst(n130), .createdump(createdump), .file_id({1'b0, 1'b0, 1'b1, 1'b0, 
        1'b1}) );
  memv_1 mem_vl ( .data_out(validbit), .addr({n146, n144, n142, n140, n138, 
        n136, n134, n132}), .data_in(valid_in), .write(n128), .clk(clk), .rst(
        n130), .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  AND2X2 U3 ( .A(comp), .B(n125), .Y(n102) );
  AND2X1 U4 ( .A(n5), .B(n103), .Y(n1) );
  NOR2X1 U5 ( .A(n1), .B(n80), .Y(n193) );
  INVX2 U6 ( .A(n192), .Y(n2) );
  INVX1 U7 ( .A(\tag_in<3> ), .Y(n121) );
  INVX1 U8 ( .A(\tag_in<0> ), .Y(n3) );
  INVX1 U9 ( .A(n143), .Y(n142) );
  INVX1 U10 ( .A(\index<5> ), .Y(n143) );
  INVX1 U11 ( .A(\tag_in<2> ), .Y(n117) );
  INVX1 U12 ( .A(\tag_in<1> ), .Y(n118) );
  INVX1 U13 ( .A(n145), .Y(n144) );
  INVX1 U14 ( .A(\index<6> ), .Y(n145) );
  INVX1 U15 ( .A(n147), .Y(n146) );
  INVX1 U16 ( .A(\index<7> ), .Y(n147) );
  INVX1 U17 ( .A(comp), .Y(n153) );
  INVX1 U18 ( .A(\offset<0> ), .Y(n122) );
  INVX1 U19 ( .A(n122), .Y(err) );
  XNOR2X1 U20 ( .A(n198), .B(n3), .Y(n150) );
  BUFX2 U21 ( .A(n108), .Y(n4) );
  INVX1 U22 ( .A(n157), .Y(n5) );
  AND2X2 U23 ( .A(write), .B(n153), .Y(n92) );
  AND2X2 U24 ( .A(n108), .B(n92), .Y(n6) );
  OR2X2 U25 ( .A(n2), .B(n110), .Y(n7) );
  INVX1 U26 ( .A(n7), .Y(n8) );
  OR2X2 U27 ( .A(n2), .B(n99), .Y(n9) );
  INVX1 U28 ( .A(n9), .Y(n10) );
  OR2X2 U29 ( .A(n15), .B(n12), .Y(n11) );
  OR2X2 U30 ( .A(n20), .B(n19), .Y(n12) );
  OR2X2 U31 ( .A(n106), .B(n97), .Y(n13) );
  INVX1 U32 ( .A(n13), .Y(n14) );
  AND2X2 U33 ( .A(n78), .B(n65), .Y(n15) );
  OR2X2 U34 ( .A(\offset<2> ), .B(n158), .Y(n16) );
  OR2X2 U35 ( .A(n2), .B(n16), .Y(n17) );
  INVX1 U36 ( .A(n17), .Y(n18) );
  OR2X2 U37 ( .A(n149), .B(n148), .Y(n19) );
  OR2X2 U38 ( .A(n151), .B(n150), .Y(n20) );
  AND2X2 U39 ( .A(n66), .B(n53), .Y(n21) );
  INVX1 U40 ( .A(n21), .Y(\data_out<0> ) );
  AND2X2 U41 ( .A(n54), .B(n67), .Y(n23) );
  INVX1 U42 ( .A(n23), .Y(\data_out<1> ) );
  AND2X2 U43 ( .A(n55), .B(n68), .Y(n25) );
  INVX1 U44 ( .A(n25), .Y(\data_out<2> ) );
  AND2X2 U45 ( .A(n56), .B(n69), .Y(n27) );
  INVX1 U46 ( .A(n27), .Y(\data_out<5> ) );
  AND2X2 U47 ( .A(n70), .B(n57), .Y(n29) );
  INVX1 U48 ( .A(n29), .Y(\data_out<7> ) );
  AND2X2 U49 ( .A(n58), .B(n71), .Y(n31) );
  INVX1 U50 ( .A(n31), .Y(\data_out<8> ) );
  AND2X2 U51 ( .A(n59), .B(n72), .Y(n33) );
  INVX1 U52 ( .A(n33), .Y(\data_out<11> ) );
  AND2X2 U53 ( .A(n60), .B(n73), .Y(n35) );
  INVX1 U54 ( .A(n35), .Y(\data_out<12> ) );
  AND2X2 U55 ( .A(n61), .B(n74), .Y(n37) );
  INVX1 U56 ( .A(n37), .Y(\data_out<13> ) );
  AND2X2 U57 ( .A(n62), .B(n75), .Y(n39) );
  INVX1 U58 ( .A(n39), .Y(\data_out<14> ) );
  AND2X2 U59 ( .A(n76), .B(n63), .Y(n41) );
  INVX1 U60 ( .A(n41), .Y(\data_out<15> ) );
  BUFX2 U61 ( .A(n165), .Y(n43) );
  BUFX2 U62 ( .A(n168), .Y(n44) );
  BUFX2 U63 ( .A(n171), .Y(n45) );
  BUFX2 U64 ( .A(n178), .Y(n46) );
  BUFX2 U65 ( .A(n180), .Y(n47) );
  BUFX2 U66 ( .A(n166), .Y(n48) );
  BUFX2 U67 ( .A(n167), .Y(n49) );
  BUFX2 U68 ( .A(n172), .Y(n50) );
  BUFX2 U69 ( .A(n177), .Y(n51) );
  BUFX2 U70 ( .A(n179), .Y(n52) );
  BUFX2 U71 ( .A(n160), .Y(n53) );
  BUFX2 U72 ( .A(n161), .Y(n54) );
  BUFX2 U73 ( .A(n163), .Y(n55) );
  BUFX2 U74 ( .A(n169), .Y(n56) );
  BUFX2 U75 ( .A(n174), .Y(n57) );
  BUFX2 U76 ( .A(n175), .Y(n58) );
  BUFX2 U77 ( .A(n181), .Y(n59) );
  BUFX2 U78 ( .A(n183), .Y(n60) );
  BUFX2 U79 ( .A(n185), .Y(n61) );
  BUFX2 U80 ( .A(n187), .Y(n62) );
  BUFX2 U81 ( .A(n191), .Y(n63) );
  AND2X2 U82 ( .A(\tag_in<4> ), .B(\tag_out<4> ), .Y(n64) );
  INVX1 U83 ( .A(n64), .Y(n65) );
  BUFX2 U84 ( .A(n159), .Y(n66) );
  BUFX2 U85 ( .A(n162), .Y(n67) );
  BUFX2 U86 ( .A(n164), .Y(n68) );
  BUFX2 U87 ( .A(n170), .Y(n69) );
  BUFX2 U88 ( .A(n173), .Y(n70) );
  BUFX2 U89 ( .A(n176), .Y(n71) );
  BUFX2 U90 ( .A(n182), .Y(n72) );
  BUFX2 U91 ( .A(n184), .Y(n73) );
  BUFX2 U92 ( .A(n186), .Y(n74) );
  BUFX2 U93 ( .A(n188), .Y(n75) );
  BUFX2 U94 ( .A(n190), .Y(n76) );
  AND2X2 U95 ( .A(n119), .B(n120), .Y(n77) );
  INVX1 U96 ( .A(n77), .Y(n78) );
  AND2X2 U97 ( .A(enable), .B(n131), .Y(n108) );
  AND2X2 U98 ( .A(dirtybit), .B(n4), .Y(n79) );
  INVX1 U99 ( .A(n79), .Y(n80) );
  BUFX2 U100 ( .A(n193), .Y(dirty) );
  AND2X2 U101 ( .A(n43), .B(n48), .Y(n82) );
  INVX1 U102 ( .A(n82), .Y(\data_out<3> ) );
  AND2X2 U103 ( .A(n49), .B(n44), .Y(n84) );
  INVX1 U104 ( .A(n84), .Y(\data_out<4> ) );
  AND2X2 U105 ( .A(n45), .B(n50), .Y(n86) );
  INVX1 U106 ( .A(n86), .Y(\data_out<6> ) );
  AND2X2 U107 ( .A(n51), .B(n46), .Y(n88) );
  INVX1 U108 ( .A(n88), .Y(\data_out<9> ) );
  AND2X2 U109 ( .A(n52), .B(n47), .Y(n90) );
  INVX1 U110 ( .A(n90), .Y(\data_out<10> ) );
  INVX1 U111 ( .A(n92), .Y(n93) );
  AND2X2 U112 ( .A(n4), .B(n152), .Y(n94) );
  INVX1 U113 ( .A(n94), .Y(n95) );
  INVX1 U114 ( .A(n94), .Y(n96) );
  OR2X2 U115 ( .A(\offset<1> ), .B(n113), .Y(n97) );
  AND2X2 U116 ( .A(\offset<2> ), .B(n158), .Y(n98) );
  INVX1 U117 ( .A(n98), .Y(n99) );
  AND2X2 U118 ( .A(\offset<1> ), .B(n112), .Y(n100) );
  INVX1 U119 ( .A(n100), .Y(n101) );
  INVX1 U120 ( .A(n102), .Y(n103) );
  OR2X2 U121 ( .A(\offset<2> ), .B(n101), .Y(n104) );
  INVX1 U122 ( .A(n104), .Y(n105) );
  INVX1 U123 ( .A(\offset<2> ), .Y(n106) );
  AND2X1 U124 ( .A(n111), .B(n112), .Y(n107) );
  INVX1 U125 ( .A(n4), .Y(n109) );
  INVX1 U126 ( .A(n111), .Y(n110) );
  AND2X2 U127 ( .A(\offset<2> ), .B(\offset<1> ), .Y(n111) );
  AND2X1 U128 ( .A(n157), .B(n4), .Y(n112) );
  INVX1 U129 ( .A(n112), .Y(n113) );
  INVX8 U130 ( .A(\index<1> ), .Y(n135) );
  INVX1 U131 ( .A(\offset<1> ), .Y(n158) );
  BUFX2 U132 ( .A(n198), .Y(\tag_out<0> ) );
  INVX1 U133 ( .A(rst), .Y(n131) );
  BUFX2 U134 ( .A(n197), .Y(\tag_out<1> ) );
  BUFX2 U135 ( .A(n195), .Y(\tag_out<3> ) );
  XNOR2X1 U136 ( .A(n196), .B(n117), .Y(n149) );
  XNOR2X1 U137 ( .A(n197), .B(n118), .Y(n151) );
  INVX1 U138 ( .A(\tag_in<4> ), .Y(n119) );
  INVX1 U139 ( .A(\tag_out<4> ), .Y(n120) );
  XNOR2X1 U140 ( .A(n195), .B(n121), .Y(n148) );
  INVX1 U141 ( .A(write), .Y(n157) );
  INVX1 U142 ( .A(n133), .Y(n124) );
  BUFX2 U143 ( .A(n11), .Y(n125) );
  BUFX2 U144 ( .A(n132), .Y(n126) );
  INVX1 U145 ( .A(n133), .Y(n132) );
  BUFX2 U146 ( .A(n196), .Y(\tag_out<2> ) );
  INVX1 U147 ( .A(n96), .Y(hit) );
  INVX1 U148 ( .A(n11), .Y(n152) );
  BUFX2 U149 ( .A(n6), .Y(n128) );
  INVX1 U150 ( .A(\index<0> ), .Y(n133) );
  INVX1 U151 ( .A(n128), .Y(n154) );
  INVX1 U152 ( .A(n93), .Y(n156) );
  INVX1 U153 ( .A(n2), .Y(n129) );
  INVX8 U154 ( .A(n131), .Y(n130) );
  INVX8 U155 ( .A(n135), .Y(n134) );
  INVX8 U156 ( .A(n137), .Y(n136) );
  INVX8 U157 ( .A(\index<2> ), .Y(n137) );
  INVX8 U158 ( .A(n139), .Y(n138) );
  INVX8 U159 ( .A(\index<3> ), .Y(n139) );
  INVX8 U160 ( .A(n141), .Y(n140) );
  INVX8 U161 ( .A(\index<4> ), .Y(n141) );
  OAI21X1 U162 ( .A(n157), .B(n95), .C(n154), .Y(n192) );
  NOR3X1 U163 ( .A(\offset<2> ), .B(\offset<1> ), .C(n2), .Y(wr_word0) );
  INVX2 U164 ( .A(validbit), .Y(n155) );
  NOR3X1 U165 ( .A(n156), .B(n109), .C(n155), .Y(valid) );
  AOI22X1 U166 ( .A(n14), .B(\w2<0> ), .C(\w3<0> ), .D(n107), .Y(n160) );
  NOR3X1 U167 ( .A(\offset<2> ), .B(n113), .C(\offset<1> ), .Y(n189) );
  AOI22X1 U168 ( .A(n189), .B(\w0<0> ), .C(\w1<0> ), .D(n105), .Y(n159) );
  AOI22X1 U169 ( .A(n14), .B(\w2<1> ), .C(\w3<1> ), .D(n107), .Y(n162) );
  AOI22X1 U170 ( .A(n189), .B(\w0<1> ), .C(\w1<1> ), .D(n105), .Y(n161) );
  AOI22X1 U171 ( .A(n14), .B(\w2<2> ), .C(\w3<2> ), .D(n107), .Y(n164) );
  AOI22X1 U172 ( .A(n189), .B(\w0<2> ), .C(\w1<2> ), .D(n105), .Y(n163) );
  AOI22X1 U173 ( .A(n14), .B(\w2<3> ), .C(\w3<3> ), .D(n107), .Y(n166) );
  AOI22X1 U174 ( .A(n189), .B(\w0<3> ), .C(\w1<3> ), .D(n105), .Y(n165) );
  AOI22X1 U175 ( .A(n14), .B(\w2<4> ), .C(\w3<4> ), .D(n107), .Y(n168) );
  AOI22X1 U176 ( .A(n189), .B(\w0<4> ), .C(n105), .D(\w1<4> ), .Y(n167) );
  AOI22X1 U177 ( .A(n14), .B(\w2<5> ), .C(\w3<5> ), .D(n107), .Y(n170) );
  AOI22X1 U178 ( .A(n189), .B(\w0<5> ), .C(\w1<5> ), .D(n105), .Y(n169) );
  AOI22X1 U179 ( .A(n14), .B(\w2<6> ), .C(\w3<6> ), .D(n107), .Y(n172) );
  AOI22X1 U180 ( .A(n189), .B(\w0<6> ), .C(\w1<6> ), .D(n105), .Y(n171) );
  AOI22X1 U181 ( .A(n14), .B(\w2<7> ), .C(\w3<7> ), .D(n107), .Y(n174) );
  AOI22X1 U182 ( .A(n189), .B(\w0<7> ), .C(\w1<7> ), .D(n105), .Y(n173) );
  AOI22X1 U183 ( .A(n14), .B(\w2<8> ), .C(\w3<8> ), .D(n107), .Y(n176) );
  AOI22X1 U184 ( .A(n189), .B(\w0<8> ), .C(\w1<8> ), .D(n105), .Y(n175) );
  AOI22X1 U185 ( .A(n14), .B(\w2<9> ), .C(\w3<9> ), .D(n107), .Y(n178) );
  AOI22X1 U186 ( .A(n189), .B(\w0<9> ), .C(\w1<9> ), .D(n105), .Y(n177) );
  AOI22X1 U187 ( .A(n14), .B(\w2<10> ), .C(\w3<10> ), .D(n107), .Y(n180) );
  AOI22X1 U188 ( .A(n189), .B(\w0<10> ), .C(\w1<10> ), .D(n105), .Y(n179) );
  AOI22X1 U189 ( .A(n14), .B(\w2<11> ), .C(\w3<11> ), .D(n107), .Y(n182) );
  AOI22X1 U190 ( .A(n189), .B(\w0<11> ), .C(\w1<11> ), .D(n105), .Y(n181) );
  AOI22X1 U191 ( .A(n14), .B(\w2<12> ), .C(\w3<12> ), .D(n107), .Y(n184) );
  AOI22X1 U192 ( .A(n189), .B(\w0<12> ), .C(\w1<12> ), .D(n105), .Y(n183) );
  AOI22X1 U193 ( .A(n14), .B(\w2<13> ), .C(\w3<13> ), .D(n107), .Y(n186) );
  AOI22X1 U194 ( .A(n189), .B(\w0<13> ), .C(n105), .D(\w1<13> ), .Y(n185) );
  AOI22X1 U195 ( .A(n14), .B(\w2<14> ), .C(\w3<14> ), .D(n107), .Y(n188) );
  AOI22X1 U196 ( .A(n189), .B(\w0<14> ), .C(n105), .D(\w1<14> ), .Y(n187) );
  AOI22X1 U197 ( .A(n14), .B(\w2<15> ), .C(\w3<15> ), .D(n107), .Y(n191) );
  AOI22X1 U198 ( .A(n189), .B(\w0<15> ), .C(n105), .D(\w1<15> ), .Y(n190) );
endmodule


module cache_cache_id2 ( enable, clk, rst, createdump, .tag_in({\tag_in<4> , 
        \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), .index({
        \index<7> , \index<6> , \index<5> , \index<4> , \index<3> , \index<2> , 
        \index<1> , \index<0> }), .offset({\offset<2> , \offset<1> , 
        \offset<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), comp, write, 
        valid_in, .tag_out({\tag_out<4> , \tag_out<3> , \tag_out<2> , 
        \tag_out<1> , \tag_out<0> }), .data_out({\data_out<15> , 
        \data_out<14> , \data_out<13> , \data_out<12> , \data_out<11> , 
        \data_out<10> , \data_out<9> , \data_out<8> , \data_out<7> , 
        \data_out<6> , \data_out<5> , \data_out<4> , \data_out<3> , 
        \data_out<2> , \data_out<1> , \data_out<0> }), hit, dirty, valid, err
 );
  input enable, clk, rst, createdump, \tag_in<4> , \tag_in<3> , \tag_in<2> ,
         \tag_in<1> , \tag_in<0> , \index<7> , \index<6> , \index<5> ,
         \index<4> , \index<3> , \index<2> , \index<1> , \index<0> ,
         \offset<2> , \offset<1> , \offset<0> , \data_in<15> , \data_in<14> ,
         \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> ,
         \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> ,
         \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> ,
         comp, write, valid_in;
  output \tag_out<4> , \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , hit,
         dirty, valid, err;
  wire   \w0<15> , \w0<14> , \w0<13> , \w0<12> , \w0<11> , \w0<10> , \w0<9> ,
         \w0<8> , \w0<7> , \w0<6> , \w0<5> , \w0<4> , \w0<3> , \w0<2> ,
         \w0<1> , \w0<0> , \w1<15> , \w1<14> , \w1<13> , \w1<12> , \w1<11> ,
         \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , \w1<4> ,
         \w1<3> , \w1<2> , \w1<1> , \w1<0> , \w2<15> , \w2<14> , \w2<13> ,
         \w2<12> , \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> ,
         \w2<5> , \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> , \w3<15> ,
         \w3<14> , \w3<13> , \w3<12> , \w3<11> , \w3<10> , \w3<9> , \w3<8> ,
         \w3<7> , \w3<6> , \w3<5> , \w3<4> , \w3<3> , \w3<2> , \w3<1> ,
         \w3<0> , dirtybit, validbit, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25,
         n27, n29, n31, n33, n35, n37, n39, n41, n43, n45, n47, n49, n51, n53,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n190;

  memc_Size16_3 mem_w0 ( .data_out({\w0<15> , \w0<14> , \w0<13> , \w0<12> , 
        \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> , 
        \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> }), .addr({n138, n136, n134, 
        n132, n130, n128, n126, n113}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(n12), .clk(clk), .rst(n122), .createdump(createdump), .file_id(
        {1'b1, 1'b0, 1'b0, 1'b0, 1'b0}) );
  memc_Size16_2 mem_w1 ( .data_out({\w1<15> , \w1<14> , \w1<13> , \w1<12> , 
        \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , 
        \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> }), .addr({n138, n136, n134, 
        n132, n130, n128, n126, n114}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(n16), .clk(clk), .rst(n122), .createdump(createdump), .file_id(
        {1'b1, 1'b0, 1'b0, 1'b0, 1'b1}) );
  memc_Size16_1 mem_w2 ( .data_out({\w2<15> , \w2<14> , \w2<13> , \w2<12> , 
        \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , 
        \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> }), .addr({n138, n136, n134, 
        n132, n130, n128, n126, n114}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(n2), .clk(clk), .rst(n122), .createdump(createdump), .file_id({
        1'b1, 1'b0, 1'b0, 1'b1, 1'b0}) );
  memc_Size16_0 mem_w3 ( .data_out({\w3<15> , \w3<14> , \w3<13> , \w3<12> , 
        \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , 
        \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> }), .addr({n138, n136, n134, 
        n132, n130, n128, n126, n113}), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        .write(n3), .clk(clk), .rst(n122), .createdump(createdump), .file_id({
        1'b1, 1'b0, 1'b0, 1'b1, 1'b1}) );
  memc_Size5_0 mem_tg ( .data_out({\tag_out<4> , \tag_out<3> , \tag_out<2> , 
        \tag_out<1> , \tag_out<0> }), .addr({n138, n136, n134, n132, n130, 
        n128, n126, n124}), .data_in({\tag_in<4> , \tag_in<3> , \tag_in<2> , 
        \tag_in<1> , \tag_in<0> }), .write(n10), .clk(clk), .rst(n122), 
        .createdump(createdump), .file_id({1'b1, 1'b0, 1'b1, 1'b0, 1'b0}) );
  memc_Size1_0 mem_dr ( .data_out(dirtybit), .addr({n138, n136, n134, n132, 
        n130, n128, n126, n113}), .data_in(comp), .write(n121), .clk(clk), 
        .rst(n122), .createdump(createdump), .file_id({1'b1, 1'b0, 1'b1, 1'b0, 
        1'b1}) );
  memv_0 mem_vl ( .data_out(validbit), .addr({n138, n136, n134, n132, n130, 
        n128, n126, n114}), .data_in(valid_in), .write(n9), .clk(clk), .rst(
        n122), .createdump(createdump), .file_id({1'b1, 1'b0, 1'b0, 1'b0, 1'b0}) );
  AND2X2 U3 ( .A(comp), .B(n110), .Y(n99) );
  INVX1 U4 ( .A(\tag_in<3> ), .Y(n120) );
  INVX1 U5 ( .A(\tag_in<0> ), .Y(n7) );
  INVX1 U6 ( .A(\tag_in<2> ), .Y(n119) );
  INVX1 U7 ( .A(\tag_in<1> ), .Y(n115) );
  INVX1 U8 ( .A(n135), .Y(n134) );
  INVX1 U9 ( .A(\index<5> ), .Y(n135) );
  INVX1 U10 ( .A(n137), .Y(n136) );
  INVX1 U11 ( .A(\index<6> ), .Y(n137) );
  INVX1 U12 ( .A(n139), .Y(n138) );
  INVX1 U13 ( .A(\index<7> ), .Y(n139) );
  INVX1 U14 ( .A(rst), .Y(n123) );
  AND2X1 U15 ( .A(n111), .B(n149), .Y(n9) );
  INVX1 U16 ( .A(\offset<0> ), .Y(n117) );
  INVX1 U17 ( .A(n117), .Y(err) );
  XOR2X1 U18 ( .A(\tag_in<4> ), .B(\tag_out<4> ), .Y(n1) );
  AND2X2 U19 ( .A(n8), .B(n96), .Y(n2) );
  AND2X2 U20 ( .A(n8), .B(n22), .Y(n3) );
  INVX1 U21 ( .A(n151), .Y(n4) );
  INVX1 U22 ( .A(n147), .Y(n5) );
  INVX1 U23 ( .A(n5), .Y(n6) );
  XNOR2X1 U24 ( .A(\tag_out<0> ), .B(n7), .Y(n143) );
  INVX1 U25 ( .A(n147), .Y(n8) );
  AND2X2 U26 ( .A(n17), .B(n19), .Y(n10) );
  OR2X2 U27 ( .A(n147), .B(n107), .Y(n11) );
  INVX1 U28 ( .A(n11), .Y(n12) );
  OR2X2 U29 ( .A(n1), .B(n14), .Y(n13) );
  OR2X2 U30 ( .A(n21), .B(n20), .Y(n14) );
  OR2X2 U31 ( .A(n6), .B(n95), .Y(n15) );
  INVX1 U32 ( .A(n15), .Y(n16) );
  AND2X2 U33 ( .A(n123), .B(enable), .Y(n17) );
  INVX1 U34 ( .A(n17), .Y(n18) );
  AND2X2 U35 ( .A(write), .B(n140), .Y(n19) );
  OR2X2 U36 ( .A(n142), .B(n141), .Y(n20) );
  OR2X2 U37 ( .A(n144), .B(n143), .Y(n21) );
  AND2X2 U38 ( .A(\offset<2> ), .B(\offset<1> ), .Y(n22) );
  AND2X2 U39 ( .A(n55), .B(n71), .Y(n23) );
  INVX1 U40 ( .A(n23), .Y(\data_out<0> ) );
  AND2X2 U41 ( .A(n72), .B(n56), .Y(n25) );
  INVX1 U42 ( .A(n25), .Y(\data_out<1> ) );
  AND2X2 U43 ( .A(n73), .B(n57), .Y(n27) );
  INVX1 U44 ( .A(n27), .Y(\data_out<2> ) );
  AND2X2 U45 ( .A(n74), .B(n58), .Y(n29) );
  INVX1 U46 ( .A(n29), .Y(\data_out<3> ) );
  AND2X2 U47 ( .A(n75), .B(n59), .Y(n31) );
  INVX1 U48 ( .A(n31), .Y(\data_out<4> ) );
  AND2X2 U49 ( .A(n92), .B(n60), .Y(n33) );
  INVX1 U50 ( .A(n33), .Y(\data_out<5> ) );
  AND2X2 U51 ( .A(n76), .B(n61), .Y(n35) );
  INVX1 U52 ( .A(n35), .Y(\data_out<6> ) );
  AND2X2 U53 ( .A(n77), .B(n62), .Y(n37) );
  INVX1 U54 ( .A(n37), .Y(\data_out<7> ) );
  AND2X2 U55 ( .A(n78), .B(n63), .Y(n39) );
  INVX1 U56 ( .A(n39), .Y(\data_out<8> ) );
  AND2X2 U57 ( .A(n79), .B(n64), .Y(n41) );
  INVX1 U58 ( .A(n41), .Y(\data_out<9> ) );
  AND2X2 U59 ( .A(n80), .B(n65), .Y(n43) );
  INVX1 U60 ( .A(n43), .Y(\data_out<10> ) );
  AND2X2 U61 ( .A(n81), .B(n66), .Y(n45) );
  INVX1 U62 ( .A(n45), .Y(\data_out<11> ) );
  AND2X2 U63 ( .A(n82), .B(n67), .Y(n47) );
  INVX1 U64 ( .A(n47), .Y(\data_out<12> ) );
  AND2X2 U65 ( .A(n83), .B(n68), .Y(n49) );
  INVX1 U66 ( .A(n49), .Y(\data_out<13> ) );
  AND2X2 U67 ( .A(n84), .B(n69), .Y(n51) );
  INVX1 U68 ( .A(n51), .Y(\data_out<14> ) );
  AND2X2 U69 ( .A(n85), .B(n70), .Y(n53) );
  INVX1 U70 ( .A(n53), .Y(\data_out<15> ) );
  BUFX2 U71 ( .A(n155), .Y(n55) );
  BUFX2 U72 ( .A(n156), .Y(n56) );
  BUFX2 U73 ( .A(n158), .Y(n57) );
  BUFX2 U74 ( .A(n160), .Y(n58) );
  BUFX2 U75 ( .A(n162), .Y(n59) );
  BUFX2 U76 ( .A(n165), .Y(n60) );
  BUFX2 U77 ( .A(n166), .Y(n61) );
  BUFX2 U78 ( .A(n168), .Y(n62) );
  BUFX2 U79 ( .A(n170), .Y(n63) );
  BUFX2 U80 ( .A(n173), .Y(n64) );
  BUFX2 U81 ( .A(n174), .Y(n65) );
  BUFX2 U82 ( .A(n176), .Y(n66) );
  BUFX2 U83 ( .A(n178), .Y(n67) );
  BUFX2 U84 ( .A(n180), .Y(n68) );
  BUFX2 U85 ( .A(n182), .Y(n69) );
  BUFX2 U86 ( .A(n186), .Y(n70) );
  BUFX2 U87 ( .A(n154), .Y(n71) );
  BUFX2 U88 ( .A(n157), .Y(n72) );
  BUFX2 U89 ( .A(n159), .Y(n73) );
  BUFX2 U90 ( .A(n161), .Y(n74) );
  BUFX2 U91 ( .A(n163), .Y(n75) );
  BUFX2 U92 ( .A(n167), .Y(n76) );
  BUFX2 U93 ( .A(n169), .Y(n77) );
  BUFX2 U94 ( .A(n171), .Y(n78) );
  BUFX2 U95 ( .A(n172), .Y(n79) );
  BUFX2 U96 ( .A(n175), .Y(n80) );
  BUFX2 U97 ( .A(n177), .Y(n81) );
  BUFX2 U98 ( .A(n179), .Y(n82) );
  BUFX2 U99 ( .A(n181), .Y(n83) );
  BUFX2 U100 ( .A(n183), .Y(n84) );
  BUFX2 U101 ( .A(n187), .Y(n85) );
  AND2X2 U102 ( .A(n150), .B(dirtybit), .Y(n86) );
  INVX1 U103 ( .A(n86), .Y(n87) );
  INVX1 U104 ( .A(n93), .Y(n88) );
  AND2X2 U105 ( .A(n145), .B(n150), .Y(n93) );
  AND2X2 U106 ( .A(n150), .B(n116), .Y(n89) );
  INVX1 U107 ( .A(n89), .Y(n90) );
  INVX1 U108 ( .A(n164), .Y(n91) );
  INVX1 U109 ( .A(n91), .Y(n92) );
  INVX1 U110 ( .A(n89), .Y(n94) );
  OR2X2 U111 ( .A(\offset<2> ), .B(n152), .Y(n95) );
  AND2X2 U112 ( .A(\offset<2> ), .B(n152), .Y(n96) );
  INVX1 U113 ( .A(\offset<1> ), .Y(n152) );
  AND2X2 U114 ( .A(\offset<1> ), .B(n108), .Y(n97) );
  INVX1 U115 ( .A(n97), .Y(n98) );
  INVX1 U116 ( .A(n99), .Y(n100) );
  INVX1 U117 ( .A(n190), .Y(n101) );
  INVX1 U118 ( .A(n101), .Y(dirty) );
  OR2X2 U119 ( .A(\offset<2> ), .B(n98), .Y(n103) );
  INVX1 U120 ( .A(n103), .Y(n104) );
  INVX1 U121 ( .A(n153), .Y(n184) );
  AND2X1 U122 ( .A(n22), .B(n108), .Y(n105) );
  INVX1 U123 ( .A(n19), .Y(n106) );
  OR2X2 U124 ( .A(\offset<2> ), .B(\offset<1> ), .Y(n107) );
  AND2X1 U125 ( .A(n151), .B(n150), .Y(n108) );
  INVX1 U126 ( .A(n108), .Y(n109) );
  INVX1 U127 ( .A(n145), .Y(n110) );
  INVX1 U128 ( .A(n18), .Y(n111) );
  INVX1 U129 ( .A(n111), .Y(n112) );
  INVX1 U130 ( .A(n125), .Y(n113) );
  INVX1 U131 ( .A(n125), .Y(n114) );
  INVX1 U132 ( .A(n125), .Y(n124) );
  XNOR2X1 U133 ( .A(\tag_out<1> ), .B(n115), .Y(n144) );
  INVX1 U134 ( .A(n94), .Y(hit) );
  INVX1 U135 ( .A(n13), .Y(n116) );
  INVX4 U136 ( .A(\index<1> ), .Y(n127) );
  INVX1 U137 ( .A(write), .Y(n151) );
  INVX1 U138 ( .A(\index<0> ), .Y(n125) );
  XNOR2X1 U139 ( .A(\tag_out<2> ), .B(n119), .Y(n142) );
  XNOR2X1 U140 ( .A(\tag_out<3> ), .B(n120), .Y(n141) );
  INVX1 U141 ( .A(n13), .Y(n145) );
  OAI21X1 U142 ( .A(n88), .B(n151), .C(n146), .Y(n121) );
  INVX1 U143 ( .A(n9), .Y(n146) );
  INVX1 U144 ( .A(n112), .Y(n150) );
  INVX1 U145 ( .A(n106), .Y(n149) );
  INVX1 U146 ( .A(comp), .Y(n140) );
  INVX8 U147 ( .A(n123), .Y(n122) );
  INVX8 U148 ( .A(n127), .Y(n126) );
  INVX8 U149 ( .A(n129), .Y(n128) );
  INVX8 U150 ( .A(\index<2> ), .Y(n129) );
  INVX8 U151 ( .A(n131), .Y(n130) );
  INVX8 U152 ( .A(\index<3> ), .Y(n131) );
  INVX8 U153 ( .A(n133), .Y(n132) );
  INVX8 U154 ( .A(\index<4> ), .Y(n133) );
  OAI21X1 U155 ( .A(n151), .B(n90), .C(n146), .Y(n188) );
  INVX2 U156 ( .A(n188), .Y(n147) );
  INVX2 U157 ( .A(validbit), .Y(n148) );
  NOR3X1 U158 ( .A(n149), .B(n112), .C(n148), .Y(valid) );
  AOI21X1 U159 ( .A(n4), .B(n100), .C(n87), .Y(n190) );
  NAND3X1 U160 ( .A(\offset<2> ), .B(n108), .C(n152), .Y(n153) );
  AOI22X1 U161 ( .A(n184), .B(\w2<0> ), .C(n105), .D(\w3<0> ), .Y(n155) );
  NOR3X1 U162 ( .A(\offset<2> ), .B(n109), .C(\offset<1> ), .Y(n185) );
  AOI22X1 U163 ( .A(n185), .B(\w0<0> ), .C(n104), .D(\w1<0> ), .Y(n154) );
  AOI22X1 U164 ( .A(n184), .B(\w2<1> ), .C(n105), .D(\w3<1> ), .Y(n157) );
  AOI22X1 U165 ( .A(n185), .B(\w0<1> ), .C(n104), .D(\w1<1> ), .Y(n156) );
  AOI22X1 U166 ( .A(n184), .B(\w2<2> ), .C(n105), .D(\w3<2> ), .Y(n159) );
  AOI22X1 U167 ( .A(n185), .B(\w0<2> ), .C(n104), .D(\w1<2> ), .Y(n158) );
  AOI22X1 U168 ( .A(n184), .B(\w2<3> ), .C(n105), .D(\w3<3> ), .Y(n161) );
  AOI22X1 U169 ( .A(n185), .B(\w0<3> ), .C(n104), .D(\w1<3> ), .Y(n160) );
  AOI22X1 U170 ( .A(n184), .B(\w2<4> ), .C(n105), .D(\w3<4> ), .Y(n163) );
  AOI22X1 U171 ( .A(n185), .B(\w0<4> ), .C(n104), .D(\w1<4> ), .Y(n162) );
  AOI22X1 U172 ( .A(n184), .B(\w2<5> ), .C(n105), .D(\w3<5> ), .Y(n165) );
  AOI22X1 U173 ( .A(\w0<5> ), .B(n185), .C(\w1<5> ), .D(n104), .Y(n164) );
  AOI22X1 U174 ( .A(n184), .B(\w2<6> ), .C(n105), .D(\w3<6> ), .Y(n167) );
  AOI22X1 U175 ( .A(n185), .B(\w0<6> ), .C(n104), .D(\w1<6> ), .Y(n166) );
  AOI22X1 U176 ( .A(n184), .B(\w2<7> ), .C(n105), .D(\w3<7> ), .Y(n169) );
  AOI22X1 U177 ( .A(n185), .B(\w0<7> ), .C(n104), .D(\w1<7> ), .Y(n168) );
  AOI22X1 U178 ( .A(n184), .B(\w2<8> ), .C(n105), .D(\w3<8> ), .Y(n171) );
  AOI22X1 U179 ( .A(n185), .B(\w0<8> ), .C(n104), .D(\w1<8> ), .Y(n170) );
  AOI22X1 U180 ( .A(\w2<9> ), .B(n184), .C(n105), .D(\w3<9> ), .Y(n173) );
  AOI22X1 U181 ( .A(n185), .B(\w0<9> ), .C(n104), .D(\w1<9> ), .Y(n172) );
  AOI22X1 U182 ( .A(n184), .B(\w2<10> ), .C(\w3<10> ), .D(n105), .Y(n175) );
  AOI22X1 U183 ( .A(n185), .B(\w0<10> ), .C(n104), .D(\w1<10> ), .Y(n174) );
  AOI22X1 U184 ( .A(n184), .B(\w2<11> ), .C(n105), .D(\w3<11> ), .Y(n177) );
  AOI22X1 U185 ( .A(n185), .B(\w0<11> ), .C(n104), .D(\w1<11> ), .Y(n176) );
  AOI22X1 U186 ( .A(n184), .B(\w2<12> ), .C(n105), .D(\w3<12> ), .Y(n179) );
  AOI22X1 U187 ( .A(n185), .B(\w0<12> ), .C(n104), .D(\w1<12> ), .Y(n178) );
  AOI22X1 U188 ( .A(n184), .B(\w2<13> ), .C(\w3<13> ), .D(n105), .Y(n181) );
  AOI22X1 U189 ( .A(n185), .B(\w0<13> ), .C(n104), .D(\w1<13> ), .Y(n180) );
  AOI22X1 U190 ( .A(n184), .B(\w2<14> ), .C(n105), .D(\w3<14> ), .Y(n183) );
  AOI22X1 U191 ( .A(n185), .B(\w0<14> ), .C(n104), .D(\w1<14> ), .Y(n182) );
  AOI22X1 U192 ( .A(n184), .B(\w2<15> ), .C(n105), .D(\w3<15> ), .Y(n187) );
  AOI22X1 U193 ( .A(\w0<15> ), .B(n185), .C(n104), .D(\w1<15> ), .Y(n186) );
endmodule


module four_bank_mem ( clk, rst, createdump, .addr({\addr<15> , \addr<14> , 
        \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> , 
        \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> , 
        \addr<1> , \addr<0> }), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        wr, rd, .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), stall, .busy({\busy<3> , \busy<2> , \busy<1> , 
        \busy<0> }), err );
  input clk, rst, createdump, \addr<15> , \addr<14> , \addr<13> , \addr<12> ,
         \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> ,
         \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> ,
         \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , wr, rd;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , stall,
         \busy<3> , \busy<2> , \busy<1> , \busy<0> , err;
  wire   \en<3> , \en<2> , \en<1> , \en<0> , \data0_out<15> , \data0_out<14> ,
         \data0_out<13> , \data0_out<12> , \data0_out<11> , \data0_out<10> ,
         \data0_out<9> , \data0_out<8> , \data0_out<7> , \data0_out<6> ,
         \data0_out<5> , \data0_out<4> , \data0_out<3> , \data0_out<2> ,
         \data0_out<1> , \data0_out<0> , err0, \data1_out<15> ,
         \data1_out<14> , \data1_out<13> , \data1_out<12> , \data1_out<11> ,
         \data1_out<10> , \data1_out<9> , \data1_out<8> , \data1_out<7> ,
         \data1_out<6> , \data1_out<5> , \data1_out<4> , \data1_out<3> ,
         \data1_out<2> , \data1_out<1> , \data1_out<0> , err1, \data2_out<15> ,
         \data2_out<14> , \data2_out<13> , \data2_out<12> , \data2_out<11> ,
         \data2_out<10> , \data2_out<9> , \data2_out<8> , \data2_out<7> ,
         \data2_out<6> , \data2_out<5> , \data2_out<4> , \data2_out<3> ,
         \data2_out<2> , \data2_out<1> , \data2_out<0> , err2, \data3_out<15> ,
         \data3_out<14> , \data3_out<13> , \data3_out<12> , \data3_out<11> ,
         \data3_out<10> , \data3_out<9> , \data3_out<8> , \data3_out<7> ,
         \data3_out<6> , \data3_out<5> , \data3_out<4> , \data3_out<3> ,
         \data3_out<2> , \data3_out<1> , \data3_out<0> , err3, \bsy0<3> ,
         \bsy0<2> , \bsy0<1> , \bsy0<0> , \bsy1<3> , \bsy1<2> , \bsy1<1> ,
         \bsy1<0> , \bsy2<3> , \bsy2<2> , \bsy2<1> , \bsy2<0> , n9, n10, n11,
         n13, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n1, n2, n3, n4, n5, n6, n7,
         n8, n12, n14, n15, n17, n18, n19, n21, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85,
         n87, n89, n91, n93, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114;

  NOR3X1 U9 ( .A(n96), .B(rst), .C(n2), .Y(stall) );
  OAI21X1 U11 ( .A(\addr<1> ), .B(n11), .C(n6), .Y(n10) );
  OAI21X1 U13 ( .A(\addr<1> ), .B(n13), .C(n4), .Y(n9) );
  AOI21X1 U15 ( .A(n17), .B(n16), .C(n96), .Y(err) );
  NOR3X1 U16 ( .A(err1), .B(err3), .C(err2), .Y(n16) );
  NOR3X1 U18 ( .A(n59), .B(\busy<3> ), .C(n96), .Y(\en<3> ) );
  NOR3X1 U20 ( .A(n57), .B(n96), .C(n114), .Y(\en<2> ) );
  NOR3X1 U22 ( .A(n55), .B(n96), .C(n113), .Y(\en<1> ) );
  NOR3X1 U24 ( .A(n19), .B(\busy<0> ), .C(n96), .Y(\en<0> ) );
  NOR2X1 U28 ( .A(\data3_out<9> ), .B(\data2_out<9> ), .Y(n23) );
  NOR2X1 U29 ( .A(\data1_out<9> ), .B(\data0_out<9> ), .Y(n22) );
  NOR2X1 U31 ( .A(\data3_out<8> ), .B(\data2_out<8> ), .Y(n25) );
  NOR2X1 U32 ( .A(\data1_out<8> ), .B(\data0_out<8> ), .Y(n24) );
  NOR2X1 U34 ( .A(\data3_out<7> ), .B(\data2_out<7> ), .Y(n27) );
  NOR2X1 U35 ( .A(\data1_out<7> ), .B(\data0_out<7> ), .Y(n26) );
  NOR2X1 U37 ( .A(\data3_out<6> ), .B(\data2_out<6> ), .Y(n29) );
  NOR2X1 U38 ( .A(\data1_out<6> ), .B(\data0_out<6> ), .Y(n28) );
  NOR2X1 U40 ( .A(\data3_out<5> ), .B(\data2_out<5> ), .Y(n31) );
  NOR2X1 U41 ( .A(\data1_out<5> ), .B(\data0_out<5> ), .Y(n30) );
  NOR2X1 U43 ( .A(\data3_out<4> ), .B(\data2_out<4> ), .Y(n33) );
  NOR2X1 U44 ( .A(\data1_out<4> ), .B(\data0_out<4> ), .Y(n32) );
  NOR2X1 U46 ( .A(\data3_out<3> ), .B(\data2_out<3> ), .Y(n35) );
  NOR2X1 U47 ( .A(\data1_out<3> ), .B(\data0_out<3> ), .Y(n34) );
  NOR2X1 U49 ( .A(\data3_out<2> ), .B(\data2_out<2> ), .Y(n37) );
  NOR2X1 U50 ( .A(\data1_out<2> ), .B(\data0_out<2> ), .Y(n36) );
  NOR2X1 U52 ( .A(\data3_out<1> ), .B(\data2_out<1> ), .Y(n39) );
  NOR2X1 U53 ( .A(\data1_out<1> ), .B(\data0_out<1> ), .Y(n38) );
  NOR2X1 U55 ( .A(\data3_out<15> ), .B(\data2_out<15> ), .Y(n41) );
  NOR2X1 U56 ( .A(\data1_out<15> ), .B(\data0_out<15> ), .Y(n40) );
  NOR2X1 U58 ( .A(\data3_out<14> ), .B(\data2_out<14> ), .Y(n43) );
  NOR2X1 U59 ( .A(\data1_out<14> ), .B(\data0_out<14> ), .Y(n42) );
  NOR2X1 U61 ( .A(\data3_out<13> ), .B(\data2_out<13> ), .Y(n45) );
  NOR2X1 U62 ( .A(\data1_out<13> ), .B(\data0_out<13> ), .Y(n44) );
  NOR2X1 U64 ( .A(\data3_out<12> ), .B(\data2_out<12> ), .Y(n47) );
  NOR2X1 U65 ( .A(\data1_out<12> ), .B(\data0_out<12> ), .Y(n46) );
  NOR2X1 U67 ( .A(\data3_out<11> ), .B(\data2_out<11> ), .Y(n49) );
  NOR2X1 U68 ( .A(\data1_out<11> ), .B(\data0_out<11> ), .Y(n48) );
  NOR2X1 U70 ( .A(\data3_out<10> ), .B(\data2_out<10> ), .Y(n51) );
  NOR2X1 U71 ( .A(\data1_out<10> ), .B(\data0_out<10> ), .Y(n50) );
  NOR2X1 U73 ( .A(\data3_out<0> ), .B(\data2_out<0> ), .Y(n53) );
  NOR2X1 U74 ( .A(\data1_out<0> ), .B(\data0_out<0> ), .Y(n52) );
  NOR3X1 U75 ( .A(\bsy0<3> ), .B(\bsy2<3> ), .C(\bsy1<3> ), .Y(n54) );
  NOR3X1 U76 ( .A(\bsy0<2> ), .B(\bsy2<2> ), .C(\bsy1<2> ), .Y(n11) );
  NOR3X1 U77 ( .A(\bsy0<1> ), .B(\bsy2<1> ), .C(\bsy1<1> ), .Y(n20) );
  NOR3X1 U78 ( .A(\bsy0<0> ), .B(\bsy2<0> ), .C(\bsy1<0> ), .Y(n13) );
  final_memory_3 m0 ( .data_out({\data0_out<15> , \data0_out<14> , 
        \data0_out<13> , \data0_out<12> , \data0_out<11> , \data0_out<10> , 
        \data0_out<9> , \data0_out<8> , \data0_out<7> , \data0_out<6> , 
        \data0_out<5> , \data0_out<4> , \data0_out<3> , \data0_out<2> , 
        \data0_out<1> , \data0_out<0> }), .err(err0), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n111, n109, n107, n105, n103, n101, n99, n97}), .wr(wr), 
        .rd(rd), .enable(\en<0> ), .create_dump(createdump), .bank_id({1'b0, 
        1'b0}), .clk(clk), .rst(rst) );
  final_memory_2 m1 ( .data_out({\data1_out<15> , \data1_out<14> , 
        \data1_out<13> , \data1_out<12> , \data1_out<11> , \data1_out<10> , 
        \data1_out<9> , \data1_out<8> , \data1_out<7> , \data1_out<6> , 
        \data1_out<5> , \data1_out<4> , \data1_out<3> , \data1_out<2> , 
        \data1_out<1> , \data1_out<0> }), .err(err1), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n111, n109, n107, n105, n103, n101, n99, n97}), .wr(wr), 
        .rd(rd), .enable(\en<1> ), .create_dump(createdump), .bank_id({1'b0, 
        1'b1}), .clk(clk), .rst(rst) );
  final_memory_1 m2 ( .data_out({\data2_out<15> , \data2_out<14> , 
        \data2_out<13> , \data2_out<12> , \data2_out<11> , \data2_out<10> , 
        \data2_out<9> , \data2_out<8> , \data2_out<7> , \data2_out<6> , 
        \data2_out<5> , \data2_out<4> , \data2_out<3> , \data2_out<2> , 
        \data2_out<1> , \data2_out<0> }), .err(err2), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n111, n109, n107, n105, n103, n101, n99, n97}), .wr(wr), 
        .rd(rd), .enable(\en<2> ), .create_dump(createdump), .bank_id({1'b1, 
        1'b0}), .clk(clk), .rst(rst) );
  final_memory_0 m3 ( .data_out({\data3_out<15> , \data3_out<14> , 
        \data3_out<13> , \data3_out<12> , \data3_out<11> , \data3_out<10> , 
        \data3_out<9> , \data3_out<8> , \data3_out<7> , \data3_out<6> , 
        \data3_out<5> , \data3_out<4> , \data3_out<3> , \data3_out<2> , 
        \data3_out<1> , \data3_out<0> }), .err(err3), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , n111, n109, n107, n105, n103, n101, n99, n97}), .wr(wr), 
        .rd(rd), .enable(\en<3> ), .create_dump(createdump), .bank_id({1'b1, 
        1'b1}), .clk(clk), .rst(rst) );
  dff_212 \b0[0]  ( .q(\bsy0<0> ), .d(\en<0> ), .clk(clk), .rst(rst) );
  dff_213 \b0[1]  ( .q(\bsy0<1> ), .d(\en<1> ), .clk(clk), .rst(rst) );
  dff_214 \b0[2]  ( .q(\bsy0<2> ), .d(\en<2> ), .clk(clk), .rst(rst) );
  dff_215 \b0[3]  ( .q(\bsy0<3> ), .d(\en<3> ), .clk(clk), .rst(rst) );
  dff_208 \b1[0]  ( .q(\bsy1<0> ), .d(\bsy0<0> ), .clk(clk), .rst(rst) );
  dff_209 \b1[1]  ( .q(\bsy1<1> ), .d(\bsy0<1> ), .clk(clk), .rst(rst) );
  dff_210 \b1[2]  ( .q(\bsy1<2> ), .d(\bsy0<2> ), .clk(clk), .rst(rst) );
  dff_211 \b1[3]  ( .q(\bsy1<3> ), .d(\bsy0<3> ), .clk(clk), .rst(rst) );
  dff_204 \b2[0]  ( .q(\bsy2<0> ), .d(\bsy1<0> ), .clk(clk), .rst(rst) );
  dff_205 \b2[1]  ( .q(\bsy2<1> ), .d(\bsy1<1> ), .clk(clk), .rst(rst) );
  dff_206 \b2[2]  ( .q(\bsy2<2> ), .d(\bsy1<2> ), .clk(clk), .rst(rst) );
  dff_207 \b2[3]  ( .q(\bsy2<3> ), .d(\bsy1<3> ), .clk(clk), .rst(rst) );
  INVX4 U3 ( .A(\addr<2> ), .Y(n114) );
  INVX1 U4 ( .A(n13), .Y(\busy<0> ) );
  INVX1 U5 ( .A(n54), .Y(\busy<3> ) );
  INVX1 U6 ( .A(n98), .Y(n97) );
  INVX1 U7 ( .A(n100), .Y(n99) );
  INVX1 U8 ( .A(n102), .Y(n101) );
  INVX1 U10 ( .A(\addr<5> ), .Y(n102) );
  INVX1 U12 ( .A(n104), .Y(n103) );
  INVX1 U14 ( .A(\addr<6> ), .Y(n104) );
  INVX1 U17 ( .A(n106), .Y(n105) );
  INVX1 U19 ( .A(\addr<7> ), .Y(n106) );
  INVX1 U21 ( .A(n108), .Y(n107) );
  INVX1 U23 ( .A(\addr<8> ), .Y(n108) );
  INVX1 U25 ( .A(n110), .Y(n109) );
  INVX1 U26 ( .A(\addr<9> ), .Y(n110) );
  INVX1 U27 ( .A(n112), .Y(n111) );
  INVX1 U30 ( .A(\addr<10> ), .Y(n112) );
  OR2X1 U33 ( .A(rd), .B(wr), .Y(n95) );
  INVX1 U36 ( .A(n20), .Y(\busy<1> ) );
  OR2X1 U39 ( .A(err0), .B(\addr<0> ), .Y(n15) );
  INVX1 U42 ( .A(n11), .Y(\busy<2> ) );
  OR2X2 U45 ( .A(n8), .B(n14), .Y(n1) );
  INVX1 U48 ( .A(n1), .Y(n2) );
  AND2X2 U51 ( .A(\addr<1> ), .B(\busy<1> ), .Y(n3) );
  INVX1 U54 ( .A(n3), .Y(n4) );
  AND2X2 U57 ( .A(\addr<1> ), .B(\busy<3> ), .Y(n5) );
  INVX1 U60 ( .A(n5), .Y(n6) );
  OR2X2 U63 ( .A(n60), .B(n61), .Y(n7) );
  INVX1 U66 ( .A(n7), .Y(n8) );
  OR2X2 U69 ( .A(n62), .B(n114), .Y(n12) );
  INVX1 U72 ( .A(n12), .Y(n14) );
  INVX1 U79 ( .A(n15), .Y(n17) );
  AND2X1 U80 ( .A(n113), .B(n114), .Y(n18) );
  INVX1 U81 ( .A(n18), .Y(n19) );
  AND2X1 U82 ( .A(n20), .B(n114), .Y(n21) );
  INVX1 U83 ( .A(n21), .Y(n55) );
  AND2X1 U84 ( .A(n11), .B(n113), .Y(n56) );
  INVX1 U85 ( .A(n56), .Y(n57) );
  AND2X2 U86 ( .A(\addr<2> ), .B(\addr<1> ), .Y(n58) );
  INVX1 U87 ( .A(n58), .Y(n59) );
  INVX1 U88 ( .A(n114), .Y(n60) );
  INVX1 U89 ( .A(n9), .Y(n61) );
  INVX1 U90 ( .A(n10), .Y(n62) );
  AND2X2 U91 ( .A(n52), .B(n53), .Y(n63) );
  INVX1 U92 ( .A(n63), .Y(\data_out<0> ) );
  AND2X2 U93 ( .A(n50), .B(n51), .Y(n65) );
  INVX1 U94 ( .A(n65), .Y(\data_out<10> ) );
  AND2X2 U95 ( .A(n48), .B(n49), .Y(n67) );
  INVX1 U96 ( .A(n67), .Y(\data_out<11> ) );
  AND2X2 U97 ( .A(n46), .B(n47), .Y(n69) );
  INVX1 U98 ( .A(n69), .Y(\data_out<12> ) );
  AND2X2 U99 ( .A(n44), .B(n45), .Y(n71) );
  INVX1 U100 ( .A(n71), .Y(\data_out<13> ) );
  AND2X2 U101 ( .A(n42), .B(n43), .Y(n73) );
  INVX1 U102 ( .A(n73), .Y(\data_out<14> ) );
  AND2X2 U103 ( .A(n40), .B(n41), .Y(n75) );
  INVX1 U104 ( .A(n75), .Y(\data_out<15> ) );
  AND2X2 U105 ( .A(n38), .B(n39), .Y(n77) );
  INVX1 U106 ( .A(n77), .Y(\data_out<1> ) );
  AND2X2 U107 ( .A(n36), .B(n37), .Y(n79) );
  INVX1 U108 ( .A(n79), .Y(\data_out<2> ) );
  AND2X2 U109 ( .A(n34), .B(n35), .Y(n81) );
  INVX1 U110 ( .A(n81), .Y(\data_out<3> ) );
  AND2X2 U111 ( .A(n32), .B(n33), .Y(n83) );
  INVX1 U112 ( .A(n83), .Y(\data_out<4> ) );
  AND2X2 U113 ( .A(n30), .B(n31), .Y(n85) );
  INVX1 U114 ( .A(n85), .Y(\data_out<5> ) );
  AND2X2 U115 ( .A(n28), .B(n29), .Y(n87) );
  INVX1 U116 ( .A(n87), .Y(\data_out<6> ) );
  AND2X2 U117 ( .A(n26), .B(n27), .Y(n89) );
  INVX1 U118 ( .A(n89), .Y(\data_out<7> ) );
  AND2X2 U119 ( .A(n24), .B(n25), .Y(n91) );
  INVX1 U120 ( .A(n91), .Y(\data_out<8> ) );
  AND2X2 U121 ( .A(n22), .B(n23), .Y(n93) );
  INVX1 U122 ( .A(n93), .Y(\data_out<9> ) );
  INVX1 U123 ( .A(n95), .Y(n96) );
  INVX1 U124 ( .A(\addr<4> ), .Y(n100) );
  INVX1 U125 ( .A(\addr<1> ), .Y(n113) );
  INVX1 U126 ( .A(\addr<3> ), .Y(n98) );
endmodule


module dff_266 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_265 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_264 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_263 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_245 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_246 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_247 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_248 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_249 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_250 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_251 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_252 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_253 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_254 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_255 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_256 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_257 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_258 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_259 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_260 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_262 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_229 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_230 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_231 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_232 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_233 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_234 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_235 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_236 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_237 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_238 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_239 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_240 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_241 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_242 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_243 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_244 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_261 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_224 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_225 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_226 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_227 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_228 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_221 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_222 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_223 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_216 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_217 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_218 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_219 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_220 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module mem_system ( .DataOut({\DataOut<15> , \DataOut<14> , \DataOut<13> , 
        \DataOut<12> , \DataOut<11> , \DataOut<10> , \DataOut<9> , 
        \DataOut<8> , \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , 
        \DataOut<3> , \DataOut<2> , \DataOut<1> , \DataOut<0> }), Done, Stall, 
        CacheHit, err, .Addr({\Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , 
        \Addr<11> , \Addr<10> , \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , 
        \Addr<5> , \Addr<4> , \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> }), 
    .DataIn({\DataIn<15> , \DataIn<14> , \DataIn<13> , \DataIn<12> , 
        \DataIn<11> , \DataIn<10> , \DataIn<9> , \DataIn<8> , \DataIn<7> , 
        \DataIn<6> , \DataIn<5> , \DataIn<4> , \DataIn<3> , \DataIn<2> , 
        \DataIn<1> , \DataIn<0> }), Rd, Wr, createdump, clk, rst );
  input \Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , \Addr<11> , \Addr<10> ,
         \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , \Addr<5> , \Addr<4> ,
         \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> , \DataIn<15> ,
         \DataIn<14> , \DataIn<13> , \DataIn<12> , \DataIn<11> , \DataIn<10> ,
         \DataIn<9> , \DataIn<8> , \DataIn<7> , \DataIn<6> , \DataIn<5> ,
         \DataIn<4> , \DataIn<3> , \DataIn<2> , \DataIn<1> , \DataIn<0> , Rd,
         Wr, createdump, clk, rst;
  output \DataOut<15> , \DataOut<14> , \DataOut<13> , \DataOut<12> ,
         \DataOut<11> , \DataOut<10> , \DataOut<9> , \DataOut<8> ,
         \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , \DataOut<3> ,
         \DataOut<2> , \DataOut<1> , \DataOut<0> , Done, Stall, CacheHit, err;
  wire   \tagOut0<4> , \tagOut0<3> , \tagOut0<2> , \tagOut0<1> , \tagOut0<0> ,
         \cacheDataOut0<15> , \cacheDataOut0<14> , \cacheDataOut0<13> ,
         \cacheDataOut0<12> , \cacheDataOut0<11> , \cacheDataOut0<10> ,
         \cacheDataOut0<9> , \cacheDataOut0<8> , \cacheDataOut0<7> ,
         \cacheDataOut0<6> , \cacheDataOut0<5> , \cacheDataOut0<4> ,
         \cacheDataOut0<3> , \cacheDataOut0<2> , \cacheDataOut0<1> ,
         \cacheDataOut0<0> , cacheHit0, dirty0, valid0, \cacheOff<2> ,
         \cacheOff<0> , \cacheDataIn<15> , \cacheDataIn<14> ,
         \cacheDataIn<13> , \cacheDataIn<12> , \cacheDataIn<11> ,
         \cacheDataIn<10> , \cacheDataIn<9> , \cacheDataIn<8> ,
         \cacheDataIn<7> , \cacheDataIn<6> , \cacheDataIn<5> ,
         \cacheDataIn<4> , \cacheDataIn<3> , \cacheDataIn<2> ,
         \cacheDataIn<1> , \cacheDataIn<0> , cacheComp, cacheWr,
         \cacheDataOut1<15> , \cacheDataOut1<14> , \cacheDataOut1<13> ,
         \cacheDataOut1<12> , \cacheDataOut1<11> , \cacheDataOut1<10> ,
         \cacheDataOut1<9> , \cacheDataOut1<8> , \cacheDataOut1<7> ,
         \cacheDataOut1<6> , \cacheDataOut1<5> , \cacheDataOut1<4> ,
         \cacheDataOut1<3> , \cacheDataOut1<2> , \cacheDataOut1<1> ,
         \cacheDataOut1<0> , cacheHit1, dirty1, valid1, memAddr_0,
         \memDataIn<15> , \memDataIn<14> , \memDataIn<13> , \memDataIn<12> ,
         \memDataIn<11> , \memDataIn<10> , \memDataIn<9> , \memDataIn<8> ,
         \memDataIn<7> , \memDataIn<6> , \memDataIn<5> , \memDataIn<4> ,
         \memDataIn<3> , \memDataIn<2> , \memDataIn<1> , \memDataIn<0> , memWr,
         \memDataOut<15> , \memDataOut<14> , \memDataOut<13> ,
         \memDataOut<12> , \memDataOut<11> , \memDataOut<10> , \memDataOut<9> ,
         \memDataOut<8> , \memDataOut<7> , \memDataOut<6> , \memDataOut<5> ,
         \memDataOut<4> , \memDataOut<3> , \memDataOut<2> , \memDataOut<1> ,
         \memDataOut<0> , memStall, victimWay, victimWay_in, victimWrite,
         victimWrite_in, stallWait_in, doneWait_in, \memDataOut_flop<15> ,
         \memDataOut_flop<14> , \memDataOut_flop<13> , \memDataOut_flop<12> ,
         \memDataOut_flop<11> , \memDataOut_flop<10> , \memDataOut_flop<9> ,
         \memDataOut_flop<8> , \memDataOut_flop<7> , \memDataOut_flop<6> ,
         \memDataOut_flop<5> , \memDataOut_flop<4> , \memDataOut_flop<3> ,
         \memDataOut_flop<2> , \memDataOut_flop<1> , \memDataOut_flop<0> ,
         waitMem_flop, \cacheDataOut_flop<15> , \cacheDataOut_flop<14> ,
         \cacheDataOut_flop<13> , \cacheDataOut_flop<12> ,
         \cacheDataOut_flop<11> , \cacheDataOut_flop<10> ,
         \cacheDataOut_flop<9> , \cacheDataOut_flop<8> ,
         \cacheDataOut_flop<7> , \cacheDataOut_flop<6> ,
         \cacheDataOut_flop<5> , \cacheDataOut_flop<4> ,
         \cacheDataOut_flop<3> , \cacheDataOut_flop<2> ,
         \cacheDataOut_flop<1> , \cacheDataOut_flop<0> , waitCacheHit_in,
         \nxtState<4> , \nxtState<3> , \nxtState<2> , \nxtState<1> ,
         \nxtState<0> , \state<4> , \state<3> , \state<2> , \state<1> ,
         \state<0> , \wait4Cycles_flop<0> , \wait4Cycles_in<2> ,
         \wait4Cycles_in<1> , \wait4Cycles_in<0> , \nextEvictState_in<4> ,
         \nxtEvict<4> , \nxtEvict<3> , \nxtEvict<2> , \nxtEvict<1> ,
         \nxtEvict<0> , n6, n9, n11, n265, n276, n277, n291, n293, n296, n297,
         n304, n307, n308, n309, n310, n335, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941;

  XOR2X1 U8 ( .A(n396), .B(n715), .Y(n6) );
  MUX2X1 U27 ( .B(n908), .A(n941), .S(n9), .Y(\cacheDataIn<0> ) );
  MUX2X1 U30 ( .B(n909), .A(n940), .S(n11), .Y(\cacheDataIn<1> ) );
  MUX2X1 U32 ( .B(n910), .A(n939), .S(n733), .Y(\cacheDataIn<2> ) );
  MUX2X1 U33 ( .B(n911), .A(n938), .S(n733), .Y(\cacheDataIn<3> ) );
  MUX2X1 U34 ( .B(n912), .A(n937), .S(n733), .Y(\cacheDataIn<4> ) );
  MUX2X1 U35 ( .B(n913), .A(n936), .S(n733), .Y(\cacheDataIn<5> ) );
  MUX2X1 U36 ( .B(n914), .A(n935), .S(n733), .Y(\cacheDataIn<6> ) );
  MUX2X1 U37 ( .B(n915), .A(n934), .S(n733), .Y(\cacheDataIn<7> ) );
  MUX2X1 U38 ( .B(n916), .A(n933), .S(n733), .Y(\cacheDataIn<8> ) );
  MUX2X1 U39 ( .B(n917), .A(n932), .S(n734), .Y(\cacheDataIn<9> ) );
  MUX2X1 U40 ( .B(n918), .A(n931), .S(n734), .Y(\cacheDataIn<10> ) );
  MUX2X1 U41 ( .B(n919), .A(n930), .S(n734), .Y(\cacheDataIn<11> ) );
  MUX2X1 U42 ( .B(n920), .A(n929), .S(n734), .Y(\cacheDataIn<12> ) );
  MUX2X1 U43 ( .B(n921), .A(n928), .S(n734), .Y(\cacheDataIn<13> ) );
  MUX2X1 U44 ( .B(n922), .A(n927), .S(n734), .Y(\cacheDataIn<14> ) );
  MUX2X1 U45 ( .B(n923), .A(n926), .S(n734), .Y(\cacheDataIn<15> ) );
  AND2X2 U148 ( .A(\Addr<0> ), .B(n685), .Y(memAddr_0) );
  AND2X2 U156 ( .A(\Addr<0> ), .B(n683), .Y(\cacheOff<0> ) );
  XNOR2X1 U255 ( .A(victimWay), .B(n661), .Y(victimWay_in) );
  NAND3X1 U300 ( .A(n699), .B(n924), .C(\Addr<1> ), .Y(n265) );
  NAND3X1 U309 ( .A(n699), .B(n925), .C(\Addr<2> ), .Y(n277) );
  AOI21X1 U327 ( .A(\Addr<2> ), .B(n685), .C(n866), .Y(n291) );
  AOI21X1 U329 ( .A(\Addr<1> ), .B(n685), .C(n675), .Y(n297) );
  AOI22X1 U334 ( .A(\Addr<15> ), .B(n566), .C(\tagOut0<4> ), .D(n582), .Y(n304) );
  AOI22X1 U335 ( .A(n730), .B(n566), .C(\tagOut0<3> ), .D(n582), .Y(n307) );
  AOI22X1 U336 ( .A(n729), .B(n566), .C(\tagOut0<2> ), .D(n582), .Y(n308) );
  AOI22X1 U337 ( .A(n728), .B(n566), .C(\tagOut0<1> ), .D(n582), .Y(n309) );
  AOI22X1 U338 ( .A(n727), .B(n566), .C(\tagOut0<0> ), .D(n582), .Y(n310) );
  AOI22X1 U432 ( .A(waitMem_flop), .B(\cacheDataOut_flop<9> ), .C(
        \memDataOut_flop<9> ), .D(n906), .Y(n368) );
  AOI22X1 U433 ( .A(\cacheDataOut_flop<8> ), .B(waitMem_flop), .C(
        \memDataOut_flop<8> ), .D(n906), .Y(n369) );
  AOI22X1 U434 ( .A(\cacheDataOut_flop<7> ), .B(waitMem_flop), .C(
        \memDataOut_flop<7> ), .D(n906), .Y(n370) );
  AOI22X1 U435 ( .A(\cacheDataOut_flop<6> ), .B(waitMem_flop), .C(
        \memDataOut_flop<6> ), .D(n906), .Y(n371) );
  AOI22X1 U436 ( .A(\cacheDataOut_flop<5> ), .B(waitMem_flop), .C(
        \memDataOut_flop<5> ), .D(n906), .Y(n372) );
  AOI22X1 U437 ( .A(\cacheDataOut_flop<4> ), .B(waitMem_flop), .C(
        \memDataOut_flop<4> ), .D(n906), .Y(n373) );
  AOI22X1 U438 ( .A(\cacheDataOut_flop<3> ), .B(waitMem_flop), .C(
        \memDataOut_flop<3> ), .D(n906), .Y(n374) );
  AOI22X1 U439 ( .A(\cacheDataOut_flop<2> ), .B(waitMem_flop), .C(
        \memDataOut_flop<2> ), .D(n906), .Y(n375) );
  AOI22X1 U440 ( .A(\cacheDataOut_flop<1> ), .B(waitMem_flop), .C(
        \memDataOut_flop<1> ), .D(n906), .Y(n376) );
  AOI22X1 U441 ( .A(\cacheDataOut_flop<15> ), .B(waitMem_flop), .C(
        \memDataOut_flop<15> ), .D(n906), .Y(n377) );
  AOI22X1 U442 ( .A(\cacheDataOut_flop<14> ), .B(waitMem_flop), .C(
        \memDataOut_flop<14> ), .D(n906), .Y(n378) );
  AOI22X1 U443 ( .A(\cacheDataOut_flop<13> ), .B(waitMem_flop), .C(
        \memDataOut_flop<13> ), .D(n906), .Y(n379) );
  AOI22X1 U444 ( .A(\cacheDataOut_flop<12> ), .B(waitMem_flop), .C(
        \memDataOut_flop<12> ), .D(n906), .Y(n380) );
  AOI22X1 U445 ( .A(\cacheDataOut_flop<11> ), .B(waitMem_flop), .C(
        \memDataOut_flop<11> ), .D(n906), .Y(n381) );
  AOI22X1 U446 ( .A(\cacheDataOut_flop<10> ), .B(waitMem_flop), .C(
        \memDataOut_flop<10> ), .D(n906), .Y(n382) );
  AOI22X1 U447 ( .A(\cacheDataOut_flop<0> ), .B(waitMem_flop), .C(
        \memDataOut_flop<0> ), .D(n906), .Y(n383) );
  cache_cache_id0 c0 ( .enable(n438), .clk(clk), .rst(n731), .createdump(
        createdump), .tag_in({\Addr<15> , n730, n729, n728, n727}), .index({
        n750, n748, n746, n744, n742, n740, n738, n736}), .offset({n506, n704, 
        \cacheOff<0> }), .data_in({\cacheDataIn<15> , \cacheDataIn<14> , 
        \cacheDataIn<13> , \cacheDataIn<12> , \cacheDataIn<11> , 
        \cacheDataIn<10> , \cacheDataIn<9> , \cacheDataIn<8> , 
        \cacheDataIn<7> , \cacheDataIn<6> , \cacheDataIn<5> , \cacheDataIn<4> , 
        \cacheDataIn<3> , \cacheDataIn<2> , \cacheDataIn<1> , \cacheDataIn<0> }), .comp(cacheComp), .write(cacheWr), .valid_in(n688), .tag_out({\tagOut0<4> , 
        \tagOut0<3> , \tagOut0<2> , \tagOut0<1> , \tagOut0<0> }), .data_out({
        \cacheDataOut0<15> , \cacheDataOut0<14> , \cacheDataOut0<13> , 
        \cacheDataOut0<12> , \cacheDataOut0<11> , \cacheDataOut0<10> , 
        \cacheDataOut0<9> , \cacheDataOut0<8> , \cacheDataOut0<7> , 
        \cacheDataOut0<6> , \cacheDataOut0<5> , \cacheDataOut0<4> , 
        \cacheDataOut0<3> , \cacheDataOut0<2> , \cacheDataOut0<1> , 
        \cacheDataOut0<0> }), .hit(cacheHit0), .dirty(dirty0), .valid(valid0), 
        .err() );
  cache_cache_id2 c1 ( .enable(n391), .clk(clk), .rst(n731), .createdump(
        createdump), .tag_in({\Addr<15> , n730, n729, n728, n727}), .index({
        n750, n748, n746, n744, n742, n740, n738, n736}), .offset({n506, n704, 
        \cacheOff<0> }), .data_in({\cacheDataIn<15> , \cacheDataIn<14> , 
        \cacheDataIn<13> , \cacheDataIn<12> , \cacheDataIn<11> , 
        \cacheDataIn<10> , \cacheDataIn<9> , \cacheDataIn<8> , 
        \cacheDataIn<7> , \cacheDataIn<6> , \cacheDataIn<5> , \cacheDataIn<4> , 
        \cacheDataIn<3> , \cacheDataIn<2> , \cacheDataIn<1> , \cacheDataIn<0> }), .comp(cacheComp), .write(n407), .valid_in(n688), .tag_out(), .data_out({
        \cacheDataOut1<15> , \cacheDataOut1<14> , \cacheDataOut1<13> , 
        \cacheDataOut1<12> , \cacheDataOut1<11> , \cacheDataOut1<10> , 
        \cacheDataOut1<9> , \cacheDataOut1<8> , \cacheDataOut1<7> , 
        \cacheDataOut1<6> , \cacheDataOut1<5> , \cacheDataOut1<4> , 
        \cacheDataOut1<3> , \cacheDataOut1<2> , \cacheDataOut1<1> , 
        \cacheDataOut1<0> }), .hit(cacheHit1), .dirty(dirty1), .valid(valid1), 
        .err() );
  four_bank_mem fmem ( .clk(clk), .rst(n732), .createdump(createdump), .addr({
        n889, n888, n887, n886, n885, n750, n748, n746, n744, n742, n740, n738, 
        n736, n450, n452, memAddr_0}), .data_in({\memDataIn<15> , 
        \memDataIn<14> , \memDataIn<13> , \memDataIn<12> , \memDataIn<11> , 
        \memDataIn<10> , \memDataIn<9> , \memDataIn<8> , \memDataIn<7> , 
        \memDataIn<6> , \memDataIn<5> , \memDataIn<4> , \memDataIn<3> , 
        \memDataIn<2> , \memDataIn<1> , \memDataIn<0> }), .wr(memWr), .rd(n707), .data_out({\memDataOut<15> , \memDataOut<14> , \memDataOut<13> , 
        \memDataOut<12> , \memDataOut<11> , \memDataOut<10> , \memDataOut<9> , 
        \memDataOut<8> , \memDataOut<7> , \memDataOut<6> , \memDataOut<5> , 
        \memDataOut<4> , \memDataOut<3> , \memDataOut<2> , \memDataOut<1> , 
        \memDataOut<0> }), .stall(memStall), .busy(), .err() );
  dff_266 ff6 ( .q(victimWay), .d(victimWay_in), .clk(clk), .rst(n732) );
  dff_265 ff7 ( .q(victimWrite), .d(victimWrite_in), .clk(clk), .rst(n732) );
  dff_264 waitStall ( .q(Stall), .d(n554), .clk(clk), .rst(n731) );
  dff_263 waitDone ( .q(Done), .d(n552), .clk(clk), .rst(n732) );
  dff_245 \memDataOutWait[0]  ( .q(\memDataOut_flop<0> ), .d(\memDataOut<0> ), 
        .clk(clk), .rst(n732) );
  dff_246 \memDataOutWait[1]  ( .q(\memDataOut_flop<1> ), .d(\memDataOut<1> ), 
        .clk(clk), .rst(n732) );
  dff_247 \memDataOutWait[2]  ( .q(\memDataOut_flop<2> ), .d(\memDataOut<2> ), 
        .clk(clk), .rst(n732) );
  dff_248 \memDataOutWait[3]  ( .q(\memDataOut_flop<3> ), .d(\memDataOut<3> ), 
        .clk(clk), .rst(n732) );
  dff_249 \memDataOutWait[4]  ( .q(\memDataOut_flop<4> ), .d(\memDataOut<4> ), 
        .clk(clk), .rst(n731) );
  dff_250 \memDataOutWait[5]  ( .q(\memDataOut_flop<5> ), .d(\memDataOut<5> ), 
        .clk(clk), .rst(n732) );
  dff_251 \memDataOutWait[6]  ( .q(\memDataOut_flop<6> ), .d(\memDataOut<6> ), 
        .clk(clk), .rst(n732) );
  dff_252 \memDataOutWait[7]  ( .q(\memDataOut_flop<7> ), .d(\memDataOut<7> ), 
        .clk(clk), .rst(n732) );
  dff_253 \memDataOutWait[8]  ( .q(\memDataOut_flop<8> ), .d(\memDataOut<8> ), 
        .clk(clk), .rst(n732) );
  dff_254 \memDataOutWait[9]  ( .q(\memDataOut_flop<9> ), .d(\memDataOut<9> ), 
        .clk(clk), .rst(n731) );
  dff_255 \memDataOutWait[10]  ( .q(\memDataOut_flop<10> ), .d(
        \memDataOut<10> ), .clk(clk), .rst(n731) );
  dff_256 \memDataOutWait[11]  ( .q(\memDataOut_flop<11> ), .d(
        \memDataOut<11> ), .clk(clk), .rst(n732) );
  dff_257 \memDataOutWait[12]  ( .q(\memDataOut_flop<12> ), .d(
        \memDataOut<12> ), .clk(clk), .rst(n732) );
  dff_258 \memDataOutWait[13]  ( .q(\memDataOut_flop<13> ), .d(
        \memDataOut<13> ), .clk(clk), .rst(n732) );
  dff_259 \memDataOutWait[14]  ( .q(\memDataOut_flop<14> ), .d(
        \memDataOut<14> ), .clk(clk), .rst(n732) );
  dff_260 \memDataOutWait[15]  ( .q(\memDataOut_flop<15> ), .d(
        \memDataOut<15> ), .clk(clk), .rst(n731) );
  dff_262 waitMem ( .q(waitMem_flop), .d(n520), .clk(clk), .rst(n732) );
  dff_229 \cacheDataOutWait[0]  ( .q(\cacheDataOut_flop<0> ), .d(n869), .clk(
        clk), .rst(n732) );
  dff_230 \cacheDataOutWait[1]  ( .q(\cacheDataOut_flop<1> ), .d(n870), .clk(
        clk), .rst(n731) );
  dff_231 \cacheDataOutWait[2]  ( .q(\cacheDataOut_flop<2> ), .d(n871), .clk(
        clk), .rst(n732) );
  dff_232 \cacheDataOutWait[3]  ( .q(\cacheDataOut_flop<3> ), .d(n872), .clk(
        clk), .rst(n731) );
  dff_233 \cacheDataOutWait[4]  ( .q(\cacheDataOut_flop<4> ), .d(n873), .clk(
        clk), .rst(n732) );
  dff_234 \cacheDataOutWait[5]  ( .q(\cacheDataOut_flop<5> ), .d(n874), .clk(
        clk), .rst(n732) );
  dff_235 \cacheDataOutWait[6]  ( .q(\cacheDataOut_flop<6> ), .d(n875), .clk(
        clk), .rst(n732) );
  dff_236 \cacheDataOutWait[7]  ( .q(\cacheDataOut_flop<7> ), .d(n876), .clk(
        clk), .rst(n732) );
  dff_237 \cacheDataOutWait[8]  ( .q(\cacheDataOut_flop<8> ), .d(n877), .clk(
        clk), .rst(n732) );
  dff_238 \cacheDataOutWait[9]  ( .q(\cacheDataOut_flop<9> ), .d(n878), .clk(
        clk), .rst(n731) );
  dff_239 \cacheDataOutWait[10]  ( .q(\cacheDataOut_flop<10> ), .d(n879), 
        .clk(clk), .rst(n732) );
  dff_240 \cacheDataOutWait[11]  ( .q(\cacheDataOut_flop<11> ), .d(n880), 
        .clk(clk), .rst(n732) );
  dff_241 \cacheDataOutWait[12]  ( .q(\cacheDataOut_flop<12> ), .d(n881), 
        .clk(clk), .rst(n731) );
  dff_242 \cacheDataOutWait[13]  ( .q(\cacheDataOut_flop<13> ), .d(n882), 
        .clk(clk), .rst(n732) );
  dff_243 \cacheDataOutWait[14]  ( .q(\cacheDataOut_flop<14> ), .d(n883), 
        .clk(clk), .rst(n732) );
  dff_244 \cacheDataOutWait[15]  ( .q(\cacheDataOut_flop<15> ), .d(n884), 
        .clk(clk), .rst(n731) );
  dff_261 WaitCacheHit_in ( .q(CacheHit), .d(waitCacheHit_in), .clk(clk), 
        .rst(n731) );
  dff_224 \stateReg[0]  ( .q(\state<0> ), .d(\nxtState<0> ), .clk(clk), .rst(
        n732) );
  dff_225 \stateReg[1]  ( .q(\state<1> ), .d(n550), .clk(clk), .rst(n732) );
  dff_226 \stateReg[2]  ( .q(\state<2> ), .d(\nxtState<2> ), .clk(clk), .rst(
        n731) );
  dff_227 \stateReg[3]  ( .q(\state<3> ), .d(\nxtState<3> ), .clk(clk), .rst(
        n732) );
  dff_228 \stateReg[4]  ( .q(\state<4> ), .d(n548), .clk(clk), .rst(n732) );
  dff_221 \wait4CycleFlop[0]  ( .q(\wait4Cycles_flop<0> ), .d(
        \wait4Cycles_in<0> ), .clk(clk), .rst(n731) );
  dff_222 \wait4CycleFlop[1]  ( .q(\wait4Cycles_in<0> ), .d(
        \wait4Cycles_in<1> ), .clk(clk), .rst(n731) );
  dff_223 \wait4CycleFlop[2]  ( .q(\wait4Cycles_in<1> ), .d(
        \wait4Cycles_in<2> ), .clk(clk), .rst(n732) );
  dff_216 \evictWait[0]  ( .q(\nxtEvict<0> ), .d(n569), .clk(clk), .rst(n732)
         );
  dff_217 \evictWait[1]  ( .q(\nxtEvict<1> ), .d(n567), .clk(clk), .rst(n732)
         );
  dff_218 \evictWait[2]  ( .q(\nxtEvict<2> ), .d(n665), .clk(clk), .rst(n732)
         );
  dff_219 \evictWait[3]  ( .q(\nxtEvict<3> ), .d(n663), .clk(clk), .rst(n731)
         );
  dff_220 \evictWait[4]  ( .q(\nxtEvict<4> ), .d(n687), .clk(clk), .rst(n731)
         );
  AND2X2 U448 ( .A(n524), .B(n458), .Y(n692) );
  INVX2 U449 ( .A(n702), .Y(n703) );
  AND2X2 U450 ( .A(n530), .B(n816), .Y(n702) );
  INVX2 U451 ( .A(n694), .Y(n695) );
  AND2X2 U452 ( .A(n816), .B(n542), .Y(n694) );
  AND2X2 U453 ( .A(n561), .B(n530), .Y(n696) );
  INVX2 U454 ( .A(n752), .Y(n867) );
  AND2X2 U455 ( .A(n691), .B(n697), .Y(n586) );
  AND2X2 U456 ( .A(n524), .B(n857), .Y(n690) );
  OR2X2 U457 ( .A(n403), .B(n516), .Y(n384) );
  INVX8 U458 ( .A(n705), .Y(n704) );
  AND2X2 U459 ( .A(n725), .B(n797), .Y(n677) );
  INVX1 U460 ( .A(n507), .Y(n385) );
  INVX1 U461 ( .A(n507), .Y(n508) );
  AND2X2 U462 ( .A(cacheComp), .B(waitCacheHit_in), .Y(n646) );
  INVX2 U463 ( .A(n413), .Y(n396) );
  INVX1 U464 ( .A(n855), .Y(n856) );
  OR2X1 U465 ( .A(n601), .B(n692), .Y(n648) );
  BUFX2 U466 ( .A(n865), .Y(n733) );
  BUFX2 U467 ( .A(n865), .Y(n734) );
  INVX1 U468 ( .A(\DataIn<0> ), .Y(n941) );
  INVX1 U469 ( .A(\DataIn<1> ), .Y(n940) );
  INVX1 U470 ( .A(\DataIn<2> ), .Y(n939) );
  INVX1 U471 ( .A(\DataIn<3> ), .Y(n938) );
  INVX1 U472 ( .A(\DataIn<4> ), .Y(n937) );
  INVX1 U473 ( .A(\DataIn<5> ), .Y(n936) );
  INVX1 U474 ( .A(\DataIn<6> ), .Y(n935) );
  INVX1 U475 ( .A(\DataIn<7> ), .Y(n934) );
  INVX1 U476 ( .A(\DataIn<8> ), .Y(n933) );
  INVX1 U477 ( .A(\DataIn<9> ), .Y(n932) );
  INVX1 U478 ( .A(\DataIn<10> ), .Y(n931) );
  INVX1 U479 ( .A(\DataIn<11> ), .Y(n930) );
  INVX1 U480 ( .A(\DataIn<12> ), .Y(n929) );
  INVX1 U481 ( .A(\DataIn<13> ), .Y(n928) );
  INVX1 U482 ( .A(\DataIn<14> ), .Y(n927) );
  INVX1 U483 ( .A(\DataIn<15> ), .Y(n926) );
  OR2X1 U484 ( .A(Wr), .B(Rd), .Y(n862) );
  INVX1 U485 ( .A(victimWrite), .Y(n841) );
  INVX1 U486 ( .A(\nxtEvict<3> ), .Y(n767) );
  INVX1 U487 ( .A(\nxtEvict<4> ), .Y(n828) );
  OR2X1 U488 ( .A(n533), .B(n386), .Y(n441) );
  INVX1 U489 ( .A(\Addr<2> ), .Y(n924) );
  INVX1 U490 ( .A(\Addr<1> ), .Y(n925) );
  INVX1 U491 ( .A(victimWay), .Y(n724) );
  OR2X1 U492 ( .A(\wait4Cycles_in<1> ), .B(\wait4Cycles_in<0> ), .Y(n773) );
  INVX1 U493 ( .A(Wr), .Y(n765) );
  OR2X1 U494 ( .A(n517), .B(n533), .Y(n446) );
  INVX1 U495 ( .A(\wait4Cycles_in<1> ), .Y(n755) );
  AND2X1 U496 ( .A(n464), .B(n689), .Y(n604) );
  INVX1 U497 ( .A(\memDataOut<7> ), .Y(n915) );
  INVX1 U498 ( .A(\memDataOut<14> ), .Y(n922) );
  INVX1 U499 ( .A(\memDataOut<0> ), .Y(n908) );
  INVX1 U500 ( .A(\memDataOut<1> ), .Y(n909) );
  INVX1 U501 ( .A(\memDataOut<2> ), .Y(n910) );
  INVX1 U502 ( .A(\memDataOut<3> ), .Y(n911) );
  INVX1 U503 ( .A(\memDataOut<4> ), .Y(n912) );
  INVX1 U504 ( .A(\memDataOut<5> ), .Y(n913) );
  INVX1 U505 ( .A(\memDataOut<6> ), .Y(n914) );
  INVX1 U506 ( .A(\memDataOut<8> ), .Y(n916) );
  INVX1 U507 ( .A(\memDataOut<9> ), .Y(n917) );
  INVX1 U508 ( .A(\memDataOut<10> ), .Y(n918) );
  INVX1 U509 ( .A(\memDataOut<11> ), .Y(n919) );
  INVX1 U510 ( .A(\memDataOut<12> ), .Y(n920) );
  INVX1 U511 ( .A(\memDataOut<13> ), .Y(n921) );
  INVX1 U512 ( .A(\memDataOut<15> ), .Y(n923) );
  AND2X1 U513 ( .A(n492), .B(n440), .Y(n671) );
  OR2X1 U514 ( .A(n571), .B(n602), .Y(n621) );
  INVX1 U515 ( .A(\Addr<6> ), .Y(n743) );
  INVX1 U516 ( .A(\Addr<7> ), .Y(n745) );
  INVX1 U517 ( .A(n747), .Y(n746) );
  INVX1 U518 ( .A(\Addr<8> ), .Y(n747) );
  INVX1 U519 ( .A(n749), .Y(n748) );
  INVX1 U520 ( .A(\Addr<9> ), .Y(n749) );
  INVX1 U521 ( .A(n751), .Y(n750) );
  INVX1 U522 ( .A(\Addr<10> ), .Y(n751) );
  BUFX2 U523 ( .A(\Addr<11> ), .Y(n727) );
  BUFX2 U524 ( .A(\Addr<12> ), .Y(n728) );
  BUFX2 U525 ( .A(\Addr<13> ), .Y(n729) );
  BUFX2 U526 ( .A(\Addr<14> ), .Y(n730) );
  OR2X1 U527 ( .A(n420), .B(n517), .Y(n386) );
  OR2X2 U528 ( .A(n526), .B(n838), .Y(n387) );
  INVX1 U529 ( .A(n429), .Y(n420) );
  OR2X1 U530 ( .A(n585), .B(n603), .Y(n673) );
  OR2X2 U531 ( .A(n420), .B(n535), .Y(n388) );
  AND2X1 U532 ( .A(n715), .B(n713), .Y(n389) );
  AND2X1 U533 ( .A(n449), .B(n867), .Y(n453) );
  INVX1 U534 ( .A(rst), .Y(n735) );
  INVX2 U535 ( .A(memStall), .Y(n759) );
  NOR3X1 U536 ( .A(n489), .B(n501), .C(n757), .Y(n390) );
  OR2X2 U537 ( .A(n477), .B(cacheComp), .Y(n391) );
  INVX1 U538 ( .A(n829), .Y(n392) );
  XNOR2X1 U539 ( .A(\state<2> ), .B(\state<1> ), .Y(n834) );
  INVX2 U540 ( .A(\state<4> ), .Y(n839) );
  INVX2 U541 ( .A(\state<3> ), .Y(n527) );
  MUX2X1 U542 ( .B(dirty1), .A(dirty0), .S(n724), .Y(n393) );
  INVX1 U543 ( .A(\cacheDataOut0<0> ), .Y(n394) );
  MUX2X1 U544 ( .B(n801), .A(n844), .S(n723), .Y(n882) );
  MUX2X1 U545 ( .B(n804), .A(n847), .S(n722), .Y(n879) );
  INVX4 U546 ( .A(n814), .Y(n722) );
  MUX2X1 U547 ( .B(n807), .A(n849), .S(n421), .Y(n876) );
  INVX1 U548 ( .A(n814), .Y(n421) );
  NOR3X1 U549 ( .A(n489), .B(n501), .C(n757), .Y(n395) );
  INVX4 U550 ( .A(n759), .Y(n397) );
  AND2X2 U551 ( .A(n434), .B(n399), .Y(n398) );
  INVX1 U552 ( .A(n398), .Y(n861) );
  INVX1 U553 ( .A(\state<4> ), .Y(n399) );
  INVX1 U554 ( .A(n399), .Y(n400) );
  MUX2X1 U555 ( .B(n813), .A(n712), .S(n401), .Y(n870) );
  INVX1 U556 ( .A(n814), .Y(n401) );
  MUX2X1 U557 ( .B(n800), .A(n710), .S(n401), .Y(n883) );
  INVX1 U558 ( .A(n839), .Y(n402) );
  BUFX2 U559 ( .A(n428), .Y(n403) );
  INVX1 U560 ( .A(n833), .Y(n428) );
  INVX1 U561 ( .A(cacheComp), .Y(n404) );
  INVX8 U562 ( .A(n726), .Y(cacheComp) );
  INVX1 U563 ( .A(n512), .Y(n405) );
  INVX1 U564 ( .A(\state<1> ), .Y(n833) );
  BUFX2 U565 ( .A(n454), .Y(n406) );
  OR2X2 U566 ( .A(n483), .B(n822), .Y(n407) );
  INVX1 U567 ( .A(\state<3> ), .Y(n425) );
  INVX1 U568 ( .A(\cacheDataOut0<13> ), .Y(n408) );
  INVX1 U569 ( .A(\cacheDataOut0<12> ), .Y(n409) );
  INVX1 U570 ( .A(\cacheDataOut0<11> ), .Y(n410) );
  INVX1 U571 ( .A(\cacheDataOut0<5> ), .Y(n411) );
  INVX1 U572 ( .A(\cacheDataOut0<2> ), .Y(n412) );
  INVX1 U573 ( .A(\state<2> ), .Y(n413) );
  INVX1 U574 ( .A(n413), .Y(n414) );
  INVX1 U575 ( .A(\cacheDataOut0<14> ), .Y(n415) );
  INVX1 U576 ( .A(\cacheDataOut0<8> ), .Y(n416) );
  INVX1 U577 ( .A(\cacheDataOut0<7> ), .Y(n417) );
  INVX1 U578 ( .A(\cacheDataOut0<15> ), .Y(n418) );
  INVX1 U579 ( .A(\cacheDataOut0<1> ), .Y(n419) );
  INVX1 U580 ( .A(\state<0> ), .Y(n429) );
  MUX2X1 U581 ( .B(n806), .A(n714), .S(n421), .Y(n877) );
  MUX2X1 U582 ( .B(n812), .A(n717), .S(n722), .Y(n871) );
  MUX2X1 U583 ( .B(n815), .A(n854), .S(n723), .Y(n869) );
  INVX4 U584 ( .A(n798), .Y(n814) );
  INVX4 U585 ( .A(n814), .Y(n723) );
  OR2X1 U586 ( .A(n393), .B(n422), .Y(n479) );
  OR2X2 U587 ( .A(n485), .B(n792), .Y(n422) );
  INVX1 U588 ( .A(n863), .Y(n423) );
  BUFX2 U589 ( .A(n863), .Y(n424) );
  XOR2X1 U590 ( .A(n425), .B(\state<4> ), .Y(n863) );
  INVX1 U591 ( .A(\state<3> ), .Y(n829) );
  INVX2 U592 ( .A(n457), .Y(n866) );
  OR2X2 U593 ( .A(n535), .B(n433), .Y(n426) );
  OR2X2 U594 ( .A(n434), .B(n426), .Y(n427) );
  MUX2X1 U595 ( .B(n511), .A(n498), .S(n429), .Y(n835) );
  AND2X2 U596 ( .A(n403), .B(n864), .Y(n430) );
  INVX1 U597 ( .A(n430), .Y(n431) );
  INVX1 U598 ( .A(n430), .Y(n432) );
  INVX1 U599 ( .A(n864), .Y(n433) );
  INVX1 U600 ( .A(\state<0> ), .Y(n434) );
  INVX4 U601 ( .A(n510), .Y(n864) );
  AND2X2 U602 ( .A(n787), .B(n573), .Y(n435) );
  INVX1 U603 ( .A(n435), .Y(n436) );
  AND2X2 U604 ( .A(n837), .B(n726), .Y(n437) );
  INVX1 U605 ( .A(n437), .Y(n438) );
  OR2X2 U606 ( .A(n861), .B(n514), .Y(n439) );
  OR2X1 U607 ( .A(n517), .B(n384), .Y(n440) );
  OR2X2 U608 ( .A(n468), .B(n443), .Y(n442) );
  OR2X2 U609 ( .A(n607), .B(n467), .Y(n443) );
  OR2X2 U610 ( .A(n527), .B(n387), .Y(n444) );
  OR2X2 U611 ( .A(n405), .B(n532), .Y(n445) );
  OR2X2 U612 ( .A(n536), .B(n388), .Y(n447) );
  OR2X2 U613 ( .A(n700), .B(n578), .Y(n448) );
  INVX1 U614 ( .A(n448), .Y(n449) );
  OR2X2 U615 ( .A(n680), .B(n579), .Y(n450) );
  AND2X2 U616 ( .A(n478), .B(n453), .Y(n451) );
  INVX1 U617 ( .A(n451), .Y(n452) );
  AND2X2 U618 ( .A(\state<2> ), .B(n833), .Y(n454) );
  AND2X2 U619 ( .A(n868), .B(n713), .Y(n455) );
  AND2X2 U620 ( .A(n455), .B(n476), .Y(n456) );
  INVX1 U621 ( .A(n456), .Y(n457) );
  AND2X2 U622 ( .A(n760), .B(n405), .Y(n458) );
  AND2X2 U623 ( .A(n530), .B(n458), .Y(n459) );
  INVX1 U624 ( .A(n459), .Y(n460) );
  AND2X2 U625 ( .A(n458), .B(n398), .Y(n461) );
  INVX1 U626 ( .A(n461), .Y(n462) );
  AND2X2 U627 ( .A(n403), .B(n563), .Y(n463) );
  INVX1 U628 ( .A(n463), .Y(n464) );
  AND2X2 U629 ( .A(n868), .B(n528), .Y(n465) );
  AND2X2 U630 ( .A(n527), .B(n862), .Y(n466) );
  AND2X2 U631 ( .A(n405), .B(n539), .Y(n467) );
  OR2X2 U632 ( .A(n835), .B(n465), .Y(n468) );
  AND2X2 U633 ( .A(n838), .B(n866), .Y(n469) );
  OR2X2 U634 ( .A(n713), .B(n403), .Y(n470) );
  INVX1 U635 ( .A(n470), .Y(n471) );
  BUFX2 U636 ( .A(n825), .Y(n472) );
  AND2X2 U637 ( .A(cacheHit1), .B(valid1), .Y(n473) );
  INVX1 U638 ( .A(n473), .Y(n474) );
  OR2X2 U639 ( .A(n400), .B(n512), .Y(n475) );
  INVX1 U640 ( .A(n475), .Y(n476) );
  AND2X2 U641 ( .A(n442), .B(victimWrite), .Y(n477) );
  BUFX2 U642 ( .A(n297), .Y(n478) );
  INVX1 U643 ( .A(n479), .Y(n480) );
  AND2X2 U644 ( .A(n460), .B(n792), .Y(n481) );
  INVX1 U645 ( .A(n481), .Y(n482) );
  BUFX2 U646 ( .A(n821), .Y(n483) );
  AND2X2 U647 ( .A(valid0), .B(n721), .Y(n484) );
  INVX1 U648 ( .A(n484), .Y(n485) );
  BUFX2 U649 ( .A(n762), .Y(n486) );
  BUFX2 U650 ( .A(n827), .Y(n487) );
  INVX1 U651 ( .A(n563), .Y(n488) );
  AND2X2 U652 ( .A(n455), .B(n398), .Y(n563) );
  OR2X2 U653 ( .A(n461), .B(n537), .Y(n489) );
  OR2X2 U654 ( .A(n688), .B(n860), .Y(n490) );
  INVX1 U655 ( .A(n490), .Y(n491) );
  OR2X2 U656 ( .A(n534), .B(n446), .Y(n492) );
  OR2X2 U657 ( .A(n420), .B(n403), .Y(n493) );
  INVX1 U658 ( .A(n493), .Y(n494) );
  AND2X2 U659 ( .A(n713), .B(n528), .Y(n495) );
  INVX1 U660 ( .A(n495), .Y(n496) );
  AND2X2 U661 ( .A(n834), .B(n423), .Y(n497) );
  INVX1 U662 ( .A(n497), .Y(n498) );
  AND2X2 U663 ( .A(\nxtEvict<4> ), .B(n537), .Y(n499) );
  INVX1 U664 ( .A(n499), .Y(n500) );
  OR2X2 U665 ( .A(n519), .B(n389), .Y(n501) );
  AND2X2 U666 ( .A(\nxtEvict<0> ), .B(n793), .Y(n502) );
  INVX1 U667 ( .A(n502), .Y(n503) );
  AND2X2 U668 ( .A(n772), .B(n771), .Y(n504) );
  INVX1 U669 ( .A(n504), .Y(n505) );
  BUFX2 U670 ( .A(\cacheOff<2> ), .Y(n506) );
  AND2X2 U671 ( .A(n458), .B(n542), .Y(n507) );
  AND2X2 U672 ( .A(n414), .B(n829), .Y(n509) );
  INVX1 U673 ( .A(n509), .Y(n510) );
  INVX1 U674 ( .A(n509), .Y(n511) );
  INVX1 U675 ( .A(n833), .Y(n512) );
  INVX1 U676 ( .A(n529), .Y(n513) );
  NOR2X1 U677 ( .A(n428), .B(n513), .Y(n515) );
  INVX1 U678 ( .A(n515), .Y(n514) );
  INVX1 U679 ( .A(n542), .Y(n516) );
  INVX1 U680 ( .A(n529), .Y(n517) );
  AND2X2 U681 ( .A(n508), .B(n444), .Y(n518) );
  INVX1 U682 ( .A(n518), .Y(n519) );
  INVX1 U683 ( .A(n518), .Y(n520) );
  AND2X2 U684 ( .A(cacheHit0), .B(valid0), .Y(n521) );
  INVX1 U685 ( .A(n521), .Y(n522) );
  INVX1 U686 ( .A(n458), .Y(n523) );
  AND2X2 U687 ( .A(n402), .B(n838), .Y(n524) );
  INVX1 U688 ( .A(n524), .Y(n525) );
  INVX1 U689 ( .A(n465), .Y(n526) );
  AND2X2 U690 ( .A(n428), .B(n839), .Y(n528) );
  AND2X2 U691 ( .A(n396), .B(n392), .Y(n529) );
  AND2X2 U692 ( .A(n400), .B(\state<0> ), .Y(n530) );
  INVX1 U693 ( .A(n530), .Y(n531) );
  INVX1 U694 ( .A(n760), .Y(n532) );
  INVX1 U695 ( .A(n414), .Y(n868) );
  INVX1 U696 ( .A(n528), .Y(n533) );
  INVX1 U697 ( .A(n420), .Y(n534) );
  INVX1 U698 ( .A(n528), .Y(n535) );
  INVX1 U699 ( .A(n864), .Y(n536) );
  INVX4 U700 ( .A(\state<0> ), .Y(n838) );
  AND2X2 U701 ( .A(n524), .B(n816), .Y(n537) );
  AND2X2 U702 ( .A(n420), .B(n866), .Y(n538) );
  AND2X2 U703 ( .A(n396), .B(n839), .Y(n539) );
  AND2X2 U704 ( .A(n420), .B(n403), .Y(n540) );
  BUFX2 U705 ( .A(n763), .Y(n541) );
  INVX1 U706 ( .A(n541), .Y(n542) );
  INVX1 U707 ( .A(n541), .Y(n543) );
  AND2X2 U708 ( .A(n402), .B(n864), .Y(n544) );
  INVX1 U709 ( .A(n544), .Y(n545) );
  INVX1 U710 ( .A(n455), .Y(n546) );
  INVX1 U711 ( .A(\nxtState<4> ), .Y(n547) );
  INVX1 U712 ( .A(n547), .Y(n548) );
  INVX1 U713 ( .A(\nxtState<1> ), .Y(n549) );
  INVX1 U714 ( .A(n549), .Y(n550) );
  INVX1 U715 ( .A(doneWait_in), .Y(n551) );
  INVX1 U716 ( .A(n551), .Y(n552) );
  INVX1 U717 ( .A(stallWait_in), .Y(n553) );
  INVX1 U718 ( .A(n553), .Y(n554) );
  INVX1 U719 ( .A(n858), .Y(n555) );
  INVX1 U720 ( .A(n555), .Y(n556) );
  OR2X2 U721 ( .A(n480), .B(n584), .Y(n557) );
  INVX1 U722 ( .A(n557), .Y(n558) );
  AND2X2 U723 ( .A(n770), .B(n677), .Y(n559) );
  INVX1 U724 ( .A(n559), .Y(n560) );
  AND2X2 U725 ( .A(n527), .B(n406), .Y(n561) );
  INVX1 U726 ( .A(n561), .Y(n562) );
  INVX1 U727 ( .A(n563), .Y(n564) );
  AND2X1 U728 ( .A(n460), .B(n581), .Y(n565) );
  INVX1 U729 ( .A(n565), .Y(n566) );
  OR2X1 U730 ( .A(n754), .B(n568), .Y(n567) );
  OR2X1 U731 ( .A(n538), .B(n587), .Y(n568) );
  OR2X1 U732 ( .A(n752), .B(n570), .Y(n569) );
  OR2X1 U733 ( .A(n469), .B(n754), .Y(n570) );
  OR2X1 U734 ( .A(n597), .B(n572), .Y(n571) );
  OR2X1 U735 ( .A(n643), .B(n632), .Y(n572) );
  AND2X2 U736 ( .A(n464), .B(n447), .Y(n573) );
  OR2X1 U737 ( .A(n663), .B(n575), .Y(n574) );
  OR2X1 U738 ( .A(n625), .B(n626), .Y(n575) );
  OR2X1 U739 ( .A(n864), .B(n577), .Y(n576) );
  OR2X1 U740 ( .A(n466), .B(n528), .Y(n577) );
  OR2X1 U741 ( .A(n667), .B(n538), .Y(n578) );
  OR2X1 U742 ( .A(n679), .B(n587), .Y(n579) );
  INVX1 U743 ( .A(n537), .Y(n580) );
  AND2X1 U744 ( .A(n664), .B(n662), .Y(n581) );
  OR2X1 U745 ( .A(n589), .B(n583), .Y(n582) );
  OR2X1 U746 ( .A(n588), .B(n276), .Y(n583) );
  OR2X1 U747 ( .A(n766), .B(n597), .Y(n584) );
  AND2X1 U748 ( .A(n668), .B(n696), .Y(n585) );
  INVX1 U749 ( .A(n586), .Y(n587) );
  OR2X1 U750 ( .A(n596), .B(n605), .Y(n588) );
  OR2X1 U751 ( .A(n670), .B(n672), .Y(n589) );
  OR2X1 U752 ( .A(n594), .B(n694), .Y(n590) );
  INVX1 U753 ( .A(n590), .Y(n591) );
  BUFX2 U754 ( .A(n775), .Y(n592) );
  AND2X1 U755 ( .A(n693), .B(n720), .Y(n593) );
  INVX1 U756 ( .A(n593), .Y(n594) );
  AND2X1 U757 ( .A(n701), .B(n695), .Y(n595) );
  INVX1 U758 ( .A(n595), .Y(n596) );
  INVX1 U759 ( .A(n440), .Y(n597) );
  AND2X1 U760 ( .A(n691), .B(n703), .Y(n598) );
  INVX1 U761 ( .A(n598), .Y(n599) );
  AND2X2 U762 ( .A(n492), .B(n464), .Y(n600) );
  INVX1 U763 ( .A(n600), .Y(n601) );
  BUFX2 U764 ( .A(n782), .Y(n602) );
  BUFX2 U765 ( .A(n795), .Y(n603) );
  INVX1 U766 ( .A(n604), .Y(n605) );
  BUFX2 U767 ( .A(n794), .Y(n606) );
  INVX1 U768 ( .A(n836), .Y(n607) );
  INVX1 U769 ( .A(n557), .Y(n608) );
  OR2X1 U770 ( .A(n866), .B(n816), .Y(n609) );
  INVX1 U771 ( .A(n609), .Y(n610) );
  INVX1 U772 ( .A(n383), .Y(\DataOut<0> ) );
  INVX1 U773 ( .A(n382), .Y(\DataOut<10> ) );
  INVX1 U774 ( .A(n381), .Y(\DataOut<11> ) );
  INVX1 U775 ( .A(n380), .Y(\DataOut<12> ) );
  INVX1 U776 ( .A(n379), .Y(\DataOut<13> ) );
  INVX1 U777 ( .A(n378), .Y(\DataOut<14> ) );
  INVX1 U778 ( .A(n377), .Y(\DataOut<15> ) );
  INVX1 U779 ( .A(n376), .Y(\DataOut<1> ) );
  INVX1 U780 ( .A(n375), .Y(\DataOut<2> ) );
  INVX1 U781 ( .A(n374), .Y(\DataOut<3> ) );
  INVX1 U782 ( .A(n373), .Y(\DataOut<4> ) );
  INVX1 U783 ( .A(n372), .Y(\DataOut<5> ) );
  INVX1 U784 ( .A(n371), .Y(\DataOut<6> ) );
  INVX1 U785 ( .A(n370), .Y(\DataOut<7> ) );
  INVX1 U786 ( .A(n369), .Y(\DataOut<8> ) );
  INVX1 U787 ( .A(n368), .Y(\DataOut<9> ) );
  INVX1 U788 ( .A(waitMem_flop), .Y(n906) );
  BUFX2 U789 ( .A(n310), .Y(n611) );
  INVX1 U790 ( .A(n611), .Y(n885) );
  BUFX2 U791 ( .A(n309), .Y(n612) );
  INVX1 U792 ( .A(n612), .Y(n886) );
  BUFX2 U793 ( .A(n308), .Y(n613) );
  INVX1 U794 ( .A(n613), .Y(n887) );
  BUFX2 U795 ( .A(n307), .Y(n614) );
  INVX1 U796 ( .A(n614), .Y(n888) );
  INVX1 U797 ( .A(n304), .Y(n889) );
  AND2X2 U798 ( .A(n562), .B(n445), .Y(n615) );
  AND2X1 U799 ( .A(\Addr<2> ), .B(\Addr<1> ), .Y(n616) );
  INVX1 U800 ( .A(n546), .Y(n907) );
  AND2X1 U801 ( .A(n839), .B(n855), .Y(n617) );
  INVX1 U802 ( .A(n617), .Y(n618) );
  AND2X1 U803 ( .A(n676), .B(n715), .Y(n619) );
  INVX1 U804 ( .A(n619), .Y(n620) );
  INVX1 U805 ( .A(n621), .Y(n622) );
  OR2X1 U806 ( .A(n424), .B(n6), .Y(n623) );
  INVX1 U807 ( .A(n623), .Y(n624) );
  INVX1 U808 ( .A(n756), .Y(n625) );
  INVX1 U809 ( .A(n492), .Y(n626) );
  BUFX2 U810 ( .A(n791), .Y(n627) );
  AND2X2 U811 ( .A(n427), .B(n586), .Y(n628) );
  INVX1 U812 ( .A(n628), .Y(n629) );
  AND2X2 U813 ( .A(n864), .B(n533), .Y(n630) );
  INVX1 U814 ( .A(n630), .Y(n631) );
  INVX1 U815 ( .A(n633), .Y(n632) );
  BUFX2 U816 ( .A(n781), .Y(n633) );
  OR2X1 U817 ( .A(\Addr<1> ), .B(\Addr<2> ), .Y(n634) );
  INVX1 U818 ( .A(n634), .Y(n635) );
  AND2X1 U819 ( .A(Rd), .B(n461), .Y(n636) );
  INVX1 U820 ( .A(n636), .Y(n637) );
  AND2X2 U821 ( .A(n471), .B(n817), .Y(n638) );
  INVX1 U822 ( .A(n638), .Y(n639) );
  INVX1 U823 ( .A(n447), .Y(n754) );
  BUFX2 U824 ( .A(n769), .Y(n640) );
  OR2X2 U825 ( .A(n482), .B(n673), .Y(n641) );
  INVX1 U826 ( .A(n641), .Y(n642) );
  AND2X1 U827 ( .A(n669), .B(n696), .Y(n643) );
  OR2X2 U828 ( .A(n599), .B(n436), .Y(n644) );
  INVX1 U829 ( .A(n644), .Y(n645) );
  INVX1 U830 ( .A(n646), .Y(n647) );
  INVX1 U831 ( .A(n648), .Y(n649) );
  AND2X2 U832 ( .A(n693), .B(n492), .Y(n650) );
  INVX1 U833 ( .A(n650), .Y(n651) );
  OR2X2 U834 ( .A(n861), .B(n562), .Y(n652) );
  INVX1 U835 ( .A(n652), .Y(n653) );
  AND2X1 U836 ( .A(n701), .B(n778), .Y(n654) );
  INVX1 U837 ( .A(n654), .Y(n655) );
  OR2X1 U838 ( .A(n715), .B(n540), .Y(n656) );
  INVX1 U839 ( .A(n656), .Y(n657) );
  OR2X1 U840 ( .A(n540), .B(n715), .Y(n658) );
  INVX1 U841 ( .A(n658), .Y(n659) );
  AND2X1 U842 ( .A(n461), .B(n862), .Y(n660) );
  INVX1 U843 ( .A(n660), .Y(n661) );
  AND2X2 U844 ( .A(n457), .B(n427), .Y(n662) );
  INVX1 U845 ( .A(n662), .Y(n663) );
  AND2X2 U846 ( .A(n686), .B(n447), .Y(n664) );
  INVX1 U847 ( .A(n664), .Y(n665) );
  INVX1 U848 ( .A(n448), .Y(n666) );
  INVX1 U849 ( .A(n789), .Y(n667) );
  INVX1 U850 ( .A(n669), .Y(n668) );
  BUFX2 U851 ( .A(n277), .Y(n669) );
  INVX1 U852 ( .A(n395), .Y(n670) );
  INVX1 U853 ( .A(n671), .Y(n672) );
  AND2X2 U854 ( .A(n693), .B(n441), .Y(n674) );
  INVX1 U855 ( .A(n674), .Y(n675) );
  BUFX2 U856 ( .A(n265), .Y(n676) );
  INVX1 U857 ( .A(n677), .Y(n678) );
  INVX1 U858 ( .A(n293), .Y(n679) );
  INVX1 U859 ( .A(n291), .Y(n680) );
  INVX1 U860 ( .A(n335), .Y(n681) );
  INVX1 U861 ( .A(n681), .Y(n682) );
  INVX1 U862 ( .A(n681), .Y(n683) );
  INVX1 U863 ( .A(n296), .Y(n684) );
  INVX1 U864 ( .A(n684), .Y(n685) );
  INVX1 U865 ( .A(n687), .Y(n686) );
  BUFX2 U866 ( .A(\nextEvictState_in<4> ), .Y(n687) );
  AND2X1 U867 ( .A(n857), .B(n530), .Y(n688) );
  INVX1 U868 ( .A(n688), .Y(n689) );
  INVX1 U869 ( .A(n445), .Y(n816) );
  INVX1 U870 ( .A(n580), .Y(n793) );
  INVX1 U871 ( .A(n690), .Y(n691) );
  INVX1 U872 ( .A(n692), .Y(n693) );
  INVX1 U873 ( .A(n696), .Y(n697) );
  OR2X2 U874 ( .A(n774), .B(\Addr<0> ), .Y(n698) );
  INVX1 U875 ( .A(n698), .Y(n699) );
  AND2X1 U876 ( .A(n561), .B(n543), .Y(n700) );
  INVX1 U877 ( .A(n700), .Y(n701) );
  AND2X2 U878 ( .A(n591), .B(n472), .Y(n705) );
  AND2X2 U879 ( .A(n859), .B(n556), .Y(n706) );
  INVX1 U880 ( .A(n706), .Y(n707) );
  INVX1 U881 ( .A(\Addr<5> ), .Y(n741) );
  INVX1 U882 ( .A(n786), .Y(n787) );
  INVX1 U883 ( .A(n786), .Y(n764) );
  MUX2X1 U884 ( .B(n809), .A(n851), .S(n722), .Y(n874) );
  INVX1 U885 ( .A(\cacheDataOut0<3> ), .Y(n708) );
  AND2X2 U886 ( .A(n725), .B(n757), .Y(n709) );
  INVX1 U887 ( .A(n709), .Y(n792) );
  INVX1 U888 ( .A(\cacheDataOut0<14> ), .Y(n710) );
  INVX1 U889 ( .A(\cacheDataOut0<10> ), .Y(n711) );
  INVX1 U890 ( .A(\cacheDataOut0<1> ), .Y(n712) );
  INVX1 U891 ( .A(n527), .Y(n713) );
  INVX1 U892 ( .A(n431), .Y(n857) );
  INVX2 U893 ( .A(\Addr<4> ), .Y(n739) );
  INVX1 U894 ( .A(\cacheDataOut0<8> ), .Y(n714) );
  BUFX2 U895 ( .A(n402), .Y(n715) );
  INVX1 U896 ( .A(\cacheDataOut0<4> ), .Y(n716) );
  INVX1 U897 ( .A(\cacheDataOut0<2> ), .Y(n717) );
  INVX1 U898 ( .A(\cacheDataOut0<6> ), .Y(n718) );
  INVX1 U899 ( .A(\cacheDataOut0<9> ), .Y(n719) );
  BUFX2 U900 ( .A(n564), .Y(n720) );
  INVX1 U901 ( .A(n840), .Y(n721) );
  INVX1 U902 ( .A(valid1), .Y(n840) );
  MUX2X1 U903 ( .B(n805), .A(n848), .S(n723), .Y(n878) );
  MUX2X1 U904 ( .B(n811), .A(n853), .S(n723), .Y(n872) );
  MUX2X1 U905 ( .B(n803), .A(n846), .S(n722), .Y(n880) );
  MUX2X1 U906 ( .B(n802), .A(n845), .S(n722), .Y(n881) );
  MUX2X1 U907 ( .B(n799), .A(n843), .S(n723), .Y(n884) );
  MUX2X1 U908 ( .B(dirty1), .A(dirty0), .S(n724), .Y(n758) );
  INVX1 U909 ( .A(\cacheDataOut1<9> ), .Y(n805) );
  INVX1 U910 ( .A(\cacheDataOut1<15> ), .Y(n799) );
  INVX1 U911 ( .A(\cacheDataOut1<14> ), .Y(n800) );
  INVX1 U912 ( .A(\cacheDataOut1<13> ), .Y(n801) );
  INVX1 U913 ( .A(\cacheDataOut1<12> ), .Y(n802) );
  INVX1 U914 ( .A(\cacheDataOut1<5> ), .Y(n809) );
  INVX1 U915 ( .A(\cacheDataOut0<12> ), .Y(n845) );
  AND2X2 U916 ( .A(n522), .B(n474), .Y(n725) );
  INVX1 U917 ( .A(n725), .Y(waitCacheHit_in) );
  INVX1 U918 ( .A(\cacheDataOut1<11> ), .Y(n803) );
  INVX1 U919 ( .A(\cacheDataOut1<10> ), .Y(n804) );
  INVX1 U920 ( .A(\cacheDataOut1<8> ), .Y(n806) );
  INVX1 U921 ( .A(\cacheDataOut1<7> ), .Y(n807) );
  INVX1 U922 ( .A(\cacheDataOut1<6> ), .Y(n808) );
  INVX1 U923 ( .A(\cacheDataOut0<13> ), .Y(n844) );
  INVX1 U924 ( .A(\cacheDataOut0<10> ), .Y(n847) );
  INVX1 U925 ( .A(\cacheDataOut0<15> ), .Y(n843) );
  INVX1 U926 ( .A(\cacheDataOut1<4> ), .Y(n810) );
  INVX1 U927 ( .A(\cacheDataOut0<11> ), .Y(n846) );
  INVX1 U928 ( .A(\cacheDataOut0<9> ), .Y(n848) );
  INVX1 U929 ( .A(\cacheDataOut1<3> ), .Y(n811) );
  INVX1 U930 ( .A(n508), .Y(n797) );
  INVX1 U931 ( .A(\cacheDataOut0<7> ), .Y(n849) );
  INVX1 U932 ( .A(n737), .Y(n736) );
  INVX1 U933 ( .A(\Addr<3> ), .Y(n737) );
  INVX1 U934 ( .A(\cacheDataOut1<2> ), .Y(n812) );
  INVX1 U935 ( .A(\cacheDataOut1<1> ), .Y(n813) );
  INVX1 U936 ( .A(\cacheDataOut1<0> ), .Y(n815) );
  INVX1 U937 ( .A(\cacheDataOut0<6> ), .Y(n850) );
  INVX1 U938 ( .A(\cacheDataOut0<5> ), .Y(n851) );
  INVX1 U939 ( .A(\cacheDataOut0<4> ), .Y(n852) );
  INVX1 U940 ( .A(n439), .Y(n757) );
  INVX1 U941 ( .A(\cacheDataOut0<3> ), .Y(n853) );
  AND2X2 U942 ( .A(n439), .B(n385), .Y(n726) );
  INVX1 U943 ( .A(\cacheDataOut0<0> ), .Y(n854) );
  INVX8 U944 ( .A(n735), .Y(n731) );
  INVX8 U945 ( .A(n735), .Y(n732) );
  INVX8 U946 ( .A(n460), .Y(n860) );
  INVX8 U947 ( .A(n739), .Y(n738) );
  INVX8 U948 ( .A(n741), .Y(n740) );
  INVX8 U949 ( .A(n743), .Y(n742) );
  INVX8 U950 ( .A(n745), .Y(n744) );
  OAI21X1 U951 ( .A(n562), .B(n525), .C(n691), .Y(n752) );
  NAND3X1 U952 ( .A(n867), .B(n703), .C(n697), .Y(\nextEvictState_in<4> ) );
  NOR2X1 U953 ( .A(\wait4Cycles_in<0> ), .B(\wait4Cycles_flop<0> ), .Y(n753)
         );
  NAND3X1 U954 ( .A(n755), .B(n754), .C(n753), .Y(n756) );
  OR2X2 U955 ( .A(n758), .B(n485), .Y(n770) );
  AOI22X1 U956 ( .A(n759), .B(n574), .C(n709), .D(n770), .Y(n762) );
  NOR2X1 U957 ( .A(n392), .B(n396), .Y(n760) );
  NOR3X1 U958 ( .A(n692), .B(n860), .C(n687), .Y(n761) );
  NAND3X1 U959 ( .A(n761), .B(n500), .C(n486), .Y(\nxtState<4> ) );
  NAND2X1 U960 ( .A(n839), .B(\state<0> ), .Y(n763) );
  OAI21X1 U961 ( .A(n492), .B(n759), .C(n441), .Y(n786) );
  OAI21X1 U962 ( .A(n462), .B(n765), .C(n764), .Y(n766) );
  NOR2X1 U963 ( .A(n580), .B(n767), .Y(n768) );
  AOI21X1 U964 ( .A(n397), .B(n866), .C(n768), .Y(n769) );
  NAND3X1 U965 ( .A(n464), .B(n640), .C(n608), .Y(\nxtState<3> ) );
  AOI21X1 U966 ( .A(\nxtEvict<2> ), .B(n537), .C(n585), .Y(n772) );
  MUX2X1 U967 ( .B(n694), .A(n629), .S(memStall), .Y(n771) );
  NOR3X1 U968 ( .A(n773), .B(n397), .C(\wait4Cycles_flop<0> ), .Y(n776) );
  NOR2X1 U969 ( .A(n773), .B(\wait4Cycles_flop<0> ), .Y(n774) );
  NAND3X1 U970 ( .A(n690), .B(n699), .C(n616), .Y(n775) );
  OAI21X1 U971 ( .A(n776), .B(n447), .C(n592), .Y(n779) );
  NOR2X1 U972 ( .A(n562), .B(n420), .Y(n777) );
  OAI21X1 U973 ( .A(n620), .B(n397), .C(n777), .Y(n778) );
  NOR3X1 U974 ( .A(n505), .B(n779), .C(n655), .Y(n780) );
  NAND3X1 U975 ( .A(n560), .B(n780), .C(n558), .Y(\nxtState<2> ) );
  OAI21X1 U976 ( .A(n861), .B(n445), .C(n427), .Y(n785) );
  NAND3X1 U977 ( .A(n524), .B(n561), .C(n676), .Y(n781) );
  NAND3X1 U978 ( .A(n701), .B(n457), .C(n460), .Y(n782) );
  MUX2X1 U979 ( .B(n622), .A(n695), .S(n397), .Y(n784) );
  AND2X2 U980 ( .A(\nxtEvict<1> ), .B(n537), .Y(n783) );
  NOR3X1 U981 ( .A(n785), .B(n784), .C(n783), .Y(n788) );
  NAND3X1 U982 ( .A(n788), .B(n678), .C(n645), .Y(\nxtState<1> ) );
  OAI21X1 U983 ( .A(n615), .B(n861), .C(n674), .Y(n276) );
  AND2X2 U984 ( .A(n427), .B(n695), .Y(n789) );
  AND2X2 U985 ( .A(n703), .B(n697), .Y(n790) );
  NAND3X1 U986 ( .A(n666), .B(n790), .C(n671), .Y(n791) );
  MUX2X1 U987 ( .B(n276), .A(n627), .S(n397), .Y(n796) );
  NAND3X1 U988 ( .A(n699), .B(n635), .C(n702), .Y(n794) );
  NAND3X1 U989 ( .A(n606), .B(n637), .C(n503), .Y(n795) );
  NAND3X1 U990 ( .A(n464), .B(n796), .C(n642), .Y(\nxtState<0> ) );
  MUX2X1 U991 ( .B(victimWrite), .A(n522), .S(n797), .Y(n798) );
  MUX2X1 U992 ( .B(n850), .A(n808), .S(n814), .Y(n875) );
  MUX2X1 U993 ( .B(n852), .A(n810), .S(n814), .Y(n873) );
  NAND3X1 U994 ( .A(n444), .B(n689), .C(n647), .Y(doneWait_in) );
  OAI21X1 U995 ( .A(waitCacheHit_in), .B(n838), .C(n839), .Y(n817) );
  NAND2X1 U996 ( .A(n838), .B(waitCacheHit_in), .Y(n818) );
  AOI22X1 U997 ( .A(n838), .B(n576), .C(n539), .D(n818), .Y(n819) );
  NAND3X1 U998 ( .A(n610), .B(n639), .C(n819), .Y(stallWait_in) );
  OAI21X1 U999 ( .A(n838), .B(n432), .C(n545), .Y(n822) );
  NAND3X1 U1000 ( .A(n713), .B(n398), .C(n405), .Y(n820) );
  NAND3X1 U1001 ( .A(n488), .B(n820), .C(n457), .Y(n821) );
  OR2X2 U1002 ( .A(n483), .B(n822), .Y(cacheWr) );
  AND2X2 U1003 ( .A(n703), .B(n447), .Y(n823) );
  NAND3X1 U1004 ( .A(n390), .B(n460), .C(n823), .Y(n335) );
  MUX2X1 U1005 ( .B(n496), .A(n631), .S(n420), .Y(n824) );
  AOI21X1 U1006 ( .A(\Addr<1> ), .B(n682), .C(n824), .Y(n825) );
  AOI21X1 U1007 ( .A(\Addr<2> ), .B(n683), .C(n538), .Y(n827) );
  MUX2X1 U1008 ( .B(n561), .A(n857), .S(n715), .Y(n826) );
  NAND3X1 U1009 ( .A(n487), .B(n826), .C(n649), .Y(\cacheOff<2> ) );
  NAND3X1 U1010 ( .A(n527), .B(n828), .C(n454), .Y(n830) );
  NOR2X1 U1011 ( .A(\nxtEvict<3> ), .B(n830), .Y(n832) );
  NOR3X1 U1012 ( .A(\nxtEvict<0> ), .B(\nxtEvict<2> ), .C(\nxtEvict<1> ), .Y(
        n831) );
  AOI21X1 U1013 ( .A(n831), .B(n832), .C(n543), .Y(n836) );
  NAND2X1 U1014 ( .A(n841), .B(n442), .Y(n837) );
  OAI21X1 U1015 ( .A(n494), .B(n517), .C(n615), .Y(n855) );
  AOI21X1 U1016 ( .A(n460), .B(n618), .C(n397), .Y(\wait4Cycles_in<2> ) );
  OAI21X1 U1017 ( .A(n840), .B(victimWay), .C(valid0), .Y(n842) );
  MUX2X1 U1018 ( .B(n842), .A(n841), .S(n404), .Y(victimWrite_in) );
  MUX2X1 U1019 ( .B(n418), .A(n926), .S(n860), .Y(\memDataIn<15> ) );
  MUX2X1 U1020 ( .B(n415), .A(n927), .S(n860), .Y(\memDataIn<14> ) );
  MUX2X1 U1021 ( .B(n408), .A(n928), .S(n860), .Y(\memDataIn<13> ) );
  MUX2X1 U1022 ( .B(n409), .A(n929), .S(n860), .Y(\memDataIn<12> ) );
  MUX2X1 U1023 ( .B(n410), .A(n930), .S(n860), .Y(\memDataIn<11> ) );
  MUX2X1 U1024 ( .B(n711), .A(n931), .S(n860), .Y(\memDataIn<10> ) );
  MUX2X1 U1025 ( .B(n719), .A(n932), .S(n860), .Y(\memDataIn<9> ) );
  MUX2X1 U1026 ( .B(n416), .A(n933), .S(n860), .Y(\memDataIn<8> ) );
  MUX2X1 U1027 ( .B(n417), .A(n934), .S(n860), .Y(\memDataIn<7> ) );
  MUX2X1 U1028 ( .B(n718), .A(n935), .S(n860), .Y(\memDataIn<6> ) );
  MUX2X1 U1029 ( .B(n411), .A(n936), .S(n860), .Y(\memDataIn<5> ) );
  MUX2X1 U1030 ( .B(n716), .A(n937), .S(n860), .Y(\memDataIn<4> ) );
  MUX2X1 U1031 ( .B(n708), .A(n938), .S(n860), .Y(\memDataIn<3> ) );
  MUX2X1 U1032 ( .B(n412), .A(n939), .S(n860), .Y(\memDataIn<2> ) );
  MUX2X1 U1033 ( .B(n419), .A(n940), .S(n860), .Y(\memDataIn<1> ) );
  MUX2X1 U1034 ( .B(n394), .A(n941), .S(n860), .Y(\memDataIn<0> ) );
  MUX2X1 U1035 ( .B(n856), .A(n523), .S(n715), .Y(memWr) );
  AND2X2 U1036 ( .A(n703), .B(n457), .Y(n859) );
  AOI22X1 U1037 ( .A(n715), .B(n561), .C(n857), .D(n531), .Y(n858) );
  NAND3X1 U1038 ( .A(n491), .B(n395), .C(n464), .Y(n296) );
  NOR3X1 U1039 ( .A(n651), .B(n653), .C(n700), .Y(n293) );
  MUX2X1 U1040 ( .B(n864), .A(n907), .S(n657), .Y(n865) );
  MUX2X1 U1041 ( .B(n864), .A(n907), .S(n659), .Y(n11) );
  MUX2X1 U1042 ( .B(n624), .A(n864), .S(n540), .Y(n9) );
endmodule

