
module dff_203 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_202 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_185 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_186 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_187 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_188 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_189 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_190 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_191 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_192 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_193 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_194 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_195 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_196 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_197 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_169 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_170 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_171 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_172 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_173 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_174 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_175 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_176 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_177 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_178 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_179 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_180 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_181 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_182 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_183 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_184 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_161 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_162 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_163 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_164 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_165 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_166 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_167 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_168 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_201 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_200 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_199 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_198 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X1 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(rst), .Y(n1) );
  AND2X2 U4 ( .A(d), .B(n1), .Y(N3) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module memc_Size16_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n214, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1162), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1161), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1160), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1159), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1158), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1157), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1156), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1155), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1154), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1153), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1152), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1151), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1150), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1149), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1148), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1147), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1146), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1145), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1144), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1143), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1142), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1141), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1140), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1139), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1138), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1137), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1136), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1135), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1134), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1133), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1132), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1131), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1130), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1129), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1128), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1127), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1126), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1125), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1124), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1123), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1122), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1121), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1120), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1119), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1118), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1117), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1116), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1115), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1114), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1113), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1112), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1111), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1110), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1109), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1108), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1107), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1106), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1105), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1104), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1103), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1102), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1101), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1100), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1099), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1098), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1097), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1096), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1095), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1094), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1093), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1092), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1091), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1090), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1089), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1088), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1087), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1086), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1085), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1084), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1083), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1082), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1081), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1080), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1079), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1078), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1077), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1076), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1075), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1074), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1073), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1072), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1071), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1070), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1069), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1068), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1067), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1066), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1065), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1064), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1063), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1062), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1061), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1060), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1059), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1058), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1057), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1056), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1055), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1054), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1053), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1052), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1051), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1050), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1049), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1048), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1047), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1046), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1045), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1044), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1043), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1042), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1041), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1040), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1039), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1038), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1037), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1036), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1035), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1034), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1033), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1032), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1031), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1030), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1029), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1028), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1027), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1026), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1025), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1024), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1023), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1022), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1021), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1020), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1019), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1018), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1017), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1016), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1015), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n1014), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n1013), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n1012), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n1011), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1010), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1009), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1008), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1007), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1006), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1005), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1004), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1003), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n1002), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n1001), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n1000), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n999), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n998), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n997), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n996), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n995), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n994), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n993), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n992), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n991), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n990), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n989), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n988), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n987), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n986), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n985), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n984), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n983), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n982), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n981), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n980), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n979), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n978), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n977), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n976), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n975), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n974), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n973), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n972), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n971), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n970), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n969), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n968), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n967), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n966), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n965), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n964), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n963), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n962), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n961), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n960), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n959), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n958), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n957), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n956), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n955), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n954), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n953), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n952), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n951), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n950), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n949), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n948), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n947), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n946), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n945), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n944), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n943), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n942), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n941), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n940), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n939), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n938), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n937), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n936), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n935), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n934), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n933), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n932), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n931), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n930), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n929), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n928), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n927), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n926), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n925), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n924), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n923), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n922), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n921), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n920), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n919), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n918), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n917), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n916), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n915), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n914), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n913), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n912), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n911), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n910), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n909), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n908), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n907), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n906), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n905), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n904), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n903), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n902), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n901), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n900), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n899), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n898), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n897), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n896), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n895), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n894), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n893), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n892), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n891), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n890), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n889), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n888), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n887), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n886), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n885), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n884), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n883), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n882), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n881), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n880), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n879), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n878), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n877), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n876), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n875), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n874), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n873), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n872), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n871), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n870), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n869), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n868), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n867), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n866), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n865), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n864), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n863), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n862), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n861), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n860), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n859), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n858), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n857), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n856), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n855), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n854), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n853), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n852), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n851), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n850), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n849), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n848), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n847), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n846), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n845), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n844), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n843), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n842), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n841), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n840), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n839), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n838), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n837), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n836), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n835), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n834), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n833), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n832), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n831), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n830), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n829), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n828), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n827), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n826), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n825), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n824), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n823), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n822), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n821), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n820), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n819), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n818), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n817), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n816), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n815), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n814), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n813), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n812), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n811), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n810), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n809), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n808), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n807), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n806), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n805), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n804), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n803), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n802), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n801), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n800), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n799), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n798), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n797), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n796), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n795), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n794), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n793), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n792), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n791), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n790), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n789), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n788), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n787), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n786), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n785), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n784), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n783), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n782), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n781), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n780), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n779), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n778), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n777), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n776), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n775), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n774), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n773), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n772), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n771), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n770), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n769), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n768), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n767), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n766), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n765), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n764), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n763), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n762), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n761), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n760), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n759), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n758), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n757), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n756), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n755), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n754), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n753), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n752), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n751), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n750), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n749), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n748), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n747), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n746), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n745), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n744), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n743), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n742), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n741), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n740), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n739), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n738), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n737), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n736), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n735), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n734), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n733), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n732), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n731), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n730), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n729), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n728), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n727), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n726), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n725), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n724), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n723), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n722), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n721), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n720), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n719), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n718), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n717), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n716), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n715), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n714), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n713), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n712), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n711), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n710), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n709), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n708), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n707), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n706), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n705), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n704), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n703), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n702), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n701), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n700), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n699), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n698), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n697), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n696), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n695), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n694), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n693), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n692), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n691), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n690), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n689), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n688), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n687), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n686), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n685), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n684), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n683), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n682), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n681), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n680), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n679), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n678), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n677), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n676), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n675), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n674), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n673), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n672), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n671), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n670), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n669), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n668), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n667), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n666), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n665), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n664), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n663), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n662), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n661), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n660), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n659), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n658), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n657), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n656), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n655), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n654), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n653), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n652), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n651), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n214) );
  INVX4 U2 ( .A(n1344), .Y(n1345) );
  INVX2 U3 ( .A(n1344), .Y(n1346) );
  INVX1 U4 ( .A(n1342), .Y(n1357) );
  INVX1 U5 ( .A(n1342), .Y(n1356) );
  INVX2 U6 ( .A(n1904), .Y(n1409) );
  INVX4 U7 ( .A(n147), .Y(n237) );
  INVX4 U8 ( .A(n146), .Y(n234) );
  INVX1 U9 ( .A(n1303), .Y(N32) );
  INVX1 U10 ( .A(n1304), .Y(N31) );
  INVX1 U11 ( .A(n1305), .Y(N30) );
  INVX1 U12 ( .A(n1306), .Y(N29) );
  INVX1 U13 ( .A(n1307), .Y(N28) );
  INVX1 U14 ( .A(n1308), .Y(N27) );
  INVX1 U15 ( .A(n1309), .Y(N26) );
  INVX1 U16 ( .A(n1311), .Y(N24) );
  INVX1 U17 ( .A(n1312), .Y(N23) );
  INVX1 U18 ( .A(n1313), .Y(N22) );
  INVX1 U19 ( .A(n1314), .Y(N21) );
  INVX1 U20 ( .A(n1315), .Y(N20) );
  INVX1 U21 ( .A(n1316), .Y(N19) );
  INVX1 U22 ( .A(n1317), .Y(N18) );
  INVX1 U23 ( .A(n1318), .Y(N17) );
  INVX1 U24 ( .A(n1359), .Y(n1344) );
  INVX1 U25 ( .A(n1358), .Y(n1342) );
  INVX1 U26 ( .A(n1358), .Y(n1343) );
  INVX1 U27 ( .A(n1438), .Y(n1322) );
  INVX1 U28 ( .A(n1329), .Y(n1330) );
  INVX1 U29 ( .A(n1329), .Y(n1331) );
  INVX2 U30 ( .A(n1329), .Y(n1332) );
  INVX1 U31 ( .A(n1341), .Y(n1333) );
  INVX1 U32 ( .A(n1343), .Y(n1348) );
  INVX1 U33 ( .A(n1341), .Y(n1334) );
  INVX1 U34 ( .A(n1343), .Y(n1349) );
  INVX2 U35 ( .A(n1343), .Y(n1350) );
  INVX1 U36 ( .A(n1341), .Y(n1335) );
  INVX2 U37 ( .A(n1343), .Y(n1351) );
  INVX1 U38 ( .A(n1328), .Y(n1336) );
  INVX2 U39 ( .A(n1343), .Y(n1353) );
  INVX1 U40 ( .A(n1342), .Y(n1354) );
  INVX1 U41 ( .A(n1328), .Y(n1337) );
  INVX1 U42 ( .A(n1322), .Y(n1325) );
  INVX1 U43 ( .A(n1342), .Y(n1355) );
  INVX2 U44 ( .A(n1328), .Y(n1338) );
  INVX2 U45 ( .A(n1328), .Y(n1339) );
  INVX1 U46 ( .A(n1322), .Y(n1324) );
  INVX2 U47 ( .A(n1343), .Y(n1347) );
  INVX2 U48 ( .A(n1343), .Y(n1352) );
  INVX2 U49 ( .A(n1329), .Y(n1340) );
  INVX1 U50 ( .A(n1310), .Y(N25) );
  BUFX2 U51 ( .A(n181), .Y(n1388) );
  INVX1 U52 ( .A(n1322), .Y(n1323) );
  INVX1 U53 ( .A(n1439), .Y(n1326) );
  INVX1 U54 ( .A(n1439), .Y(n1327) );
  INVX1 U55 ( .A(n1436), .Y(n1341) );
  INVX1 U56 ( .A(n1435), .Y(n1359) );
  INVX1 U57 ( .A(N14), .Y(n1441) );
  INVX1 U58 ( .A(n1435), .Y(n1358) );
  INVX1 U59 ( .A(n1441), .Y(n1319) );
  INVX1 U60 ( .A(n1440), .Y(n1321) );
  INVX1 U61 ( .A(n1440), .Y(n1320) );
  INVX1 U62 ( .A(n228), .Y(n1362) );
  INVX1 U63 ( .A(n229), .Y(n1369) );
  INVX1 U64 ( .A(n230), .Y(n1386) );
  INVX1 U65 ( .A(n231), .Y(n1403) );
  INVX1 U66 ( .A(n1436), .Y(n1329) );
  INVX1 U67 ( .A(n1436), .Y(n1328) );
  INVX1 U68 ( .A(rst), .Y(n1434) );
  INVX8 U69 ( .A(n1), .Y(n1408) );
  BUFX2 U70 ( .A(n179), .Y(n1385) );
  BUFX2 U71 ( .A(n177), .Y(n1383) );
  BUFX2 U72 ( .A(n175), .Y(n1381) );
  BUFX2 U73 ( .A(n173), .Y(n1379) );
  BUFX2 U74 ( .A(n171), .Y(n1377) );
  BUFX2 U75 ( .A(n169), .Y(n1375) );
  BUFX2 U76 ( .A(n167), .Y(n1373) );
  BUFX2 U77 ( .A(n163), .Y(n1368) );
  BUFX2 U78 ( .A(n161), .Y(n1366) );
  BUFX2 U79 ( .A(n159), .Y(n1364) );
  BUFX2 U80 ( .A(n165), .Y(n1371) );
  BUFX2 U81 ( .A(n197), .Y(n1405) );
  INVX4 U82 ( .A(n1409), .Y(n1406) );
  AND2X2 U83 ( .A(\data_in<11> ), .B(n1406), .Y(n211) );
  INVX1 U84 ( .A(n144), .Y(n1) );
  INVX1 U85 ( .A(n212), .Y(n2) );
  INVX1 U86 ( .A(n212), .Y(n3) );
  INVX1 U87 ( .A(n212), .Y(n4) );
  INVX1 U88 ( .A(n212), .Y(n5) );
  INVX1 U89 ( .A(n212), .Y(n6) );
  INVX1 U90 ( .A(n212), .Y(n7) );
  INVX1 U91 ( .A(n212), .Y(n8) );
  INVX1 U92 ( .A(n212), .Y(n9) );
  BUFX4 U93 ( .A(n2), .Y(n10) );
  BUFX4 U94 ( .A(n2), .Y(n11) );
  BUFX4 U95 ( .A(n3), .Y(n12) );
  BUFX4 U96 ( .A(n3), .Y(n13) );
  INVX1 U97 ( .A(n227), .Y(n14) );
  INVX1 U98 ( .A(n227), .Y(n15) );
  INVX1 U99 ( .A(n227), .Y(n16) );
  INVX1 U100 ( .A(n227), .Y(n17) );
  INVX1 U101 ( .A(n227), .Y(n18) );
  INVX1 U102 ( .A(n227), .Y(n19) );
  INVX1 U103 ( .A(n227), .Y(n20) );
  INVX1 U104 ( .A(n227), .Y(n21) );
  BUFX4 U105 ( .A(n15), .Y(n22) );
  BUFX4 U106 ( .A(n15), .Y(n23) );
  INVX1 U107 ( .A(n226), .Y(n24) );
  INVX1 U108 ( .A(n226), .Y(n25) );
  INVX1 U109 ( .A(n226), .Y(n26) );
  INVX1 U110 ( .A(n226), .Y(n27) );
  INVX1 U111 ( .A(n226), .Y(n28) );
  INVX1 U112 ( .A(n226), .Y(n29) );
  INVX1 U113 ( .A(n226), .Y(n30) );
  INVX1 U114 ( .A(n226), .Y(n31) );
  BUFX4 U115 ( .A(n25), .Y(n32) );
  BUFX4 U116 ( .A(n25), .Y(n33) );
  INVX1 U117 ( .A(n225), .Y(n34) );
  INVX1 U118 ( .A(n225), .Y(n35) );
  INVX1 U119 ( .A(n225), .Y(n36) );
  INVX1 U120 ( .A(n225), .Y(n37) );
  INVX1 U121 ( .A(n225), .Y(n38) );
  INVX1 U122 ( .A(n225), .Y(n39) );
  INVX1 U123 ( .A(n225), .Y(n40) );
  INVX1 U124 ( .A(n225), .Y(n41) );
  BUFX4 U125 ( .A(n35), .Y(n42) );
  BUFX4 U126 ( .A(n35), .Y(n43) );
  BUFX2 U127 ( .A(n159), .Y(n1363) );
  BUFX2 U128 ( .A(n161), .Y(n1365) );
  BUFX2 U129 ( .A(n163), .Y(n1367) );
  BUFX2 U130 ( .A(n165), .Y(n1370) );
  BUFX2 U131 ( .A(n167), .Y(n1372) );
  BUFX2 U132 ( .A(n169), .Y(n1374) );
  BUFX2 U133 ( .A(n171), .Y(n1376) );
  BUFX2 U134 ( .A(n173), .Y(n1378) );
  BUFX2 U135 ( .A(n175), .Y(n1380) );
  BUFX2 U136 ( .A(n177), .Y(n1382) );
  BUFX2 U137 ( .A(n179), .Y(n1384) );
  BUFX2 U138 ( .A(n181), .Y(n1387) );
  AND2X2 U139 ( .A(\mem<7><1> ), .B(n1389), .Y(n44) );
  INVX1 U140 ( .A(n44), .Y(n45) );
  AND2X2 U141 ( .A(\mem<7><2> ), .B(n1389), .Y(n46) );
  INVX1 U142 ( .A(n46), .Y(n47) );
  AND2X2 U143 ( .A(\mem<7><3> ), .B(n1389), .Y(n48) );
  INVX1 U144 ( .A(n48), .Y(n49) );
  AND2X2 U145 ( .A(\mem<7><4> ), .B(n1389), .Y(n50) );
  INVX1 U146 ( .A(n50), .Y(n51) );
  AND2X2 U147 ( .A(\mem<7><5> ), .B(n1389), .Y(n52) );
  INVX1 U148 ( .A(n52), .Y(n53) );
  AND2X2 U149 ( .A(\mem<7><6> ), .B(n1389), .Y(n54) );
  INVX1 U150 ( .A(n54), .Y(n55) );
  AND2X2 U151 ( .A(\mem<7><7> ), .B(n1389), .Y(n56) );
  INVX1 U152 ( .A(n56), .Y(n57) );
  BUFX2 U153 ( .A(n183), .Y(n1389) );
  BUFX2 U154 ( .A(n183), .Y(n1390) );
  AND2X2 U155 ( .A(\mem<6><1> ), .B(n1391), .Y(n58) );
  INVX1 U156 ( .A(n58), .Y(n59) );
  AND2X2 U157 ( .A(\mem<6><2> ), .B(n1391), .Y(n60) );
  INVX1 U158 ( .A(n60), .Y(n61) );
  AND2X2 U159 ( .A(\mem<6><3> ), .B(n1391), .Y(n62) );
  INVX1 U160 ( .A(n62), .Y(n63) );
  AND2X2 U161 ( .A(\mem<6><4> ), .B(n1391), .Y(n64) );
  INVX1 U162 ( .A(n64), .Y(n65) );
  AND2X2 U163 ( .A(\mem<6><5> ), .B(n1391), .Y(n66) );
  INVX1 U164 ( .A(n66), .Y(n67) );
  AND2X2 U165 ( .A(\mem<6><6> ), .B(n1391), .Y(n68) );
  INVX1 U166 ( .A(n68), .Y(n69) );
  AND2X2 U167 ( .A(\mem<6><7> ), .B(n1391), .Y(n70) );
  INVX1 U168 ( .A(n70), .Y(n71) );
  BUFX2 U169 ( .A(n185), .Y(n1391) );
  BUFX2 U170 ( .A(n185), .Y(n1392) );
  AND2X2 U171 ( .A(\mem<5><1> ), .B(n1393), .Y(n72) );
  INVX1 U172 ( .A(n72), .Y(n73) );
  AND2X2 U173 ( .A(\mem<5><2> ), .B(n1393), .Y(n74) );
  INVX1 U174 ( .A(n74), .Y(n75) );
  AND2X2 U175 ( .A(\mem<5><3> ), .B(n1393), .Y(n76) );
  INVX1 U176 ( .A(n76), .Y(n77) );
  AND2X2 U177 ( .A(\mem<5><4> ), .B(n1393), .Y(n78) );
  INVX1 U178 ( .A(n78), .Y(n79) );
  AND2X2 U179 ( .A(\mem<5><5> ), .B(n1393), .Y(n80) );
  INVX1 U180 ( .A(n80), .Y(n81) );
  AND2X2 U181 ( .A(\mem<5><6> ), .B(n1393), .Y(n82) );
  INVX1 U182 ( .A(n82), .Y(n83) );
  AND2X2 U183 ( .A(\mem<5><7> ), .B(n1393), .Y(n84) );
  INVX1 U184 ( .A(n84), .Y(n85) );
  BUFX2 U185 ( .A(n187), .Y(n1393) );
  BUFX2 U186 ( .A(n187), .Y(n1394) );
  AND2X2 U187 ( .A(\mem<4><1> ), .B(n1395), .Y(n86) );
  INVX1 U188 ( .A(n86), .Y(n87) );
  AND2X2 U189 ( .A(\mem<4><2> ), .B(n1395), .Y(n88) );
  INVX1 U190 ( .A(n88), .Y(n89) );
  AND2X2 U191 ( .A(\mem<4><3> ), .B(n1395), .Y(n90) );
  INVX1 U192 ( .A(n90), .Y(n91) );
  AND2X2 U193 ( .A(\mem<4><4> ), .B(n1395), .Y(n92) );
  INVX1 U194 ( .A(n92), .Y(n93) );
  AND2X2 U195 ( .A(\mem<4><5> ), .B(n1395), .Y(n94) );
  INVX1 U196 ( .A(n94), .Y(n95) );
  AND2X2 U197 ( .A(\mem<4><6> ), .B(n1395), .Y(n96) );
  INVX1 U198 ( .A(n96), .Y(n97) );
  AND2X2 U199 ( .A(\mem<4><7> ), .B(n1395), .Y(n98) );
  INVX1 U200 ( .A(n98), .Y(n99) );
  BUFX2 U201 ( .A(n189), .Y(n1395) );
  BUFX2 U202 ( .A(n189), .Y(n1396) );
  AND2X2 U203 ( .A(\mem<3><1> ), .B(n1397), .Y(n100) );
  INVX1 U204 ( .A(n100), .Y(n101) );
  AND2X2 U205 ( .A(\mem<3><2> ), .B(n1397), .Y(n102) );
  INVX1 U206 ( .A(n102), .Y(n103) );
  AND2X2 U207 ( .A(\mem<3><3> ), .B(n1397), .Y(n104) );
  INVX1 U208 ( .A(n104), .Y(n105) );
  AND2X2 U209 ( .A(\mem<3><4> ), .B(n1397), .Y(n106) );
  INVX1 U210 ( .A(n106), .Y(n107) );
  AND2X2 U211 ( .A(\mem<3><5> ), .B(n1397), .Y(n108) );
  INVX1 U212 ( .A(n108), .Y(n109) );
  AND2X2 U213 ( .A(\mem<3><6> ), .B(n1397), .Y(n110) );
  INVX1 U214 ( .A(n110), .Y(n111) );
  AND2X2 U215 ( .A(\mem<3><7> ), .B(n1397), .Y(n112) );
  INVX1 U216 ( .A(n112), .Y(n113) );
  BUFX2 U217 ( .A(n191), .Y(n1397) );
  BUFX2 U218 ( .A(n191), .Y(n1398) );
  AND2X2 U219 ( .A(\mem<2><1> ), .B(n1399), .Y(n114) );
  INVX1 U220 ( .A(n114), .Y(n115) );
  AND2X2 U221 ( .A(\mem<2><2> ), .B(n1399), .Y(n116) );
  INVX1 U222 ( .A(n116), .Y(n117) );
  AND2X2 U223 ( .A(\mem<2><3> ), .B(n1399), .Y(n118) );
  INVX1 U224 ( .A(n118), .Y(n119) );
  AND2X2 U225 ( .A(\mem<2><4> ), .B(n1399), .Y(n120) );
  INVX1 U226 ( .A(n120), .Y(n121) );
  AND2X2 U227 ( .A(\mem<2><5> ), .B(n1399), .Y(n122) );
  INVX1 U228 ( .A(n122), .Y(n123) );
  AND2X2 U229 ( .A(\mem<2><6> ), .B(n1399), .Y(n124) );
  INVX1 U230 ( .A(n124), .Y(n125) );
  AND2X2 U231 ( .A(\mem<2><7> ), .B(n1399), .Y(n126) );
  INVX1 U232 ( .A(n126), .Y(n127) );
  BUFX2 U233 ( .A(n193), .Y(n1399) );
  BUFX2 U234 ( .A(n193), .Y(n1400) );
  AND2X2 U235 ( .A(\mem<1><1> ), .B(n1401), .Y(n128) );
  INVX1 U236 ( .A(n128), .Y(n129) );
  AND2X2 U237 ( .A(\mem<1><2> ), .B(n1401), .Y(n130) );
  INVX1 U238 ( .A(n130), .Y(n131) );
  AND2X2 U239 ( .A(\mem<1><3> ), .B(n1401), .Y(n132) );
  INVX1 U240 ( .A(n132), .Y(n133) );
  AND2X2 U241 ( .A(\mem<1><4> ), .B(n1401), .Y(n134) );
  INVX1 U242 ( .A(n134), .Y(n135) );
  AND2X2 U243 ( .A(\mem<1><5> ), .B(n1401), .Y(n136) );
  INVX1 U244 ( .A(n136), .Y(n137) );
  AND2X2 U245 ( .A(\mem<1><6> ), .B(n1401), .Y(n138) );
  INVX1 U246 ( .A(n138), .Y(n139) );
  AND2X2 U247 ( .A(\mem<1><7> ), .B(n1401), .Y(n140) );
  INVX1 U248 ( .A(n140), .Y(n141) );
  BUFX2 U249 ( .A(n195), .Y(n1401) );
  BUFX2 U250 ( .A(n195), .Y(n1402) );
  BUFX2 U251 ( .A(n197), .Y(n1404) );
  BUFX2 U252 ( .A(write), .Y(n142) );
  OR2X2 U253 ( .A(write), .B(rst), .Y(n143) );
  AND2X2 U254 ( .A(n142), .B(n1434), .Y(n144) );
  INVX1 U255 ( .A(n144), .Y(n145) );
  AND2X2 U256 ( .A(n1406), .B(n232), .Y(n146) );
  AND2X2 U257 ( .A(n1406), .B(n235), .Y(n147) );
  AND2X2 U258 ( .A(n1406), .B(n238), .Y(n148) );
  AND2X2 U259 ( .A(n1406), .B(n242), .Y(n149) );
  AND2X2 U260 ( .A(n1406), .B(n246), .Y(n150) );
  AND2X2 U261 ( .A(n1406), .B(n250), .Y(n151) );
  AND2X2 U262 ( .A(n1406), .B(n254), .Y(n152) );
  AND2X2 U263 ( .A(n1406), .B(n228), .Y(n153) );
  AND2X2 U264 ( .A(n1406), .B(n260), .Y(n154) );
  AND2X2 U265 ( .A(n1406), .B(n264), .Y(n155) );
  AND2X2 U266 ( .A(n1406), .B(n268), .Y(n156) );
  AND2X2 U267 ( .A(n1406), .B(n272), .Y(n157) );
  AND2X2 U268 ( .A(n1407), .B(n276), .Y(n158) );
  INVX1 U269 ( .A(n158), .Y(n159) );
  AND2X2 U270 ( .A(n1407), .B(n278), .Y(n160) );
  INVX1 U271 ( .A(n160), .Y(n161) );
  AND2X2 U272 ( .A(n1407), .B(n280), .Y(n162) );
  INVX1 U273 ( .A(n162), .Y(n163) );
  AND2X2 U274 ( .A(n1407), .B(n229), .Y(n164) );
  INVX1 U275 ( .A(n164), .Y(n165) );
  AND2X2 U276 ( .A(n1407), .B(n282), .Y(n166) );
  INVX1 U277 ( .A(n166), .Y(n167) );
  AND2X2 U278 ( .A(n1407), .B(n284), .Y(n168) );
  INVX1 U279 ( .A(n168), .Y(n169) );
  AND2X2 U280 ( .A(n1407), .B(n286), .Y(n170) );
  INVX1 U281 ( .A(n170), .Y(n171) );
  AND2X2 U282 ( .A(n1407), .B(n288), .Y(n172) );
  INVX1 U283 ( .A(n172), .Y(n173) );
  AND2X2 U284 ( .A(n1407), .B(n290), .Y(n174) );
  INVX1 U285 ( .A(n174), .Y(n175) );
  AND2X2 U286 ( .A(n1407), .B(n292), .Y(n176) );
  INVX1 U287 ( .A(n176), .Y(n177) );
  AND2X2 U288 ( .A(n1407), .B(n294), .Y(n178) );
  INVX1 U289 ( .A(n178), .Y(n179) );
  AND2X2 U290 ( .A(n1408), .B(n230), .Y(n180) );
  INVX1 U291 ( .A(n180), .Y(n181) );
  AND2X2 U292 ( .A(n1408), .B(n296), .Y(n182) );
  INVX1 U293 ( .A(n182), .Y(n183) );
  AND2X2 U294 ( .A(n1408), .B(n298), .Y(n184) );
  INVX1 U295 ( .A(n184), .Y(n185) );
  AND2X2 U296 ( .A(n1408), .B(n300), .Y(n186) );
  INVX1 U297 ( .A(n186), .Y(n187) );
  AND2X2 U298 ( .A(n1408), .B(n302), .Y(n188) );
  INVX1 U299 ( .A(n188), .Y(n189) );
  AND2X2 U300 ( .A(n1408), .B(n304), .Y(n190) );
  INVX1 U301 ( .A(n190), .Y(n191) );
  AND2X2 U302 ( .A(n1408), .B(n306), .Y(n192) );
  INVX1 U303 ( .A(n192), .Y(n193) );
  AND2X2 U304 ( .A(n1408), .B(n308), .Y(n194) );
  INVX1 U305 ( .A(n194), .Y(n195) );
  AND2X2 U306 ( .A(n1407), .B(n231), .Y(n196) );
  INVX1 U307 ( .A(n196), .Y(n197) );
  INVX1 U308 ( .A(n1437), .Y(n1436) );
  INVX1 U309 ( .A(N13), .Y(n1440) );
  AND2X1 U310 ( .A(n1438), .B(n1436), .Y(n198) );
  INVX1 U311 ( .A(n1439), .Y(n1438) );
  AND2X1 U312 ( .A(n214), .B(N14), .Y(n199) );
  BUFX2 U313 ( .A(n1474), .Y(n200) );
  INVX1 U314 ( .A(n200), .Y(n1852) );
  BUFX2 U315 ( .A(n1491), .Y(n201) );
  INVX1 U316 ( .A(n201), .Y(n1862) );
  BUFX2 U317 ( .A(n1508), .Y(n202) );
  INVX1 U318 ( .A(n202), .Y(n1872) );
  BUFX2 U319 ( .A(n1525), .Y(n203) );
  INVX1 U320 ( .A(n203), .Y(n1882) );
  BUFX2 U321 ( .A(n1542), .Y(n204) );
  INVX1 U322 ( .A(n204), .Y(n1892) );
  BUFX2 U323 ( .A(n1703), .Y(n205) );
  INVX1 U324 ( .A(n205), .Y(n1816) );
  BUFX2 U325 ( .A(n1833), .Y(n206) );
  INVX1 U326 ( .A(n206), .Y(n1902) );
  AND2X1 U327 ( .A(n1348), .B(n198), .Y(n207) );
  AND2X1 U328 ( .A(n1320), .B(n199), .Y(n208) );
  INVX1 U329 ( .A(n145), .Y(n1904) );
  AND2X1 U330 ( .A(n1435), .B(n198), .Y(n209) );
  AND2X1 U331 ( .A(n1440), .B(n199), .Y(n210) );
  AND2X2 U332 ( .A(\data_in<0> ), .B(n1408), .Y(n212) );
  AND2X2 U333 ( .A(\data_in<1> ), .B(n1408), .Y(n213) );
  AND2X2 U334 ( .A(\data_in<2> ), .B(n1408), .Y(n215) );
  AND2X2 U335 ( .A(\data_in<3> ), .B(n1408), .Y(n216) );
  AND2X2 U336 ( .A(\data_in<4> ), .B(n1408), .Y(n217) );
  AND2X2 U337 ( .A(\data_in<5> ), .B(n1408), .Y(n218) );
  AND2X2 U338 ( .A(\data_in<6> ), .B(n1408), .Y(n219) );
  AND2X2 U339 ( .A(\data_in<7> ), .B(n1408), .Y(n220) );
  AND2X2 U340 ( .A(\data_in<8> ), .B(n1408), .Y(n221) );
  AND2X2 U341 ( .A(\data_in<9> ), .B(n1408), .Y(n222) );
  AND2X2 U342 ( .A(\data_in<10> ), .B(n1408), .Y(n223) );
  AND2X2 U343 ( .A(\data_in<12> ), .B(n1408), .Y(n224) );
  AND2X2 U344 ( .A(\data_in<13> ), .B(n1406), .Y(n225) );
  AND2X2 U345 ( .A(\data_in<14> ), .B(n1408), .Y(n226) );
  AND2X2 U346 ( .A(\data_in<15> ), .B(n1408), .Y(n227) );
  AND2X1 U347 ( .A(n208), .B(n1903), .Y(n228) );
  AND2X1 U348 ( .A(n1903), .B(n210), .Y(n229) );
  AND2X1 U349 ( .A(n1903), .B(n1816), .Y(n230) );
  AND2X1 U350 ( .A(n1903), .B(n1902), .Y(n231) );
  AND2X1 U351 ( .A(n207), .B(n208), .Y(n232) );
  INVX1 U352 ( .A(n232), .Y(n233) );
  AND2X1 U353 ( .A(n208), .B(n209), .Y(n235) );
  INVX1 U354 ( .A(n235), .Y(n236) );
  AND2X1 U355 ( .A(n208), .B(n1852), .Y(n238) );
  INVX1 U356 ( .A(n238), .Y(n239) );
  INVX1 U357 ( .A(n148), .Y(n240) );
  INVX1 U358 ( .A(n148), .Y(n241) );
  AND2X1 U359 ( .A(n208), .B(n1862), .Y(n242) );
  INVX1 U360 ( .A(n242), .Y(n243) );
  INVX1 U361 ( .A(n149), .Y(n244) );
  INVX1 U362 ( .A(n149), .Y(n245) );
  AND2X1 U363 ( .A(n208), .B(n1872), .Y(n246) );
  INVX1 U364 ( .A(n246), .Y(n247) );
  INVX1 U365 ( .A(n150), .Y(n248) );
  INVX1 U366 ( .A(n150), .Y(n249) );
  AND2X1 U367 ( .A(n208), .B(n1882), .Y(n250) );
  INVX1 U368 ( .A(n250), .Y(n251) );
  INVX1 U369 ( .A(n151), .Y(n252) );
  INVX1 U370 ( .A(n151), .Y(n253) );
  AND2X1 U371 ( .A(n208), .B(n1892), .Y(n254) );
  INVX1 U372 ( .A(n254), .Y(n255) );
  INVX1 U373 ( .A(n152), .Y(n256) );
  INVX1 U374 ( .A(n152), .Y(n257) );
  INVX1 U375 ( .A(n153), .Y(n258) );
  INVX1 U376 ( .A(n153), .Y(n259) );
  AND2X1 U377 ( .A(n207), .B(n210), .Y(n260) );
  INVX1 U378 ( .A(n260), .Y(n261) );
  INVX1 U379 ( .A(n154), .Y(n262) );
  INVX1 U380 ( .A(n154), .Y(n263) );
  AND2X1 U381 ( .A(n209), .B(n210), .Y(n264) );
  INVX1 U382 ( .A(n264), .Y(n265) );
  INVX1 U383 ( .A(n155), .Y(n266) );
  INVX1 U384 ( .A(n155), .Y(n267) );
  AND2X1 U385 ( .A(n1852), .B(n210), .Y(n268) );
  INVX1 U386 ( .A(n268), .Y(n269) );
  INVX1 U387 ( .A(n156), .Y(n270) );
  INVX1 U388 ( .A(n156), .Y(n271) );
  AND2X1 U389 ( .A(n1862), .B(n210), .Y(n272) );
  INVX1 U390 ( .A(n272), .Y(n273) );
  INVX1 U391 ( .A(n157), .Y(n274) );
  INVX1 U392 ( .A(n157), .Y(n275) );
  AND2X1 U393 ( .A(n1872), .B(n210), .Y(n276) );
  INVX1 U394 ( .A(n276), .Y(n277) );
  AND2X1 U395 ( .A(n1882), .B(n210), .Y(n278) );
  INVX1 U396 ( .A(n278), .Y(n279) );
  AND2X1 U397 ( .A(n1892), .B(n210), .Y(n280) );
  INVX1 U398 ( .A(n280), .Y(n281) );
  AND2X1 U399 ( .A(n207), .B(n1816), .Y(n282) );
  INVX1 U400 ( .A(n282), .Y(n283) );
  AND2X1 U401 ( .A(n209), .B(n1816), .Y(n284) );
  INVX1 U402 ( .A(n284), .Y(n285) );
  AND2X1 U403 ( .A(n1852), .B(n1816), .Y(n286) );
  INVX1 U404 ( .A(n286), .Y(n287) );
  AND2X1 U405 ( .A(n1862), .B(n1816), .Y(n288) );
  INVX1 U406 ( .A(n288), .Y(n289) );
  AND2X1 U407 ( .A(n1872), .B(n1816), .Y(n290) );
  INVX1 U408 ( .A(n290), .Y(n291) );
  AND2X1 U409 ( .A(n1882), .B(n1816), .Y(n292) );
  INVX1 U410 ( .A(n292), .Y(n293) );
  AND2X1 U411 ( .A(n1892), .B(n1816), .Y(n294) );
  INVX1 U412 ( .A(n294), .Y(n295) );
  AND2X1 U413 ( .A(n207), .B(n1902), .Y(n296) );
  INVX1 U414 ( .A(n296), .Y(n297) );
  AND2X1 U415 ( .A(n209), .B(n1902), .Y(n298) );
  INVX1 U416 ( .A(n298), .Y(n299) );
  AND2X1 U417 ( .A(n1852), .B(n1902), .Y(n300) );
  INVX1 U418 ( .A(n300), .Y(n301) );
  AND2X1 U419 ( .A(n1862), .B(n1902), .Y(n302) );
  INVX1 U420 ( .A(n302), .Y(n303) );
  AND2X1 U421 ( .A(n1872), .B(n1902), .Y(n304) );
  INVX1 U422 ( .A(n304), .Y(n305) );
  AND2X1 U423 ( .A(n1882), .B(n1902), .Y(n306) );
  INVX1 U424 ( .A(n306), .Y(n307) );
  AND2X1 U425 ( .A(n1892), .B(n1902), .Y(n308) );
  INVX1 U426 ( .A(n308), .Y(n309) );
  INVX2 U427 ( .A(n143), .Y(n310) );
  MUX2X1 U428 ( .B(n312), .A(n313), .S(n1330), .Y(n311) );
  MUX2X1 U429 ( .B(n315), .A(n316), .S(n1330), .Y(n314) );
  MUX2X1 U430 ( .B(n318), .A(n319), .S(n1330), .Y(n317) );
  MUX2X1 U431 ( .B(n321), .A(n322), .S(n1330), .Y(n320) );
  MUX2X1 U432 ( .B(n324), .A(n325), .S(n1321), .Y(n323) );
  MUX2X1 U433 ( .B(n327), .A(n328), .S(n1330), .Y(n326) );
  MUX2X1 U434 ( .B(n330), .A(n331), .S(n1330), .Y(n329) );
  MUX2X1 U435 ( .B(n333), .A(n334), .S(n1330), .Y(n332) );
  MUX2X1 U436 ( .B(n336), .A(n337), .S(n1330), .Y(n335) );
  MUX2X1 U437 ( .B(n339), .A(n340), .S(n1321), .Y(n338) );
  MUX2X1 U438 ( .B(n342), .A(n343), .S(n1331), .Y(n341) );
  MUX2X1 U439 ( .B(n345), .A(n346), .S(n1331), .Y(n344) );
  MUX2X1 U440 ( .B(n348), .A(n349), .S(n1331), .Y(n347) );
  MUX2X1 U441 ( .B(n351), .A(n352), .S(n1331), .Y(n350) );
  MUX2X1 U442 ( .B(n354), .A(n355), .S(n1321), .Y(n353) );
  MUX2X1 U443 ( .B(n357), .A(n358), .S(n1331), .Y(n356) );
  MUX2X1 U444 ( .B(n360), .A(n361), .S(n1331), .Y(n359) );
  MUX2X1 U445 ( .B(n363), .A(n364), .S(n1331), .Y(n362) );
  MUX2X1 U446 ( .B(n366), .A(n367), .S(n1331), .Y(n365) );
  MUX2X1 U447 ( .B(n369), .A(n370), .S(n1321), .Y(n368) );
  MUX2X1 U448 ( .B(n372), .A(n373), .S(n1331), .Y(n371) );
  MUX2X1 U449 ( .B(n375), .A(n376), .S(n1331), .Y(n374) );
  MUX2X1 U450 ( .B(n378), .A(n379), .S(n1331), .Y(n377) );
  MUX2X1 U451 ( .B(n381), .A(n382), .S(n1331), .Y(n380) );
  MUX2X1 U452 ( .B(n384), .A(n385), .S(n1321), .Y(n383) );
  MUX2X1 U453 ( .B(n387), .A(n388), .S(n1332), .Y(n386) );
  MUX2X1 U454 ( .B(n390), .A(n391), .S(n1332), .Y(n389) );
  MUX2X1 U455 ( .B(n393), .A(n394), .S(n1332), .Y(n392) );
  MUX2X1 U456 ( .B(n396), .A(n397), .S(n1332), .Y(n395) );
  MUX2X1 U457 ( .B(n399), .A(n400), .S(n1321), .Y(n398) );
  MUX2X1 U458 ( .B(n402), .A(n403), .S(n1332), .Y(n401) );
  MUX2X1 U459 ( .B(n405), .A(n406), .S(n1332), .Y(n404) );
  MUX2X1 U460 ( .B(n408), .A(n409), .S(n1332), .Y(n407) );
  MUX2X1 U461 ( .B(n411), .A(n412), .S(n1332), .Y(n410) );
  MUX2X1 U462 ( .B(n414), .A(n415), .S(n1321), .Y(n413) );
  MUX2X1 U463 ( .B(n417), .A(n418), .S(n1332), .Y(n416) );
  MUX2X1 U464 ( .B(n420), .A(n421), .S(n1332), .Y(n419) );
  MUX2X1 U465 ( .B(n423), .A(n424), .S(n1332), .Y(n422) );
  MUX2X1 U466 ( .B(n426), .A(n427), .S(n1332), .Y(n425) );
  MUX2X1 U467 ( .B(n429), .A(n430), .S(n1321), .Y(n428) );
  MUX2X1 U468 ( .B(n432), .A(n433), .S(n1333), .Y(n431) );
  MUX2X1 U469 ( .B(n435), .A(n436), .S(n1333), .Y(n434) );
  MUX2X1 U470 ( .B(n438), .A(n439), .S(n1333), .Y(n437) );
  MUX2X1 U471 ( .B(n441), .A(n442), .S(n1333), .Y(n440) );
  MUX2X1 U472 ( .B(n444), .A(n445), .S(n1321), .Y(n443) );
  MUX2X1 U473 ( .B(n447), .A(n448), .S(n1333), .Y(n446) );
  MUX2X1 U474 ( .B(n450), .A(n451), .S(n1333), .Y(n449) );
  MUX2X1 U475 ( .B(n453), .A(n454), .S(n1333), .Y(n452) );
  MUX2X1 U476 ( .B(n456), .A(n457), .S(n1333), .Y(n455) );
  MUX2X1 U477 ( .B(n459), .A(n460), .S(n1321), .Y(n458) );
  MUX2X1 U478 ( .B(n462), .A(n463), .S(n1333), .Y(n461) );
  MUX2X1 U479 ( .B(n465), .A(n466), .S(n1333), .Y(n464) );
  MUX2X1 U480 ( .B(n468), .A(n469), .S(n1333), .Y(n467) );
  MUX2X1 U481 ( .B(n471), .A(n472), .S(n1333), .Y(n470) );
  MUX2X1 U482 ( .B(n474), .A(n475), .S(n1321), .Y(n473) );
  MUX2X1 U483 ( .B(n477), .A(n478), .S(n1334), .Y(n476) );
  MUX2X1 U484 ( .B(n480), .A(n481), .S(n1334), .Y(n479) );
  MUX2X1 U485 ( .B(n483), .A(n484), .S(n1334), .Y(n482) );
  MUX2X1 U486 ( .B(n486), .A(n487), .S(n1334), .Y(n485) );
  MUX2X1 U487 ( .B(n489), .A(n490), .S(n1321), .Y(n488) );
  MUX2X1 U488 ( .B(n492), .A(n493), .S(n1334), .Y(n491) );
  MUX2X1 U489 ( .B(n495), .A(n496), .S(n1334), .Y(n494) );
  MUX2X1 U490 ( .B(n498), .A(n499), .S(n1334), .Y(n497) );
  MUX2X1 U491 ( .B(n501), .A(n502), .S(n1334), .Y(n500) );
  MUX2X1 U492 ( .B(n504), .A(n505), .S(n1320), .Y(n503) );
  MUX2X1 U493 ( .B(n507), .A(n508), .S(n1334), .Y(n506) );
  MUX2X1 U494 ( .B(n510), .A(n511), .S(n1334), .Y(n509) );
  MUX2X1 U495 ( .B(n513), .A(n514), .S(n1334), .Y(n512) );
  MUX2X1 U496 ( .B(n516), .A(n517), .S(n1334), .Y(n515) );
  MUX2X1 U497 ( .B(n519), .A(n520), .S(n1320), .Y(n518) );
  MUX2X1 U498 ( .B(n522), .A(n523), .S(n1335), .Y(n521) );
  MUX2X1 U499 ( .B(n525), .A(n526), .S(n1335), .Y(n524) );
  MUX2X1 U500 ( .B(n528), .A(n529), .S(n1335), .Y(n527) );
  MUX2X1 U501 ( .B(n531), .A(n532), .S(n1335), .Y(n530) );
  MUX2X1 U502 ( .B(n534), .A(n535), .S(n1320), .Y(n533) );
  MUX2X1 U503 ( .B(n537), .A(n538), .S(n1335), .Y(n536) );
  MUX2X1 U504 ( .B(n540), .A(n541), .S(n1335), .Y(n539) );
  MUX2X1 U505 ( .B(n543), .A(n544), .S(n1335), .Y(n542) );
  MUX2X1 U506 ( .B(n546), .A(n547), .S(n1335), .Y(n545) );
  MUX2X1 U507 ( .B(n549), .A(n550), .S(n1320), .Y(n548) );
  MUX2X1 U508 ( .B(n552), .A(n553), .S(n1335), .Y(n551) );
  MUX2X1 U509 ( .B(n555), .A(n556), .S(n1335), .Y(n554) );
  MUX2X1 U510 ( .B(n558), .A(n559), .S(n1335), .Y(n557) );
  MUX2X1 U511 ( .B(n561), .A(n562), .S(n1335), .Y(n560) );
  MUX2X1 U512 ( .B(n564), .A(n565), .S(n1320), .Y(n563) );
  MUX2X1 U513 ( .B(n567), .A(n568), .S(n1336), .Y(n566) );
  MUX2X1 U514 ( .B(n570), .A(n571), .S(n1336), .Y(n569) );
  MUX2X1 U515 ( .B(n573), .A(n574), .S(n1336), .Y(n572) );
  MUX2X1 U516 ( .B(n576), .A(n577), .S(n1336), .Y(n575) );
  MUX2X1 U517 ( .B(n579), .A(n580), .S(n1320), .Y(n578) );
  MUX2X1 U518 ( .B(n582), .A(n583), .S(n1336), .Y(n581) );
  MUX2X1 U519 ( .B(n585), .A(n586), .S(n1336), .Y(n584) );
  MUX2X1 U520 ( .B(n588), .A(n589), .S(n1336), .Y(n587) );
  MUX2X1 U521 ( .B(n591), .A(n592), .S(n1336), .Y(n590) );
  MUX2X1 U522 ( .B(n594), .A(n595), .S(n1320), .Y(n593) );
  MUX2X1 U523 ( .B(n597), .A(n598), .S(n1336), .Y(n596) );
  MUX2X1 U524 ( .B(n600), .A(n601), .S(n1336), .Y(n599) );
  MUX2X1 U525 ( .B(n603), .A(n604), .S(n1336), .Y(n602) );
  MUX2X1 U526 ( .B(n606), .A(n607), .S(n1336), .Y(n605) );
  MUX2X1 U527 ( .B(n609), .A(n610), .S(n1320), .Y(n608) );
  MUX2X1 U528 ( .B(n612), .A(n613), .S(n1337), .Y(n611) );
  MUX2X1 U529 ( .B(n615), .A(n616), .S(n1337), .Y(n614) );
  MUX2X1 U530 ( .B(n618), .A(n619), .S(n1337), .Y(n617) );
  MUX2X1 U531 ( .B(n621), .A(n622), .S(n1337), .Y(n620) );
  MUX2X1 U532 ( .B(n624), .A(n625), .S(n1320), .Y(n623) );
  MUX2X1 U533 ( .B(n627), .A(n628), .S(n1337), .Y(n626) );
  MUX2X1 U534 ( .B(n630), .A(n631), .S(n1337), .Y(n629) );
  MUX2X1 U535 ( .B(n633), .A(n634), .S(n1337), .Y(n632) );
  MUX2X1 U536 ( .B(n636), .A(n637), .S(n1337), .Y(n635) );
  MUX2X1 U537 ( .B(n639), .A(n640), .S(n1320), .Y(n638) );
  MUX2X1 U538 ( .B(n642), .A(n643), .S(n1337), .Y(n641) );
  MUX2X1 U539 ( .B(n645), .A(n646), .S(n1337), .Y(n644) );
  MUX2X1 U540 ( .B(n648), .A(n649), .S(n1337), .Y(n647) );
  MUX2X1 U541 ( .B(n1163), .A(n1164), .S(n1337), .Y(n650) );
  MUX2X1 U542 ( .B(n1166), .A(n1167), .S(n1320), .Y(n1165) );
  MUX2X1 U543 ( .B(n1169), .A(n1170), .S(n1338), .Y(n1168) );
  MUX2X1 U544 ( .B(n1172), .A(n1173), .S(n1338), .Y(n1171) );
  MUX2X1 U545 ( .B(n1175), .A(n1176), .S(n1338), .Y(n1174) );
  MUX2X1 U546 ( .B(n1178), .A(n1179), .S(n1338), .Y(n1177) );
  MUX2X1 U547 ( .B(n1181), .A(n1182), .S(n1320), .Y(n1180) );
  MUX2X1 U548 ( .B(n1184), .A(n1185), .S(n1338), .Y(n1183) );
  MUX2X1 U549 ( .B(n1187), .A(n1188), .S(n1338), .Y(n1186) );
  MUX2X1 U550 ( .B(n1190), .A(n1191), .S(n1338), .Y(n1189) );
  MUX2X1 U551 ( .B(n1193), .A(n1194), .S(n1338), .Y(n1192) );
  MUX2X1 U552 ( .B(n1196), .A(n1197), .S(n1321), .Y(n1195) );
  MUX2X1 U553 ( .B(n1199), .A(n1200), .S(n1338), .Y(n1198) );
  MUX2X1 U554 ( .B(n1202), .A(n1203), .S(n1338), .Y(n1201) );
  MUX2X1 U555 ( .B(n1205), .A(n1206), .S(n1338), .Y(n1204) );
  MUX2X1 U556 ( .B(n1208), .A(n1209), .S(n1338), .Y(n1207) );
  MUX2X1 U557 ( .B(n1211), .A(n1212), .S(n1321), .Y(n1210) );
  MUX2X1 U558 ( .B(n1214), .A(n1215), .S(n1339), .Y(n1213) );
  MUX2X1 U559 ( .B(n1217), .A(n1218), .S(n1339), .Y(n1216) );
  MUX2X1 U560 ( .B(n1220), .A(n1221), .S(n1339), .Y(n1219) );
  MUX2X1 U561 ( .B(n1223), .A(n1224), .S(n1339), .Y(n1222) );
  MUX2X1 U562 ( .B(n1226), .A(n1227), .S(n1320), .Y(n1225) );
  MUX2X1 U563 ( .B(n1229), .A(n1230), .S(n1339), .Y(n1228) );
  MUX2X1 U564 ( .B(n1232), .A(n1233), .S(n1339), .Y(n1231) );
  MUX2X1 U565 ( .B(n1235), .A(n1236), .S(n1339), .Y(n1234) );
  MUX2X1 U566 ( .B(n1238), .A(n1239), .S(n1339), .Y(n1237) );
  MUX2X1 U567 ( .B(n1241), .A(n1242), .S(n1321), .Y(n1240) );
  MUX2X1 U568 ( .B(n1244), .A(n1245), .S(n1339), .Y(n1243) );
  MUX2X1 U569 ( .B(n1247), .A(n1248), .S(n1339), .Y(n1246) );
  MUX2X1 U570 ( .B(n1250), .A(n1251), .S(n1339), .Y(n1249) );
  MUX2X1 U571 ( .B(n1253), .A(n1254), .S(n1339), .Y(n1252) );
  MUX2X1 U572 ( .B(n1256), .A(n1257), .S(n1321), .Y(n1255) );
  MUX2X1 U573 ( .B(n1259), .A(n1260), .S(n1340), .Y(n1258) );
  MUX2X1 U574 ( .B(n1262), .A(n1263), .S(n1340), .Y(n1261) );
  MUX2X1 U575 ( .B(n1265), .A(n1266), .S(n1340), .Y(n1264) );
  MUX2X1 U576 ( .B(n1268), .A(n1269), .S(n1340), .Y(n1267) );
  MUX2X1 U577 ( .B(n1271), .A(n1272), .S(n1321), .Y(n1270) );
  MUX2X1 U578 ( .B(n1274), .A(n1275), .S(n1340), .Y(n1273) );
  MUX2X1 U579 ( .B(n1277), .A(n1278), .S(n1340), .Y(n1276) );
  MUX2X1 U580 ( .B(n1280), .A(n1281), .S(n1340), .Y(n1279) );
  MUX2X1 U581 ( .B(n1283), .A(n1284), .S(n1340), .Y(n1282) );
  MUX2X1 U582 ( .B(n1286), .A(n1287), .S(n1321), .Y(n1285) );
  MUX2X1 U583 ( .B(n1289), .A(n1290), .S(n1340), .Y(n1288) );
  MUX2X1 U584 ( .B(n1292), .A(n1293), .S(n1340), .Y(n1291) );
  MUX2X1 U585 ( .B(n1295), .A(n1296), .S(n1340), .Y(n1294) );
  MUX2X1 U586 ( .B(n1298), .A(n1299), .S(n1340), .Y(n1297) );
  MUX2X1 U587 ( .B(n1301), .A(n1302), .S(n1321), .Y(n1300) );
  MUX2X1 U588 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1351), .Y(n313) );
  MUX2X1 U589 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1356), .Y(n312) );
  MUX2X1 U590 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1345), .Y(n316) );
  MUX2X1 U591 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1354), .Y(n315) );
  MUX2X1 U592 ( .B(n314), .A(n311), .S(n1327), .Y(n325) );
  MUX2X1 U593 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1345), .Y(n319) );
  MUX2X1 U594 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1349), .Y(n318) );
  MUX2X1 U595 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1347), .Y(n322) );
  MUX2X1 U596 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1353), .Y(n321) );
  MUX2X1 U597 ( .B(n320), .A(n317), .S(n1327), .Y(n324) );
  MUX2X1 U598 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1350), .Y(n328) );
  MUX2X1 U599 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1352), .Y(n327) );
  MUX2X1 U600 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1345), .Y(n331) );
  MUX2X1 U601 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1353), .Y(n330) );
  MUX2X1 U602 ( .B(n329), .A(n326), .S(n1327), .Y(n340) );
  MUX2X1 U603 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1345), .Y(n334) );
  MUX2X1 U604 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1350), .Y(n333) );
  MUX2X1 U605 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1345), .Y(n337) );
  MUX2X1 U606 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1345), .Y(n336) );
  MUX2X1 U607 ( .B(n335), .A(n332), .S(n1327), .Y(n339) );
  MUX2X1 U608 ( .B(n338), .A(n323), .S(n1319), .Y(n1303) );
  MUX2X1 U609 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1351), .Y(n343) );
  MUX2X1 U610 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1352), .Y(n342) );
  MUX2X1 U611 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1350), .Y(n346) );
  MUX2X1 U612 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1353), .Y(n345) );
  MUX2X1 U613 ( .B(n344), .A(n341), .S(n1327), .Y(n355) );
  MUX2X1 U614 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1351), .Y(n349) );
  MUX2X1 U615 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1345), .Y(n348) );
  MUX2X1 U616 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1347), .Y(n352) );
  MUX2X1 U617 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1350), .Y(n351) );
  MUX2X1 U618 ( .B(n350), .A(n347), .S(n1327), .Y(n354) );
  MUX2X1 U619 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1347), .Y(n358) );
  MUX2X1 U620 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1353), .Y(n357) );
  MUX2X1 U621 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1345), .Y(n361) );
  MUX2X1 U622 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1345), .Y(n360) );
  MUX2X1 U623 ( .B(n359), .A(n356), .S(n1327), .Y(n370) );
  MUX2X1 U624 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1347), .Y(n364) );
  MUX2X1 U625 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1353), .Y(n363) );
  MUX2X1 U626 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1345), .Y(n367) );
  MUX2X1 U627 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1345), .Y(n366) );
  MUX2X1 U628 ( .B(n365), .A(n362), .S(n1327), .Y(n369) );
  MUX2X1 U629 ( .B(n368), .A(n353), .S(n1319), .Y(n1304) );
  MUX2X1 U630 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1351), .Y(n373) );
  MUX2X1 U631 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1352), .Y(n372) );
  MUX2X1 U632 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1350), .Y(n376) );
  MUX2X1 U633 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1354), .Y(n375) );
  MUX2X1 U634 ( .B(n374), .A(n371), .S(n1327), .Y(n385) );
  MUX2X1 U635 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1350), .Y(n379) );
  MUX2X1 U636 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1353), .Y(n378) );
  MUX2X1 U637 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1351), .Y(n382) );
  MUX2X1 U638 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1350), .Y(n381) );
  MUX2X1 U639 ( .B(n380), .A(n377), .S(n1327), .Y(n384) );
  MUX2X1 U640 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1345), .Y(n388) );
  MUX2X1 U641 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1345), .Y(n387) );
  MUX2X1 U642 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1345), .Y(n391) );
  MUX2X1 U643 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1345), .Y(n390) );
  MUX2X1 U644 ( .B(n389), .A(n386), .S(n1327), .Y(n400) );
  MUX2X1 U645 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1345), .Y(n394) );
  MUX2X1 U646 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1345), .Y(n393) );
  MUX2X1 U647 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1345), .Y(n397) );
  MUX2X1 U648 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1345), .Y(n396) );
  MUX2X1 U649 ( .B(n395), .A(n392), .S(n1327), .Y(n399) );
  MUX2X1 U650 ( .B(n398), .A(n383), .S(n1319), .Y(n1305) );
  MUX2X1 U651 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1345), .Y(n403) );
  MUX2X1 U652 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1345), .Y(n402) );
  MUX2X1 U653 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1345), .Y(n406) );
  MUX2X1 U654 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1345), .Y(n405) );
  MUX2X1 U655 ( .B(n404), .A(n401), .S(n1326), .Y(n415) );
  MUX2X1 U656 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1346), .Y(n409) );
  MUX2X1 U657 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1346), .Y(n408) );
  MUX2X1 U658 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1346), .Y(n412) );
  MUX2X1 U659 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1346), .Y(n411) );
  MUX2X1 U660 ( .B(n410), .A(n407), .S(n1326), .Y(n414) );
  MUX2X1 U661 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1346), .Y(n418) );
  MUX2X1 U662 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1346), .Y(n417) );
  MUX2X1 U663 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1346), .Y(n421) );
  MUX2X1 U664 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1346), .Y(n420) );
  MUX2X1 U665 ( .B(n419), .A(n416), .S(n1326), .Y(n430) );
  MUX2X1 U666 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1346), .Y(n424) );
  MUX2X1 U667 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1346), .Y(n423) );
  MUX2X1 U668 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1346), .Y(n427) );
  MUX2X1 U669 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1346), .Y(n426) );
  MUX2X1 U670 ( .B(n425), .A(n422), .S(n1326), .Y(n429) );
  MUX2X1 U671 ( .B(n428), .A(n413), .S(n1319), .Y(n1306) );
  MUX2X1 U672 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1347), .Y(n433) );
  MUX2X1 U673 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1347), .Y(n432) );
  MUX2X1 U674 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1347), .Y(n436) );
  MUX2X1 U675 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1347), .Y(n435) );
  MUX2X1 U676 ( .B(n434), .A(n431), .S(n1326), .Y(n445) );
  MUX2X1 U677 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1347), .Y(n439) );
  MUX2X1 U678 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1347), .Y(n438) );
  MUX2X1 U679 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1347), .Y(n442) );
  MUX2X1 U680 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1347), .Y(n441) );
  MUX2X1 U681 ( .B(n440), .A(n437), .S(n1326), .Y(n444) );
  MUX2X1 U682 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1347), .Y(n448) );
  MUX2X1 U683 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1347), .Y(n447) );
  MUX2X1 U684 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1347), .Y(n451) );
  MUX2X1 U685 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1347), .Y(n450) );
  MUX2X1 U686 ( .B(n449), .A(n446), .S(n1326), .Y(n460) );
  MUX2X1 U687 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1352), .Y(n454) );
  MUX2X1 U688 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1352), .Y(n453) );
  MUX2X1 U689 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1347), .Y(n457) );
  MUX2X1 U690 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1353), .Y(n456) );
  MUX2X1 U691 ( .B(n455), .A(n452), .S(n1326), .Y(n459) );
  MUX2X1 U692 ( .B(n458), .A(n443), .S(n1319), .Y(n1307) );
  MUX2X1 U693 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1351), .Y(n463) );
  MUX2X1 U694 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1351), .Y(n462) );
  MUX2X1 U695 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1352), .Y(n466) );
  MUX2X1 U696 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1350), .Y(n465) );
  MUX2X1 U697 ( .B(n464), .A(n461), .S(n1326), .Y(n475) );
  MUX2X1 U698 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1348), .Y(n469) );
  MUX2X1 U699 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1347), .Y(n468) );
  MUX2X1 U700 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1351), .Y(n472) );
  MUX2X1 U701 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1353), .Y(n471) );
  MUX2X1 U702 ( .B(n470), .A(n467), .S(n1326), .Y(n474) );
  MUX2X1 U703 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1351), .Y(n478) );
  MUX2X1 U704 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1347), .Y(n477) );
  MUX2X1 U705 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1347), .Y(n481) );
  MUX2X1 U706 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1352), .Y(n480) );
  MUX2X1 U707 ( .B(n479), .A(n476), .S(n1326), .Y(n490) );
  MUX2X1 U708 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1355), .Y(n484) );
  MUX2X1 U709 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1353), .Y(n483) );
  MUX2X1 U710 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1351), .Y(n487) );
  MUX2X1 U711 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1345), .Y(n486) );
  MUX2X1 U712 ( .B(n485), .A(n482), .S(n1326), .Y(n489) );
  MUX2X1 U713 ( .B(n488), .A(n473), .S(n1319), .Y(n1308) );
  MUX2X1 U714 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1347), .Y(n493) );
  MUX2X1 U715 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1353), .Y(n492) );
  MUX2X1 U716 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1352), .Y(n496) );
  MUX2X1 U717 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1350), .Y(n495) );
  MUX2X1 U718 ( .B(n494), .A(n491), .S(n1327), .Y(n505) );
  MUX2X1 U719 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1348), .Y(n499) );
  MUX2X1 U720 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1348), .Y(n498) );
  MUX2X1 U721 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1348), .Y(n502) );
  MUX2X1 U722 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1348), .Y(n501) );
  MUX2X1 U723 ( .B(n500), .A(n497), .S(n1323), .Y(n504) );
  MUX2X1 U724 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1348), .Y(n508) );
  MUX2X1 U725 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1348), .Y(n507) );
  MUX2X1 U726 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1348), .Y(n511) );
  MUX2X1 U727 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1348), .Y(n510) );
  MUX2X1 U728 ( .B(n509), .A(n506), .S(n1323), .Y(n520) );
  MUX2X1 U729 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1348), .Y(n514) );
  MUX2X1 U730 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1348), .Y(n513) );
  MUX2X1 U731 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1348), .Y(n517) );
  MUX2X1 U732 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1348), .Y(n516) );
  MUX2X1 U733 ( .B(n515), .A(n512), .S(n1326), .Y(n519) );
  MUX2X1 U734 ( .B(n518), .A(n503), .S(n1319), .Y(n1309) );
  MUX2X1 U735 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1349), .Y(n523) );
  MUX2X1 U736 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1349), .Y(n522) );
  MUX2X1 U737 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1349), .Y(n526) );
  MUX2X1 U738 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1349), .Y(n525) );
  MUX2X1 U739 ( .B(n524), .A(n521), .S(n1323), .Y(n535) );
  MUX2X1 U740 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1349), .Y(n529) );
  MUX2X1 U741 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1349), .Y(n528) );
  MUX2X1 U742 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1349), .Y(n532) );
  MUX2X1 U743 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1349), .Y(n531) );
  MUX2X1 U744 ( .B(n530), .A(n527), .S(n1327), .Y(n534) );
  MUX2X1 U745 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1349), .Y(n538) );
  MUX2X1 U746 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1349), .Y(n537) );
  MUX2X1 U747 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1349), .Y(n541) );
  MUX2X1 U748 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1349), .Y(n540) );
  MUX2X1 U749 ( .B(n539), .A(n536), .S(n1323), .Y(n550) );
  MUX2X1 U750 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1350), .Y(n544) );
  MUX2X1 U751 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1350), .Y(n543) );
  MUX2X1 U752 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1350), .Y(n547) );
  MUX2X1 U753 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1350), .Y(n546) );
  MUX2X1 U754 ( .B(n545), .A(n542), .S(n1323), .Y(n549) );
  MUX2X1 U755 ( .B(n548), .A(n533), .S(n1319), .Y(n1310) );
  MUX2X1 U756 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1350), .Y(n553) );
  MUX2X1 U757 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1350), .Y(n552) );
  MUX2X1 U758 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1350), .Y(n556) );
  MUX2X1 U759 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1350), .Y(n555) );
  MUX2X1 U760 ( .B(n554), .A(n551), .S(n1325), .Y(n565) );
  MUX2X1 U761 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1350), .Y(n559) );
  MUX2X1 U762 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1350), .Y(n558) );
  MUX2X1 U763 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1350), .Y(n562) );
  MUX2X1 U764 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1350), .Y(n561) );
  MUX2X1 U765 ( .B(n560), .A(n557), .S(n1326), .Y(n564) );
  MUX2X1 U766 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1351), .Y(n568) );
  MUX2X1 U767 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1351), .Y(n567) );
  MUX2X1 U768 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1351), .Y(n571) );
  MUX2X1 U769 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1351), .Y(n570) );
  MUX2X1 U770 ( .B(n569), .A(n566), .S(n1325), .Y(n580) );
  MUX2X1 U771 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1351), .Y(n574) );
  MUX2X1 U772 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1351), .Y(n573) );
  MUX2X1 U773 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1351), .Y(n577) );
  MUX2X1 U774 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1351), .Y(n576) );
  MUX2X1 U775 ( .B(n575), .A(n572), .S(n1323), .Y(n579) );
  MUX2X1 U776 ( .B(n578), .A(n563), .S(n1319), .Y(n1311) );
  MUX2X1 U777 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1351), .Y(n583) );
  MUX2X1 U778 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1351), .Y(n582) );
  MUX2X1 U779 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1351), .Y(n586) );
  MUX2X1 U780 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1351), .Y(n585) );
  MUX2X1 U781 ( .B(n584), .A(n581), .S(n1325), .Y(n595) );
  MUX2X1 U782 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1352), .Y(n589) );
  MUX2X1 U783 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1352), .Y(n588) );
  MUX2X1 U784 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1352), .Y(n592) );
  MUX2X1 U785 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1352), .Y(n591) );
  MUX2X1 U786 ( .B(n590), .A(n587), .S(n1325), .Y(n594) );
  MUX2X1 U787 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1352), .Y(n598) );
  MUX2X1 U788 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1352), .Y(n597) );
  MUX2X1 U789 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1352), .Y(n601) );
  MUX2X1 U790 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1352), .Y(n600) );
  MUX2X1 U791 ( .B(n599), .A(n596), .S(n1325), .Y(n610) );
  MUX2X1 U792 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1352), .Y(n604) );
  MUX2X1 U793 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1352), .Y(n603) );
  MUX2X1 U794 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1352), .Y(n607) );
  MUX2X1 U795 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1352), .Y(n606) );
  MUX2X1 U796 ( .B(n605), .A(n602), .S(n1325), .Y(n609) );
  MUX2X1 U797 ( .B(n608), .A(n593), .S(n1319), .Y(n1312) );
  MUX2X1 U798 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1353), .Y(n613) );
  MUX2X1 U799 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1353), .Y(n612) );
  MUX2X1 U800 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1353), .Y(n616) );
  MUX2X1 U801 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1353), .Y(n615) );
  MUX2X1 U802 ( .B(n614), .A(n611), .S(n1325), .Y(n625) );
  MUX2X1 U803 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1353), .Y(n619) );
  MUX2X1 U804 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1353), .Y(n618) );
  MUX2X1 U805 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1353), .Y(n622) );
  MUX2X1 U806 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1353), .Y(n621) );
  MUX2X1 U807 ( .B(n620), .A(n617), .S(n1325), .Y(n624) );
  MUX2X1 U808 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1353), .Y(n628) );
  MUX2X1 U809 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1353), .Y(n627) );
  MUX2X1 U810 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1353), .Y(n631) );
  MUX2X1 U811 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1353), .Y(n630) );
  MUX2X1 U812 ( .B(n629), .A(n626), .S(n1325), .Y(n640) );
  MUX2X1 U813 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1354), .Y(n634) );
  MUX2X1 U814 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1354), .Y(n633) );
  MUX2X1 U815 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1354), .Y(n637) );
  MUX2X1 U816 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1354), .Y(n636) );
  MUX2X1 U817 ( .B(n635), .A(n632), .S(n1325), .Y(n639) );
  MUX2X1 U818 ( .B(n638), .A(n623), .S(n1319), .Y(n1313) );
  MUX2X1 U819 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1354), .Y(n643) );
  MUX2X1 U820 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1354), .Y(n642) );
  MUX2X1 U821 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1354), .Y(n646) );
  MUX2X1 U822 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1354), .Y(n645) );
  MUX2X1 U823 ( .B(n644), .A(n641), .S(n1325), .Y(n1167) );
  MUX2X1 U824 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1354), .Y(n649) );
  MUX2X1 U825 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1354), .Y(n648) );
  MUX2X1 U826 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1354), .Y(n1164) );
  MUX2X1 U827 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1354), .Y(n1163) );
  MUX2X1 U828 ( .B(n650), .A(n647), .S(n1325), .Y(n1166) );
  MUX2X1 U829 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1355), .Y(n1170) );
  MUX2X1 U830 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1355), .Y(n1169) );
  MUX2X1 U831 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1355), .Y(n1173) );
  MUX2X1 U832 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1355), .Y(n1172) );
  MUX2X1 U833 ( .B(n1171), .A(n1168), .S(n1325), .Y(n1182) );
  MUX2X1 U834 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1355), .Y(n1176) );
  MUX2X1 U835 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1355), .Y(n1175) );
  MUX2X1 U836 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1355), .Y(n1179) );
  MUX2X1 U837 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1355), .Y(n1178) );
  MUX2X1 U838 ( .B(n1177), .A(n1174), .S(n1325), .Y(n1181) );
  MUX2X1 U839 ( .B(n1180), .A(n1165), .S(n1319), .Y(n1314) );
  MUX2X1 U840 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1355), .Y(n1185) );
  MUX2X1 U841 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1355), .Y(n1184) );
  MUX2X1 U842 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1355), .Y(n1188) );
  MUX2X1 U843 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1355), .Y(n1187) );
  MUX2X1 U844 ( .B(n1186), .A(n1183), .S(n1324), .Y(n1197) );
  MUX2X1 U845 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1356), .Y(n1191) );
  MUX2X1 U846 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1356), .Y(n1190) );
  MUX2X1 U847 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1356), .Y(n1194) );
  MUX2X1 U848 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1356), .Y(n1193) );
  MUX2X1 U849 ( .B(n1192), .A(n1189), .S(n1324), .Y(n1196) );
  MUX2X1 U850 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1356), .Y(n1200) );
  MUX2X1 U851 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1356), .Y(n1199) );
  MUX2X1 U852 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1356), .Y(n1203) );
  MUX2X1 U853 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1356), .Y(n1202) );
  MUX2X1 U854 ( .B(n1201), .A(n1198), .S(n1324), .Y(n1212) );
  MUX2X1 U855 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1356), .Y(n1206) );
  MUX2X1 U856 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1356), .Y(n1205) );
  MUX2X1 U857 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1356), .Y(n1209) );
  MUX2X1 U858 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1356), .Y(n1208) );
  MUX2X1 U859 ( .B(n1207), .A(n1204), .S(n1324), .Y(n1211) );
  MUX2X1 U860 ( .B(n1210), .A(n1195), .S(n1319), .Y(n1315) );
  MUX2X1 U861 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1355), .Y(n1215) );
  MUX2X1 U862 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1345), .Y(n1214) );
  MUX2X1 U863 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1347), .Y(n1218) );
  MUX2X1 U864 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1350), .Y(n1217) );
  MUX2X1 U865 ( .B(n1216), .A(n1213), .S(n1324), .Y(n1227) );
  MUX2X1 U866 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1352), .Y(n1221) );
  MUX2X1 U867 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1353), .Y(n1220) );
  MUX2X1 U868 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1351), .Y(n1224) );
  MUX2X1 U869 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1353), .Y(n1223) );
  MUX2X1 U870 ( .B(n1222), .A(n1219), .S(n1324), .Y(n1226) );
  MUX2X1 U871 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1352), .Y(n1230) );
  MUX2X1 U872 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1345), .Y(n1229) );
  MUX2X1 U873 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1345), .Y(n1233) );
  MUX2X1 U874 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1347), .Y(n1232) );
  MUX2X1 U875 ( .B(n1231), .A(n1228), .S(n1324), .Y(n1242) );
  MUX2X1 U876 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1356), .Y(n1236) );
  MUX2X1 U877 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1356), .Y(n1235) );
  MUX2X1 U878 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1346), .Y(n1239) );
  MUX2X1 U879 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1355), .Y(n1238) );
  MUX2X1 U880 ( .B(n1237), .A(n1234), .S(n1324), .Y(n1241) );
  MUX2X1 U881 ( .B(n1240), .A(n1225), .S(n1319), .Y(n1316) );
  MUX2X1 U882 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1357), .Y(n1245) );
  MUX2X1 U883 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1346), .Y(n1244) );
  MUX2X1 U884 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1359), .Y(n1248) );
  MUX2X1 U885 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1353), .Y(n1247) );
  MUX2X1 U886 ( .B(n1246), .A(n1243), .S(n1324), .Y(n1257) );
  MUX2X1 U887 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1345), .Y(n1251) );
  MUX2X1 U888 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1357), .Y(n1250) );
  MUX2X1 U889 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1354), .Y(n1254) );
  MUX2X1 U890 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1351), .Y(n1253) );
  MUX2X1 U891 ( .B(n1252), .A(n1249), .S(n1324), .Y(n1256) );
  MUX2X1 U892 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1357), .Y(n1260) );
  MUX2X1 U893 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1357), .Y(n1259) );
  MUX2X1 U894 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1357), .Y(n1263) );
  MUX2X1 U895 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1357), .Y(n1262) );
  MUX2X1 U896 ( .B(n1261), .A(n1258), .S(n1324), .Y(n1272) );
  MUX2X1 U897 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1357), .Y(n1266) );
  MUX2X1 U898 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1357), .Y(n1265) );
  MUX2X1 U899 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1357), .Y(n1269) );
  MUX2X1 U900 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1357), .Y(n1268) );
  MUX2X1 U901 ( .B(n1267), .A(n1264), .S(n1324), .Y(n1271) );
  MUX2X1 U902 ( .B(n1270), .A(n1255), .S(n1319), .Y(n1317) );
  MUX2X1 U903 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1357), .Y(n1275) );
  MUX2X1 U904 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1357), .Y(n1274) );
  MUX2X1 U905 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1357), .Y(n1278) );
  MUX2X1 U906 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1357), .Y(n1277) );
  MUX2X1 U907 ( .B(n1276), .A(n1273), .S(n1323), .Y(n1287) );
  MUX2X1 U908 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1352), .Y(n1281) );
  MUX2X1 U909 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1352), .Y(n1280) );
  MUX2X1 U910 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1346), .Y(n1284) );
  MUX2X1 U911 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1352), .Y(n1283) );
  MUX2X1 U912 ( .B(n1282), .A(n1279), .S(n1323), .Y(n1286) );
  MUX2X1 U913 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1345), .Y(n1290) );
  MUX2X1 U914 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1347), .Y(n1289) );
  MUX2X1 U915 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1357), .Y(n1293) );
  MUX2X1 U916 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1351), .Y(n1292) );
  MUX2X1 U917 ( .B(n1291), .A(n1288), .S(n1323), .Y(n1302) );
  MUX2X1 U918 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1345), .Y(n1296) );
  MUX2X1 U919 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1350), .Y(n1295) );
  MUX2X1 U920 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1350), .Y(n1299) );
  MUX2X1 U921 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1350), .Y(n1298) );
  MUX2X1 U922 ( .B(n1297), .A(n1294), .S(n1323), .Y(n1301) );
  MUX2X1 U923 ( .B(n1300), .A(n1285), .S(n1319), .Y(n1318) );
  INVX1 U924 ( .A(N12), .Y(n1439) );
  AND2X2 U925 ( .A(n1360), .B(N29), .Y(\data_out<3> ) );
  INVX1 U926 ( .A(n143), .Y(n1360) );
  INVX1 U927 ( .A(n143), .Y(n1361) );
  INVX1 U928 ( .A(N11), .Y(n1437) );
  INVX1 U929 ( .A(N10), .Y(n1435) );
  INVX8 U930 ( .A(n1409), .Y(n1407) );
  INVX8 U931 ( .A(n213), .Y(n1410) );
  INVX8 U932 ( .A(n213), .Y(n1411) );
  INVX8 U933 ( .A(n215), .Y(n1412) );
  INVX8 U934 ( .A(n215), .Y(n1413) );
  INVX8 U935 ( .A(n216), .Y(n1414) );
  INVX8 U936 ( .A(n216), .Y(n1415) );
  INVX8 U937 ( .A(n217), .Y(n1416) );
  INVX8 U938 ( .A(n217), .Y(n1417) );
  INVX8 U939 ( .A(n218), .Y(n1418) );
  INVX8 U940 ( .A(n218), .Y(n1419) );
  INVX8 U941 ( .A(n219), .Y(n1420) );
  INVX8 U942 ( .A(n219), .Y(n1421) );
  INVX8 U943 ( .A(n220), .Y(n1422) );
  INVX8 U944 ( .A(n220), .Y(n1423) );
  INVX8 U945 ( .A(n221), .Y(n1424) );
  INVX8 U946 ( .A(n221), .Y(n1425) );
  INVX8 U947 ( .A(n222), .Y(n1426) );
  INVX8 U948 ( .A(n222), .Y(n1427) );
  INVX8 U949 ( .A(n223), .Y(n1428) );
  INVX8 U950 ( .A(n223), .Y(n1429) );
  INVX8 U951 ( .A(n211), .Y(n1430) );
  INVX8 U952 ( .A(n211), .Y(n1431) );
  INVX8 U953 ( .A(n224), .Y(n1432) );
  INVX8 U954 ( .A(n224), .Y(n1433) );
  AND2X2 U955 ( .A(n310), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U956 ( .A(n1361), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U957 ( .A(n1361), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U958 ( .A(n1361), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U959 ( .A(n310), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U960 ( .A(n310), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U961 ( .A(n1360), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U962 ( .A(n310), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U963 ( .A(n1360), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U964 ( .A(n310), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U965 ( .A(n310), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U966 ( .A(n1360), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U967 ( .A(n310), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U968 ( .A(n1361), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U969 ( .A(n310), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U970 ( .A(\mem<31><0> ), .B(n234), .Y(n1442) );
  OAI21X1 U971 ( .A(n233), .B(n4), .C(n1442), .Y(n651) );
  NAND2X1 U972 ( .A(\mem<31><1> ), .B(n234), .Y(n1443) );
  OAI21X1 U973 ( .A(n1411), .B(n233), .C(n1443), .Y(n652) );
  NAND2X1 U974 ( .A(\mem<31><2> ), .B(n234), .Y(n1444) );
  OAI21X1 U975 ( .A(n1413), .B(n233), .C(n1444), .Y(n653) );
  NAND2X1 U976 ( .A(\mem<31><3> ), .B(n234), .Y(n1445) );
  OAI21X1 U977 ( .A(n1415), .B(n233), .C(n1445), .Y(n654) );
  NAND2X1 U978 ( .A(\mem<31><4> ), .B(n234), .Y(n1446) );
  OAI21X1 U979 ( .A(n1417), .B(n233), .C(n1446), .Y(n655) );
  NAND2X1 U980 ( .A(\mem<31><5> ), .B(n234), .Y(n1447) );
  OAI21X1 U981 ( .A(n1419), .B(n233), .C(n1447), .Y(n656) );
  NAND2X1 U982 ( .A(\mem<31><6> ), .B(n234), .Y(n1448) );
  OAI21X1 U983 ( .A(n1421), .B(n233), .C(n1448), .Y(n657) );
  NAND2X1 U984 ( .A(\mem<31><7> ), .B(n234), .Y(n1449) );
  OAI21X1 U985 ( .A(n1423), .B(n233), .C(n1449), .Y(n658) );
  NAND2X1 U986 ( .A(\mem<31><8> ), .B(n234), .Y(n1450) );
  OAI21X1 U987 ( .A(n1425), .B(n233), .C(n1450), .Y(n659) );
  NAND2X1 U988 ( .A(\mem<31><9> ), .B(n234), .Y(n1451) );
  OAI21X1 U989 ( .A(n1427), .B(n233), .C(n1451), .Y(n660) );
  NAND2X1 U990 ( .A(\mem<31><10> ), .B(n234), .Y(n1452) );
  OAI21X1 U991 ( .A(n1429), .B(n233), .C(n1452), .Y(n661) );
  NAND2X1 U992 ( .A(\mem<31><11> ), .B(n234), .Y(n1453) );
  OAI21X1 U993 ( .A(n1430), .B(n233), .C(n1453), .Y(n662) );
  NAND2X1 U994 ( .A(\mem<31><12> ), .B(n234), .Y(n1454) );
  OAI21X1 U995 ( .A(n1433), .B(n233), .C(n1454), .Y(n663) );
  NAND2X1 U996 ( .A(\mem<31><13> ), .B(n234), .Y(n1455) );
  OAI21X1 U997 ( .A(n43), .B(n233), .C(n1455), .Y(n664) );
  NAND2X1 U998 ( .A(\mem<31><14> ), .B(n234), .Y(n1456) );
  OAI21X1 U999 ( .A(n33), .B(n233), .C(n1456), .Y(n665) );
  NAND2X1 U1000 ( .A(\mem<31><15> ), .B(n234), .Y(n1457) );
  OAI21X1 U1001 ( .A(n23), .B(n233), .C(n1457), .Y(n666) );
  NAND2X1 U1002 ( .A(\mem<30><0> ), .B(n237), .Y(n1458) );
  OAI21X1 U1003 ( .A(n236), .B(n8), .C(n1458), .Y(n667) );
  NAND2X1 U1004 ( .A(\mem<30><1> ), .B(n237), .Y(n1459) );
  OAI21X1 U1005 ( .A(n236), .B(n1411), .C(n1459), .Y(n668) );
  NAND2X1 U1006 ( .A(\mem<30><2> ), .B(n237), .Y(n1460) );
  OAI21X1 U1007 ( .A(n236), .B(n1413), .C(n1460), .Y(n669) );
  NAND2X1 U1008 ( .A(\mem<30><3> ), .B(n237), .Y(n1461) );
  OAI21X1 U1009 ( .A(n236), .B(n1415), .C(n1461), .Y(n670) );
  NAND2X1 U1010 ( .A(\mem<30><4> ), .B(n237), .Y(n1462) );
  OAI21X1 U1011 ( .A(n236), .B(n1417), .C(n1462), .Y(n671) );
  NAND2X1 U1012 ( .A(\mem<30><5> ), .B(n237), .Y(n1463) );
  OAI21X1 U1013 ( .A(n236), .B(n1419), .C(n1463), .Y(n672) );
  NAND2X1 U1014 ( .A(\mem<30><6> ), .B(n237), .Y(n1464) );
  OAI21X1 U1015 ( .A(n236), .B(n1421), .C(n1464), .Y(n673) );
  NAND2X1 U1016 ( .A(\mem<30><7> ), .B(n237), .Y(n1465) );
  OAI21X1 U1017 ( .A(n236), .B(n1423), .C(n1465), .Y(n674) );
  NAND2X1 U1018 ( .A(\mem<30><8> ), .B(n237), .Y(n1466) );
  OAI21X1 U1019 ( .A(n236), .B(n1424), .C(n1466), .Y(n675) );
  NAND2X1 U1020 ( .A(\mem<30><9> ), .B(n237), .Y(n1467) );
  OAI21X1 U1021 ( .A(n236), .B(n1426), .C(n1467), .Y(n676) );
  NAND2X1 U1022 ( .A(\mem<30><10> ), .B(n237), .Y(n1468) );
  OAI21X1 U1023 ( .A(n236), .B(n1428), .C(n1468), .Y(n677) );
  NAND2X1 U1024 ( .A(\mem<30><11> ), .B(n237), .Y(n1469) );
  OAI21X1 U1025 ( .A(n236), .B(n1431), .C(n1469), .Y(n678) );
  NAND2X1 U1026 ( .A(\mem<30><12> ), .B(n237), .Y(n1470) );
  OAI21X1 U1027 ( .A(n236), .B(n1432), .C(n1470), .Y(n679) );
  NAND2X1 U1028 ( .A(\mem<30><13> ), .B(n237), .Y(n1471) );
  OAI21X1 U1029 ( .A(n236), .B(n40), .C(n1471), .Y(n680) );
  NAND2X1 U1030 ( .A(\mem<30><14> ), .B(n237), .Y(n1472) );
  OAI21X1 U1031 ( .A(n236), .B(n30), .C(n1472), .Y(n681) );
  NAND2X1 U1032 ( .A(\mem<30><15> ), .B(n237), .Y(n1473) );
  OAI21X1 U1033 ( .A(n236), .B(n20), .C(n1473), .Y(n682) );
  NAND3X1 U1034 ( .A(n1351), .B(n1438), .C(n1437), .Y(n1474) );
  NAND2X1 U1035 ( .A(\mem<29><0> ), .B(n241), .Y(n1475) );
  OAI21X1 U1036 ( .A(n239), .B(n7), .C(n1475), .Y(n683) );
  NAND2X1 U1037 ( .A(\mem<29><1> ), .B(n241), .Y(n1476) );
  OAI21X1 U1038 ( .A(n239), .B(n1410), .C(n1476), .Y(n684) );
  NAND2X1 U1039 ( .A(\mem<29><2> ), .B(n241), .Y(n1477) );
  OAI21X1 U1040 ( .A(n239), .B(n1412), .C(n1477), .Y(n685) );
  NAND2X1 U1041 ( .A(\mem<29><3> ), .B(n241), .Y(n1478) );
  OAI21X1 U1042 ( .A(n239), .B(n1414), .C(n1478), .Y(n686) );
  NAND2X1 U1043 ( .A(\mem<29><4> ), .B(n241), .Y(n1479) );
  OAI21X1 U1044 ( .A(n239), .B(n1416), .C(n1479), .Y(n687) );
  NAND2X1 U1045 ( .A(\mem<29><5> ), .B(n241), .Y(n1480) );
  OAI21X1 U1046 ( .A(n239), .B(n1418), .C(n1480), .Y(n688) );
  NAND2X1 U1047 ( .A(\mem<29><6> ), .B(n241), .Y(n1481) );
  OAI21X1 U1048 ( .A(n239), .B(n1420), .C(n1481), .Y(n689) );
  NAND2X1 U1049 ( .A(\mem<29><7> ), .B(n241), .Y(n1482) );
  OAI21X1 U1050 ( .A(n239), .B(n1422), .C(n1482), .Y(n690) );
  NAND2X1 U1051 ( .A(\mem<29><8> ), .B(n240), .Y(n1483) );
  OAI21X1 U1052 ( .A(n239), .B(n1425), .C(n1483), .Y(n691) );
  NAND2X1 U1053 ( .A(\mem<29><9> ), .B(n240), .Y(n1484) );
  OAI21X1 U1054 ( .A(n239), .B(n1427), .C(n1484), .Y(n692) );
  NAND2X1 U1055 ( .A(\mem<29><10> ), .B(n240), .Y(n1485) );
  OAI21X1 U1056 ( .A(n239), .B(n1429), .C(n1485), .Y(n693) );
  NAND2X1 U1057 ( .A(\mem<29><11> ), .B(n240), .Y(n1486) );
  OAI21X1 U1058 ( .A(n239), .B(n1430), .C(n1486), .Y(n694) );
  NAND2X1 U1059 ( .A(\mem<29><12> ), .B(n240), .Y(n1487) );
  OAI21X1 U1060 ( .A(n239), .B(n1433), .C(n1487), .Y(n695) );
  NAND2X1 U1061 ( .A(\mem<29><13> ), .B(n240), .Y(n1488) );
  OAI21X1 U1062 ( .A(n239), .B(n41), .C(n1488), .Y(n696) );
  NAND2X1 U1063 ( .A(\mem<29><14> ), .B(n240), .Y(n1489) );
  OAI21X1 U1064 ( .A(n239), .B(n31), .C(n1489), .Y(n697) );
  NAND2X1 U1065 ( .A(\mem<29><15> ), .B(n240), .Y(n1490) );
  OAI21X1 U1066 ( .A(n239), .B(n21), .C(n1490), .Y(n698) );
  NAND3X1 U1067 ( .A(n1438), .B(n1437), .C(n1435), .Y(n1491) );
  NAND2X1 U1068 ( .A(\mem<28><0> ), .B(n245), .Y(n1492) );
  OAI21X1 U1069 ( .A(n243), .B(n10), .C(n1492), .Y(n699) );
  NAND2X1 U1070 ( .A(\mem<28><1> ), .B(n245), .Y(n1493) );
  OAI21X1 U1071 ( .A(n243), .B(n1411), .C(n1493), .Y(n700) );
  NAND2X1 U1072 ( .A(\mem<28><2> ), .B(n245), .Y(n1494) );
  OAI21X1 U1073 ( .A(n243), .B(n1413), .C(n1494), .Y(n701) );
  NAND2X1 U1074 ( .A(\mem<28><3> ), .B(n245), .Y(n1495) );
  OAI21X1 U1075 ( .A(n243), .B(n1415), .C(n1495), .Y(n702) );
  NAND2X1 U1076 ( .A(\mem<28><4> ), .B(n245), .Y(n1496) );
  OAI21X1 U1077 ( .A(n243), .B(n1417), .C(n1496), .Y(n703) );
  NAND2X1 U1078 ( .A(\mem<28><5> ), .B(n245), .Y(n1497) );
  OAI21X1 U1079 ( .A(n243), .B(n1419), .C(n1497), .Y(n704) );
  NAND2X1 U1080 ( .A(\mem<28><6> ), .B(n245), .Y(n1498) );
  OAI21X1 U1081 ( .A(n243), .B(n1421), .C(n1498), .Y(n705) );
  NAND2X1 U1082 ( .A(\mem<28><7> ), .B(n245), .Y(n1499) );
  OAI21X1 U1083 ( .A(n243), .B(n1423), .C(n1499), .Y(n706) );
  NAND2X1 U1084 ( .A(\mem<28><8> ), .B(n244), .Y(n1500) );
  OAI21X1 U1085 ( .A(n243), .B(n1424), .C(n1500), .Y(n707) );
  NAND2X1 U1086 ( .A(\mem<28><9> ), .B(n244), .Y(n1501) );
  OAI21X1 U1087 ( .A(n243), .B(n1426), .C(n1501), .Y(n708) );
  NAND2X1 U1088 ( .A(\mem<28><10> ), .B(n244), .Y(n1502) );
  OAI21X1 U1089 ( .A(n243), .B(n1428), .C(n1502), .Y(n709) );
  NAND2X1 U1090 ( .A(\mem<28><11> ), .B(n244), .Y(n1503) );
  OAI21X1 U1091 ( .A(n243), .B(n1431), .C(n1503), .Y(n710) );
  NAND2X1 U1092 ( .A(\mem<28><12> ), .B(n244), .Y(n1504) );
  OAI21X1 U1093 ( .A(n243), .B(n1432), .C(n1504), .Y(n711) );
  NAND2X1 U1094 ( .A(\mem<28><13> ), .B(n244), .Y(n1505) );
  OAI21X1 U1095 ( .A(n243), .B(n41), .C(n1505), .Y(n712) );
  NAND2X1 U1096 ( .A(\mem<28><14> ), .B(n244), .Y(n1506) );
  OAI21X1 U1097 ( .A(n243), .B(n31), .C(n1506), .Y(n713) );
  NAND2X1 U1098 ( .A(\mem<28><15> ), .B(n244), .Y(n1507) );
  OAI21X1 U1099 ( .A(n243), .B(n21), .C(n1507), .Y(n714) );
  NAND3X1 U1100 ( .A(n1347), .B(n1436), .C(n1439), .Y(n1508) );
  NAND2X1 U1101 ( .A(\mem<27><0> ), .B(n249), .Y(n1509) );
  OAI21X1 U1102 ( .A(n247), .B(n9), .C(n1509), .Y(n715) );
  NAND2X1 U1103 ( .A(\mem<27><1> ), .B(n249), .Y(n1510) );
  OAI21X1 U1104 ( .A(n247), .B(n1410), .C(n1510), .Y(n716) );
  NAND2X1 U1105 ( .A(\mem<27><2> ), .B(n249), .Y(n1511) );
  OAI21X1 U1106 ( .A(n247), .B(n1412), .C(n1511), .Y(n717) );
  NAND2X1 U1107 ( .A(\mem<27><3> ), .B(n249), .Y(n1512) );
  OAI21X1 U1108 ( .A(n247), .B(n1414), .C(n1512), .Y(n718) );
  NAND2X1 U1109 ( .A(\mem<27><4> ), .B(n249), .Y(n1513) );
  OAI21X1 U1110 ( .A(n247), .B(n1416), .C(n1513), .Y(n719) );
  NAND2X1 U1111 ( .A(\mem<27><5> ), .B(n249), .Y(n1514) );
  OAI21X1 U1112 ( .A(n247), .B(n1418), .C(n1514), .Y(n720) );
  NAND2X1 U1113 ( .A(\mem<27><6> ), .B(n249), .Y(n1515) );
  OAI21X1 U1114 ( .A(n247), .B(n1420), .C(n1515), .Y(n721) );
  NAND2X1 U1115 ( .A(\mem<27><7> ), .B(n249), .Y(n1516) );
  OAI21X1 U1116 ( .A(n247), .B(n1422), .C(n1516), .Y(n722) );
  NAND2X1 U1117 ( .A(\mem<27><8> ), .B(n248), .Y(n1517) );
  OAI21X1 U1118 ( .A(n247), .B(n1425), .C(n1517), .Y(n723) );
  NAND2X1 U1119 ( .A(\mem<27><9> ), .B(n248), .Y(n1518) );
  OAI21X1 U1120 ( .A(n247), .B(n1427), .C(n1518), .Y(n724) );
  NAND2X1 U1121 ( .A(\mem<27><10> ), .B(n248), .Y(n1519) );
  OAI21X1 U1122 ( .A(n247), .B(n1429), .C(n1519), .Y(n725) );
  NAND2X1 U1123 ( .A(\mem<27><11> ), .B(n248), .Y(n1520) );
  OAI21X1 U1124 ( .A(n247), .B(n1430), .C(n1520), .Y(n726) );
  NAND2X1 U1125 ( .A(\mem<27><12> ), .B(n248), .Y(n1521) );
  OAI21X1 U1126 ( .A(n247), .B(n1433), .C(n1521), .Y(n727) );
  NAND2X1 U1127 ( .A(\mem<27><13> ), .B(n248), .Y(n1522) );
  OAI21X1 U1128 ( .A(n247), .B(n34), .C(n1522), .Y(n728) );
  NAND2X1 U1129 ( .A(\mem<27><14> ), .B(n248), .Y(n1523) );
  OAI21X1 U1130 ( .A(n247), .B(n24), .C(n1523), .Y(n729) );
  NAND2X1 U1131 ( .A(\mem<27><15> ), .B(n248), .Y(n1524) );
  OAI21X1 U1132 ( .A(n247), .B(n14), .C(n1524), .Y(n730) );
  NAND3X1 U1133 ( .A(n1439), .B(n1436), .C(n1435), .Y(n1525) );
  NAND2X1 U1134 ( .A(\mem<26><0> ), .B(n253), .Y(n1526) );
  OAI21X1 U1135 ( .A(n251), .B(n8), .C(n1526), .Y(n731) );
  NAND2X1 U1136 ( .A(\mem<26><1> ), .B(n253), .Y(n1527) );
  OAI21X1 U1137 ( .A(n251), .B(n1411), .C(n1527), .Y(n732) );
  NAND2X1 U1138 ( .A(\mem<26><2> ), .B(n253), .Y(n1528) );
  OAI21X1 U1139 ( .A(n251), .B(n1413), .C(n1528), .Y(n733) );
  NAND2X1 U1140 ( .A(\mem<26><3> ), .B(n253), .Y(n1529) );
  OAI21X1 U1141 ( .A(n251), .B(n1415), .C(n1529), .Y(n734) );
  NAND2X1 U1142 ( .A(\mem<26><4> ), .B(n253), .Y(n1530) );
  OAI21X1 U1143 ( .A(n251), .B(n1417), .C(n1530), .Y(n735) );
  NAND2X1 U1144 ( .A(\mem<26><5> ), .B(n253), .Y(n1531) );
  OAI21X1 U1145 ( .A(n251), .B(n1419), .C(n1531), .Y(n736) );
  NAND2X1 U1146 ( .A(\mem<26><6> ), .B(n253), .Y(n1532) );
  OAI21X1 U1147 ( .A(n251), .B(n1421), .C(n1532), .Y(n737) );
  NAND2X1 U1148 ( .A(\mem<26><7> ), .B(n253), .Y(n1533) );
  OAI21X1 U1149 ( .A(n251), .B(n1423), .C(n1533), .Y(n738) );
  NAND2X1 U1150 ( .A(\mem<26><8> ), .B(n252), .Y(n1534) );
  OAI21X1 U1151 ( .A(n251), .B(n1424), .C(n1534), .Y(n739) );
  NAND2X1 U1152 ( .A(\mem<26><9> ), .B(n252), .Y(n1535) );
  OAI21X1 U1153 ( .A(n251), .B(n1426), .C(n1535), .Y(n740) );
  NAND2X1 U1154 ( .A(\mem<26><10> ), .B(n252), .Y(n1536) );
  OAI21X1 U1155 ( .A(n251), .B(n1428), .C(n1536), .Y(n741) );
  NAND2X1 U1156 ( .A(\mem<26><11> ), .B(n252), .Y(n1537) );
  OAI21X1 U1157 ( .A(n251), .B(n1431), .C(n1537), .Y(n742) );
  NAND2X1 U1158 ( .A(\mem<26><12> ), .B(n252), .Y(n1538) );
  OAI21X1 U1159 ( .A(n251), .B(n1432), .C(n1538), .Y(n743) );
  NAND2X1 U1160 ( .A(\mem<26><13> ), .B(n252), .Y(n1539) );
  OAI21X1 U1161 ( .A(n251), .B(n42), .C(n1539), .Y(n744) );
  NAND2X1 U1162 ( .A(\mem<26><14> ), .B(n252), .Y(n1540) );
  OAI21X1 U1163 ( .A(n251), .B(n32), .C(n1540), .Y(n745) );
  NAND2X1 U1164 ( .A(\mem<26><15> ), .B(n252), .Y(n1541) );
  OAI21X1 U1165 ( .A(n251), .B(n22), .C(n1541), .Y(n746) );
  NAND3X1 U1166 ( .A(n1352), .B(n1439), .C(n1437), .Y(n1542) );
  NAND2X1 U1167 ( .A(\mem<25><0> ), .B(n257), .Y(n1543) );
  OAI21X1 U1168 ( .A(n255), .B(n7), .C(n1543), .Y(n747) );
  NAND2X1 U1169 ( .A(\mem<25><1> ), .B(n257), .Y(n1544) );
  OAI21X1 U1170 ( .A(n255), .B(n1410), .C(n1544), .Y(n748) );
  NAND2X1 U1171 ( .A(\mem<25><2> ), .B(n257), .Y(n1545) );
  OAI21X1 U1172 ( .A(n255), .B(n1412), .C(n1545), .Y(n749) );
  NAND2X1 U1173 ( .A(\mem<25><3> ), .B(n257), .Y(n1546) );
  OAI21X1 U1174 ( .A(n255), .B(n1414), .C(n1546), .Y(n750) );
  NAND2X1 U1175 ( .A(\mem<25><4> ), .B(n257), .Y(n1547) );
  OAI21X1 U1177 ( .A(n255), .B(n1416), .C(n1547), .Y(n751) );
  NAND2X1 U1178 ( .A(\mem<25><5> ), .B(n257), .Y(n1548) );
  OAI21X1 U1179 ( .A(n255), .B(n1418), .C(n1548), .Y(n752) );
  NAND2X1 U1180 ( .A(\mem<25><6> ), .B(n257), .Y(n1549) );
  OAI21X1 U1181 ( .A(n255), .B(n1420), .C(n1549), .Y(n753) );
  NAND2X1 U1182 ( .A(\mem<25><7> ), .B(n257), .Y(n1550) );
  OAI21X1 U1183 ( .A(n255), .B(n1422), .C(n1550), .Y(n754) );
  NAND2X1 U1184 ( .A(\mem<25><8> ), .B(n256), .Y(n1551) );
  OAI21X1 U1185 ( .A(n255), .B(n1425), .C(n1551), .Y(n755) );
  NAND2X1 U1186 ( .A(\mem<25><9> ), .B(n256), .Y(n1552) );
  OAI21X1 U1187 ( .A(n255), .B(n1427), .C(n1552), .Y(n756) );
  NAND2X1 U1188 ( .A(\mem<25><10> ), .B(n256), .Y(n1553) );
  OAI21X1 U1189 ( .A(n255), .B(n1429), .C(n1553), .Y(n757) );
  NAND2X1 U1190 ( .A(\mem<25><11> ), .B(n256), .Y(n1554) );
  OAI21X1 U1191 ( .A(n255), .B(n1430), .C(n1554), .Y(n758) );
  NAND2X1 U1192 ( .A(\mem<25><12> ), .B(n256), .Y(n1555) );
  OAI21X1 U1193 ( .A(n255), .B(n1433), .C(n1555), .Y(n759) );
  NAND2X1 U1194 ( .A(\mem<25><13> ), .B(n256), .Y(n1556) );
  OAI21X1 U1195 ( .A(n255), .B(n34), .C(n1556), .Y(n760) );
  NAND2X1 U1196 ( .A(\mem<25><14> ), .B(n256), .Y(n1557) );
  OAI21X1 U1197 ( .A(n255), .B(n24), .C(n1557), .Y(n761) );
  NAND2X1 U1198 ( .A(\mem<25><15> ), .B(n256), .Y(n1558) );
  OAI21X1 U1199 ( .A(n255), .B(n14), .C(n1558), .Y(n762) );
  NOR3X1 U1200 ( .A(n1350), .B(n1436), .C(n1438), .Y(n1903) );
  NAND2X1 U1201 ( .A(\mem<24><0> ), .B(n259), .Y(n1559) );
  OAI21X1 U1202 ( .A(n1362), .B(n7), .C(n1559), .Y(n763) );
  NAND2X1 U1203 ( .A(\mem<24><1> ), .B(n259), .Y(n1560) );
  OAI21X1 U1204 ( .A(n1362), .B(n1410), .C(n1560), .Y(n764) );
  NAND2X1 U1205 ( .A(\mem<24><2> ), .B(n259), .Y(n1561) );
  OAI21X1 U1206 ( .A(n1362), .B(n1412), .C(n1561), .Y(n765) );
  NAND2X1 U1207 ( .A(\mem<24><3> ), .B(n259), .Y(n1562) );
  OAI21X1 U1208 ( .A(n1362), .B(n1414), .C(n1562), .Y(n766) );
  NAND2X1 U1209 ( .A(\mem<24><4> ), .B(n259), .Y(n1563) );
  OAI21X1 U1210 ( .A(n1362), .B(n1416), .C(n1563), .Y(n767) );
  NAND2X1 U1211 ( .A(\mem<24><5> ), .B(n259), .Y(n1564) );
  OAI21X1 U1212 ( .A(n1362), .B(n1418), .C(n1564), .Y(n768) );
  NAND2X1 U1213 ( .A(\mem<24><6> ), .B(n259), .Y(n1565) );
  OAI21X1 U1214 ( .A(n1362), .B(n1420), .C(n1565), .Y(n769) );
  NAND2X1 U1215 ( .A(\mem<24><7> ), .B(n259), .Y(n1566) );
  OAI21X1 U1216 ( .A(n1362), .B(n1422), .C(n1566), .Y(n770) );
  NAND2X1 U1217 ( .A(\mem<24><8> ), .B(n258), .Y(n1567) );
  OAI21X1 U1218 ( .A(n1362), .B(n1424), .C(n1567), .Y(n771) );
  NAND2X1 U1219 ( .A(\mem<24><9> ), .B(n258), .Y(n1568) );
  OAI21X1 U1220 ( .A(n1362), .B(n1426), .C(n1568), .Y(n772) );
  NAND2X1 U1221 ( .A(\mem<24><10> ), .B(n258), .Y(n1569) );
  OAI21X1 U1222 ( .A(n1362), .B(n1428), .C(n1569), .Y(n773) );
  NAND2X1 U1223 ( .A(\mem<24><11> ), .B(n258), .Y(n1570) );
  OAI21X1 U1224 ( .A(n1362), .B(n1431), .C(n1570), .Y(n774) );
  NAND2X1 U1225 ( .A(\mem<24><12> ), .B(n258), .Y(n1571) );
  OAI21X1 U1226 ( .A(n1362), .B(n1432), .C(n1571), .Y(n775) );
  NAND2X1 U1227 ( .A(\mem<24><13> ), .B(n258), .Y(n1572) );
  OAI21X1 U1228 ( .A(n1362), .B(n42), .C(n1572), .Y(n776) );
  NAND2X1 U1229 ( .A(\mem<24><14> ), .B(n258), .Y(n1573) );
  OAI21X1 U1230 ( .A(n1362), .B(n32), .C(n1573), .Y(n777) );
  NAND2X1 U1231 ( .A(\mem<24><15> ), .B(n258), .Y(n1574) );
  OAI21X1 U1232 ( .A(n1362), .B(n22), .C(n1574), .Y(n778) );
  NAND2X1 U1233 ( .A(\mem<23><0> ), .B(n263), .Y(n1575) );
  OAI21X1 U1234 ( .A(n261), .B(n6), .C(n1575), .Y(n779) );
  NAND2X1 U1235 ( .A(\mem<23><1> ), .B(n263), .Y(n1576) );
  OAI21X1 U1236 ( .A(n261), .B(n1411), .C(n1576), .Y(n780) );
  NAND2X1 U1237 ( .A(\mem<23><2> ), .B(n263), .Y(n1577) );
  OAI21X1 U1238 ( .A(n261), .B(n1413), .C(n1577), .Y(n781) );
  NAND2X1 U1239 ( .A(\mem<23><3> ), .B(n263), .Y(n1578) );
  OAI21X1 U1240 ( .A(n261), .B(n1415), .C(n1578), .Y(n782) );
  NAND2X1 U1241 ( .A(\mem<23><4> ), .B(n263), .Y(n1579) );
  OAI21X1 U1242 ( .A(n261), .B(n1417), .C(n1579), .Y(n783) );
  NAND2X1 U1243 ( .A(\mem<23><5> ), .B(n263), .Y(n1580) );
  OAI21X1 U1244 ( .A(n261), .B(n1419), .C(n1580), .Y(n784) );
  NAND2X1 U1245 ( .A(\mem<23><6> ), .B(n263), .Y(n1581) );
  OAI21X1 U1246 ( .A(n261), .B(n1421), .C(n1581), .Y(n785) );
  NAND2X1 U1247 ( .A(\mem<23><7> ), .B(n263), .Y(n1582) );
  OAI21X1 U1248 ( .A(n261), .B(n1423), .C(n1582), .Y(n786) );
  NAND2X1 U1249 ( .A(\mem<23><8> ), .B(n262), .Y(n1583) );
  OAI21X1 U1250 ( .A(n261), .B(n1425), .C(n1583), .Y(n787) );
  NAND2X1 U1251 ( .A(\mem<23><9> ), .B(n262), .Y(n1584) );
  OAI21X1 U1252 ( .A(n261), .B(n1427), .C(n1584), .Y(n788) );
  NAND2X1 U1253 ( .A(\mem<23><10> ), .B(n262), .Y(n1585) );
  OAI21X1 U1254 ( .A(n261), .B(n1429), .C(n1585), .Y(n789) );
  NAND2X1 U1255 ( .A(\mem<23><11> ), .B(n262), .Y(n1586) );
  OAI21X1 U1256 ( .A(n261), .B(n1431), .C(n1586), .Y(n790) );
  NAND2X1 U1257 ( .A(\mem<23><12> ), .B(n262), .Y(n1587) );
  OAI21X1 U1258 ( .A(n261), .B(n1433), .C(n1587), .Y(n791) );
  NAND2X1 U1259 ( .A(\mem<23><13> ), .B(n262), .Y(n1588) );
  OAI21X1 U1260 ( .A(n261), .B(n36), .C(n1588), .Y(n792) );
  NAND2X1 U1261 ( .A(\mem<23><14> ), .B(n262), .Y(n1589) );
  OAI21X1 U1262 ( .A(n261), .B(n26), .C(n1589), .Y(n793) );
  NAND2X1 U1263 ( .A(\mem<23><15> ), .B(n262), .Y(n1590) );
  OAI21X1 U1264 ( .A(n261), .B(n16), .C(n1590), .Y(n794) );
  NAND2X1 U1265 ( .A(\mem<22><0> ), .B(n267), .Y(n1591) );
  OAI21X1 U1266 ( .A(n265), .B(n5), .C(n1591), .Y(n795) );
  NAND2X1 U1267 ( .A(\mem<22><1> ), .B(n267), .Y(n1592) );
  OAI21X1 U1268 ( .A(n265), .B(n1411), .C(n1592), .Y(n796) );
  NAND2X1 U1269 ( .A(\mem<22><2> ), .B(n267), .Y(n1593) );
  OAI21X1 U1270 ( .A(n265), .B(n1413), .C(n1593), .Y(n797) );
  NAND2X1 U1271 ( .A(\mem<22><3> ), .B(n267), .Y(n1594) );
  OAI21X1 U1272 ( .A(n265), .B(n1415), .C(n1594), .Y(n798) );
  NAND2X1 U1273 ( .A(\mem<22><4> ), .B(n267), .Y(n1595) );
  OAI21X1 U1274 ( .A(n265), .B(n1417), .C(n1595), .Y(n799) );
  NAND2X1 U1275 ( .A(\mem<22><5> ), .B(n267), .Y(n1596) );
  OAI21X1 U1276 ( .A(n265), .B(n1419), .C(n1596), .Y(n800) );
  NAND2X1 U1277 ( .A(\mem<22><6> ), .B(n267), .Y(n1597) );
  OAI21X1 U1278 ( .A(n265), .B(n1421), .C(n1597), .Y(n801) );
  NAND2X1 U1279 ( .A(\mem<22><7> ), .B(n267), .Y(n1598) );
  OAI21X1 U1280 ( .A(n265), .B(n1423), .C(n1598), .Y(n802) );
  NAND2X1 U1281 ( .A(\mem<22><8> ), .B(n266), .Y(n1599) );
  OAI21X1 U1282 ( .A(n265), .B(n1425), .C(n1599), .Y(n803) );
  NAND2X1 U1283 ( .A(\mem<22><9> ), .B(n266), .Y(n1600) );
  OAI21X1 U1284 ( .A(n265), .B(n1427), .C(n1600), .Y(n804) );
  NAND2X1 U1285 ( .A(\mem<22><10> ), .B(n266), .Y(n1601) );
  OAI21X1 U1286 ( .A(n265), .B(n1429), .C(n1601), .Y(n805) );
  NAND2X1 U1287 ( .A(\mem<22><11> ), .B(n266), .Y(n1602) );
  OAI21X1 U1288 ( .A(n265), .B(n1431), .C(n1602), .Y(n806) );
  NAND2X1 U1289 ( .A(\mem<22><12> ), .B(n266), .Y(n1603) );
  OAI21X1 U1290 ( .A(n265), .B(n1433), .C(n1603), .Y(n807) );
  NAND2X1 U1291 ( .A(\mem<22><13> ), .B(n266), .Y(n1604) );
  OAI21X1 U1292 ( .A(n265), .B(n36), .C(n1604), .Y(n808) );
  NAND2X1 U1293 ( .A(\mem<22><14> ), .B(n266), .Y(n1605) );
  OAI21X1 U1294 ( .A(n265), .B(n27), .C(n1605), .Y(n809) );
  NAND2X1 U1295 ( .A(\mem<22><15> ), .B(n266), .Y(n1606) );
  OAI21X1 U1296 ( .A(n265), .B(n17), .C(n1606), .Y(n810) );
  NAND2X1 U1297 ( .A(\mem<21><0> ), .B(n271), .Y(n1607) );
  OAI21X1 U1298 ( .A(n269), .B(n4), .C(n1607), .Y(n811) );
  NAND2X1 U1299 ( .A(\mem<21><1> ), .B(n271), .Y(n1608) );
  OAI21X1 U1300 ( .A(n269), .B(n1411), .C(n1608), .Y(n812) );
  NAND2X1 U1301 ( .A(\mem<21><2> ), .B(n271), .Y(n1609) );
  OAI21X1 U1302 ( .A(n269), .B(n1413), .C(n1609), .Y(n813) );
  NAND2X1 U1303 ( .A(\mem<21><3> ), .B(n271), .Y(n1610) );
  OAI21X1 U1304 ( .A(n269), .B(n1415), .C(n1610), .Y(n814) );
  NAND2X1 U1305 ( .A(\mem<21><4> ), .B(n271), .Y(n1611) );
  OAI21X1 U1306 ( .A(n269), .B(n1417), .C(n1611), .Y(n815) );
  NAND2X1 U1307 ( .A(\mem<21><5> ), .B(n271), .Y(n1612) );
  OAI21X1 U1308 ( .A(n269), .B(n1419), .C(n1612), .Y(n816) );
  NAND2X1 U1309 ( .A(\mem<21><6> ), .B(n271), .Y(n1613) );
  OAI21X1 U1310 ( .A(n269), .B(n1421), .C(n1613), .Y(n817) );
  NAND2X1 U1311 ( .A(\mem<21><7> ), .B(n271), .Y(n1614) );
  OAI21X1 U1312 ( .A(n269), .B(n1423), .C(n1614), .Y(n818) );
  NAND2X1 U1313 ( .A(\mem<21><8> ), .B(n270), .Y(n1615) );
  OAI21X1 U1314 ( .A(n269), .B(n1425), .C(n1615), .Y(n819) );
  NAND2X1 U1315 ( .A(\mem<21><9> ), .B(n270), .Y(n1616) );
  OAI21X1 U1316 ( .A(n269), .B(n1427), .C(n1616), .Y(n820) );
  NAND2X1 U1317 ( .A(\mem<21><10> ), .B(n270), .Y(n1617) );
  OAI21X1 U1318 ( .A(n269), .B(n1429), .C(n1617), .Y(n821) );
  NAND2X1 U1319 ( .A(\mem<21><11> ), .B(n270), .Y(n1618) );
  OAI21X1 U1320 ( .A(n269), .B(n1431), .C(n1618), .Y(n822) );
  NAND2X1 U1321 ( .A(\mem<21><12> ), .B(n270), .Y(n1619) );
  OAI21X1 U1322 ( .A(n269), .B(n1433), .C(n1619), .Y(n823) );
  NAND2X1 U1323 ( .A(\mem<21><13> ), .B(n270), .Y(n1620) );
  OAI21X1 U1324 ( .A(n269), .B(n37), .C(n1620), .Y(n824) );
  NAND2X1 U1325 ( .A(\mem<21><14> ), .B(n270), .Y(n1621) );
  OAI21X1 U1326 ( .A(n269), .B(n27), .C(n1621), .Y(n825) );
  NAND2X1 U1327 ( .A(\mem<21><15> ), .B(n270), .Y(n1622) );
  OAI21X1 U1328 ( .A(n269), .B(n17), .C(n1622), .Y(n826) );
  NAND2X1 U1329 ( .A(\mem<20><0> ), .B(n275), .Y(n1623) );
  OAI21X1 U1330 ( .A(n273), .B(n13), .C(n1623), .Y(n827) );
  NAND2X1 U1331 ( .A(\mem<20><1> ), .B(n275), .Y(n1624) );
  OAI21X1 U1332 ( .A(n273), .B(n1411), .C(n1624), .Y(n828) );
  NAND2X1 U1333 ( .A(\mem<20><2> ), .B(n275), .Y(n1625) );
  OAI21X1 U1334 ( .A(n273), .B(n1413), .C(n1625), .Y(n829) );
  NAND2X1 U1335 ( .A(\mem<20><3> ), .B(n275), .Y(n1626) );
  OAI21X1 U1336 ( .A(n273), .B(n1415), .C(n1626), .Y(n830) );
  NAND2X1 U1337 ( .A(\mem<20><4> ), .B(n275), .Y(n1627) );
  OAI21X1 U1338 ( .A(n273), .B(n1417), .C(n1627), .Y(n831) );
  NAND2X1 U1339 ( .A(\mem<20><5> ), .B(n275), .Y(n1628) );
  OAI21X1 U1340 ( .A(n273), .B(n1419), .C(n1628), .Y(n832) );
  NAND2X1 U1341 ( .A(\mem<20><6> ), .B(n275), .Y(n1629) );
  OAI21X1 U1342 ( .A(n273), .B(n1421), .C(n1629), .Y(n833) );
  NAND2X1 U1343 ( .A(\mem<20><7> ), .B(n275), .Y(n1630) );
  OAI21X1 U1344 ( .A(n273), .B(n1423), .C(n1630), .Y(n834) );
  NAND2X1 U1345 ( .A(\mem<20><8> ), .B(n274), .Y(n1631) );
  OAI21X1 U1346 ( .A(n273), .B(n1425), .C(n1631), .Y(n835) );
  NAND2X1 U1347 ( .A(\mem<20><9> ), .B(n274), .Y(n1632) );
  OAI21X1 U1348 ( .A(n273), .B(n1427), .C(n1632), .Y(n836) );
  NAND2X1 U1349 ( .A(\mem<20><10> ), .B(n274), .Y(n1633) );
  OAI21X1 U1350 ( .A(n273), .B(n1429), .C(n1633), .Y(n837) );
  NAND2X1 U1351 ( .A(\mem<20><11> ), .B(n274), .Y(n1634) );
  OAI21X1 U1352 ( .A(n273), .B(n1431), .C(n1634), .Y(n838) );
  NAND2X1 U1353 ( .A(\mem<20><12> ), .B(n274), .Y(n1635) );
  OAI21X1 U1354 ( .A(n273), .B(n1433), .C(n1635), .Y(n839) );
  NAND2X1 U1355 ( .A(\mem<20><13> ), .B(n274), .Y(n1636) );
  OAI21X1 U1356 ( .A(n273), .B(n38), .C(n1636), .Y(n840) );
  NAND2X1 U1357 ( .A(\mem<20><14> ), .B(n274), .Y(n1637) );
  OAI21X1 U1358 ( .A(n273), .B(n28), .C(n1637), .Y(n841) );
  NAND2X1 U1359 ( .A(\mem<20><15> ), .B(n274), .Y(n1638) );
  OAI21X1 U1360 ( .A(n273), .B(n18), .C(n1638), .Y(n842) );
  NAND2X1 U1361 ( .A(\mem<19><0> ), .B(n1363), .Y(n1639) );
  OAI21X1 U1362 ( .A(n277), .B(n12), .C(n1639), .Y(n843) );
  NAND2X1 U1363 ( .A(\mem<19><1> ), .B(n1363), .Y(n1640) );
  OAI21X1 U1364 ( .A(n277), .B(n1411), .C(n1640), .Y(n844) );
  NAND2X1 U1365 ( .A(\mem<19><2> ), .B(n1363), .Y(n1641) );
  OAI21X1 U1366 ( .A(n277), .B(n1413), .C(n1641), .Y(n845) );
  NAND2X1 U1367 ( .A(\mem<19><3> ), .B(n1363), .Y(n1642) );
  OAI21X1 U1368 ( .A(n277), .B(n1415), .C(n1642), .Y(n846) );
  NAND2X1 U1369 ( .A(\mem<19><4> ), .B(n1363), .Y(n1643) );
  OAI21X1 U1370 ( .A(n277), .B(n1417), .C(n1643), .Y(n847) );
  NAND2X1 U1371 ( .A(\mem<19><5> ), .B(n1363), .Y(n1644) );
  OAI21X1 U1372 ( .A(n277), .B(n1419), .C(n1644), .Y(n848) );
  NAND2X1 U1373 ( .A(\mem<19><6> ), .B(n1363), .Y(n1645) );
  OAI21X1 U1374 ( .A(n277), .B(n1421), .C(n1645), .Y(n849) );
  NAND2X1 U1375 ( .A(\mem<19><7> ), .B(n1363), .Y(n1646) );
  OAI21X1 U1376 ( .A(n277), .B(n1423), .C(n1646), .Y(n850) );
  NAND2X1 U1377 ( .A(\mem<19><8> ), .B(n1364), .Y(n1647) );
  OAI21X1 U1378 ( .A(n277), .B(n1425), .C(n1647), .Y(n851) );
  NAND2X1 U1379 ( .A(\mem<19><9> ), .B(n1364), .Y(n1648) );
  OAI21X1 U1380 ( .A(n277), .B(n1427), .C(n1648), .Y(n852) );
  NAND2X1 U1381 ( .A(\mem<19><10> ), .B(n1364), .Y(n1649) );
  OAI21X1 U1382 ( .A(n277), .B(n1429), .C(n1649), .Y(n853) );
  NAND2X1 U1383 ( .A(\mem<19><11> ), .B(n1364), .Y(n1650) );
  OAI21X1 U1384 ( .A(n277), .B(n1431), .C(n1650), .Y(n854) );
  NAND2X1 U1385 ( .A(\mem<19><12> ), .B(n1364), .Y(n1651) );
  OAI21X1 U1386 ( .A(n277), .B(n1433), .C(n1651), .Y(n855) );
  NAND2X1 U1387 ( .A(\mem<19><13> ), .B(n1364), .Y(n1652) );
  OAI21X1 U1388 ( .A(n277), .B(n39), .C(n1652), .Y(n856) );
  NAND2X1 U1389 ( .A(\mem<19><14> ), .B(n1364), .Y(n1653) );
  OAI21X1 U1390 ( .A(n277), .B(n29), .C(n1653), .Y(n857) );
  NAND2X1 U1391 ( .A(\mem<19><15> ), .B(n1364), .Y(n1654) );
  OAI21X1 U1392 ( .A(n277), .B(n19), .C(n1654), .Y(n858) );
  NAND2X1 U1393 ( .A(\mem<18><0> ), .B(n1365), .Y(n1655) );
  OAI21X1 U1394 ( .A(n279), .B(n11), .C(n1655), .Y(n859) );
  NAND2X1 U1395 ( .A(\mem<18><1> ), .B(n1365), .Y(n1656) );
  OAI21X1 U1396 ( .A(n279), .B(n1411), .C(n1656), .Y(n860) );
  NAND2X1 U1397 ( .A(\mem<18><2> ), .B(n1365), .Y(n1657) );
  OAI21X1 U1398 ( .A(n279), .B(n1413), .C(n1657), .Y(n861) );
  NAND2X1 U1399 ( .A(\mem<18><3> ), .B(n1365), .Y(n1658) );
  OAI21X1 U1400 ( .A(n279), .B(n1415), .C(n1658), .Y(n862) );
  NAND2X1 U1401 ( .A(\mem<18><4> ), .B(n1365), .Y(n1659) );
  OAI21X1 U1402 ( .A(n279), .B(n1417), .C(n1659), .Y(n863) );
  NAND2X1 U1403 ( .A(\mem<18><5> ), .B(n1365), .Y(n1660) );
  OAI21X1 U1404 ( .A(n279), .B(n1419), .C(n1660), .Y(n864) );
  NAND2X1 U1405 ( .A(\mem<18><6> ), .B(n1365), .Y(n1661) );
  OAI21X1 U1406 ( .A(n279), .B(n1421), .C(n1661), .Y(n865) );
  NAND2X1 U1407 ( .A(\mem<18><7> ), .B(n1365), .Y(n1662) );
  OAI21X1 U1408 ( .A(n279), .B(n1423), .C(n1662), .Y(n866) );
  NAND2X1 U1409 ( .A(\mem<18><8> ), .B(n1366), .Y(n1663) );
  OAI21X1 U1410 ( .A(n279), .B(n1425), .C(n1663), .Y(n867) );
  NAND2X1 U1411 ( .A(\mem<18><9> ), .B(n1366), .Y(n1664) );
  OAI21X1 U1412 ( .A(n279), .B(n1427), .C(n1664), .Y(n868) );
  NAND2X1 U1413 ( .A(\mem<18><10> ), .B(n1366), .Y(n1665) );
  OAI21X1 U1414 ( .A(n279), .B(n1429), .C(n1665), .Y(n869) );
  NAND2X1 U1415 ( .A(\mem<18><11> ), .B(n1366), .Y(n1666) );
  OAI21X1 U1416 ( .A(n279), .B(n1431), .C(n1666), .Y(n870) );
  NAND2X1 U1417 ( .A(\mem<18><12> ), .B(n1366), .Y(n1667) );
  OAI21X1 U1418 ( .A(n279), .B(n1433), .C(n1667), .Y(n871) );
  NAND2X1 U1419 ( .A(\mem<18><13> ), .B(n1366), .Y(n1668) );
  OAI21X1 U1420 ( .A(n279), .B(n40), .C(n1668), .Y(n872) );
  NAND2X1 U1421 ( .A(\mem<18><14> ), .B(n1366), .Y(n1669) );
  OAI21X1 U1422 ( .A(n279), .B(n30), .C(n1669), .Y(n873) );
  NAND2X1 U1423 ( .A(\mem<18><15> ), .B(n1366), .Y(n1670) );
  OAI21X1 U1424 ( .A(n279), .B(n20), .C(n1670), .Y(n874) );
  NAND2X1 U1425 ( .A(\mem<17><0> ), .B(n1367), .Y(n1671) );
  OAI21X1 U1426 ( .A(n281), .B(n10), .C(n1671), .Y(n875) );
  NAND2X1 U1427 ( .A(\mem<17><1> ), .B(n1367), .Y(n1672) );
  OAI21X1 U1428 ( .A(n281), .B(n1411), .C(n1672), .Y(n876) );
  NAND2X1 U1429 ( .A(\mem<17><2> ), .B(n1367), .Y(n1673) );
  OAI21X1 U1430 ( .A(n281), .B(n1413), .C(n1673), .Y(n877) );
  NAND2X1 U1431 ( .A(\mem<17><3> ), .B(n1367), .Y(n1674) );
  OAI21X1 U1432 ( .A(n281), .B(n1415), .C(n1674), .Y(n878) );
  NAND2X1 U1433 ( .A(\mem<17><4> ), .B(n1367), .Y(n1675) );
  OAI21X1 U1434 ( .A(n281), .B(n1417), .C(n1675), .Y(n879) );
  NAND2X1 U1435 ( .A(\mem<17><5> ), .B(n1367), .Y(n1676) );
  OAI21X1 U1436 ( .A(n281), .B(n1419), .C(n1676), .Y(n880) );
  NAND2X1 U1437 ( .A(\mem<17><6> ), .B(n1367), .Y(n1677) );
  OAI21X1 U1438 ( .A(n281), .B(n1421), .C(n1677), .Y(n881) );
  NAND2X1 U1439 ( .A(\mem<17><7> ), .B(n1367), .Y(n1678) );
  OAI21X1 U1440 ( .A(n281), .B(n1423), .C(n1678), .Y(n882) );
  NAND2X1 U1441 ( .A(\mem<17><8> ), .B(n1368), .Y(n1679) );
  OAI21X1 U1442 ( .A(n281), .B(n1425), .C(n1679), .Y(n883) );
  NAND2X1 U1443 ( .A(\mem<17><9> ), .B(n1368), .Y(n1680) );
  OAI21X1 U1444 ( .A(n281), .B(n1427), .C(n1680), .Y(n884) );
  NAND2X1 U1445 ( .A(\mem<17><10> ), .B(n1368), .Y(n1681) );
  OAI21X1 U1446 ( .A(n281), .B(n1429), .C(n1681), .Y(n885) );
  NAND2X1 U1447 ( .A(\mem<17><11> ), .B(n1368), .Y(n1682) );
  OAI21X1 U1448 ( .A(n281), .B(n1431), .C(n1682), .Y(n886) );
  NAND2X1 U1449 ( .A(\mem<17><12> ), .B(n1368), .Y(n1683) );
  OAI21X1 U1450 ( .A(n281), .B(n1433), .C(n1683), .Y(n887) );
  NAND2X1 U1451 ( .A(\mem<17><13> ), .B(n1368), .Y(n1684) );
  OAI21X1 U1452 ( .A(n281), .B(n41), .C(n1684), .Y(n888) );
  NAND2X1 U1453 ( .A(\mem<17><14> ), .B(n1368), .Y(n1685) );
  OAI21X1 U1454 ( .A(n281), .B(n31), .C(n1685), .Y(n889) );
  NAND2X1 U1455 ( .A(\mem<17><15> ), .B(n1368), .Y(n1686) );
  OAI21X1 U1456 ( .A(n281), .B(n21), .C(n1686), .Y(n890) );
  NAND2X1 U1457 ( .A(\mem<16><0> ), .B(n1370), .Y(n1687) );
  OAI21X1 U1458 ( .A(n1369), .B(n6), .C(n1687), .Y(n891) );
  NAND2X1 U1459 ( .A(\mem<16><1> ), .B(n1370), .Y(n1688) );
  OAI21X1 U1460 ( .A(n1369), .B(n1411), .C(n1688), .Y(n892) );
  NAND2X1 U1461 ( .A(\mem<16><2> ), .B(n1370), .Y(n1689) );
  OAI21X1 U1462 ( .A(n1369), .B(n1413), .C(n1689), .Y(n893) );
  NAND2X1 U1463 ( .A(\mem<16><3> ), .B(n1370), .Y(n1690) );
  OAI21X1 U1464 ( .A(n1369), .B(n1415), .C(n1690), .Y(n894) );
  NAND2X1 U1465 ( .A(\mem<16><4> ), .B(n1370), .Y(n1691) );
  OAI21X1 U1466 ( .A(n1369), .B(n1417), .C(n1691), .Y(n895) );
  NAND2X1 U1467 ( .A(\mem<16><5> ), .B(n1370), .Y(n1692) );
  OAI21X1 U1468 ( .A(n1369), .B(n1419), .C(n1692), .Y(n896) );
  NAND2X1 U1469 ( .A(\mem<16><6> ), .B(n1370), .Y(n1693) );
  OAI21X1 U1470 ( .A(n1369), .B(n1421), .C(n1693), .Y(n897) );
  NAND2X1 U1471 ( .A(\mem<16><7> ), .B(n1370), .Y(n1694) );
  OAI21X1 U1472 ( .A(n1369), .B(n1423), .C(n1694), .Y(n898) );
  NAND2X1 U1473 ( .A(\mem<16><8> ), .B(n1371), .Y(n1695) );
  OAI21X1 U1474 ( .A(n1369), .B(n1425), .C(n1695), .Y(n899) );
  NAND2X1 U1475 ( .A(\mem<16><9> ), .B(n1371), .Y(n1696) );
  OAI21X1 U1476 ( .A(n1369), .B(n1427), .C(n1696), .Y(n900) );
  NAND2X1 U1477 ( .A(\mem<16><10> ), .B(n1371), .Y(n1697) );
  OAI21X1 U1478 ( .A(n1369), .B(n1429), .C(n1697), .Y(n901) );
  NAND2X1 U1479 ( .A(\mem<16><11> ), .B(n1371), .Y(n1698) );
  OAI21X1 U1480 ( .A(n1369), .B(n1430), .C(n1698), .Y(n902) );
  NAND2X1 U1481 ( .A(\mem<16><12> ), .B(n1371), .Y(n1699) );
  OAI21X1 U1482 ( .A(n1369), .B(n1433), .C(n1699), .Y(n903) );
  NAND2X1 U1483 ( .A(\mem<16><13> ), .B(n1371), .Y(n1700) );
  OAI21X1 U1484 ( .A(n1369), .B(n39), .C(n1700), .Y(n904) );
  NAND2X1 U1485 ( .A(\mem<16><14> ), .B(n1371), .Y(n1701) );
  OAI21X1 U1486 ( .A(n1369), .B(n28), .C(n1701), .Y(n905) );
  NAND2X1 U1487 ( .A(\mem<16><15> ), .B(n1371), .Y(n1702) );
  OAI21X1 U1488 ( .A(n1369), .B(n19), .C(n1702), .Y(n906) );
  NAND3X1 U1489 ( .A(n1320), .B(n214), .C(n1441), .Y(n1703) );
  NAND2X1 U1490 ( .A(\mem<15><0> ), .B(n1372), .Y(n1704) );
  OAI21X1 U1491 ( .A(n283), .B(n9), .C(n1704), .Y(n907) );
  NAND2X1 U1492 ( .A(\mem<15><1> ), .B(n1372), .Y(n1705) );
  OAI21X1 U1493 ( .A(n283), .B(n1411), .C(n1705), .Y(n908) );
  NAND2X1 U1494 ( .A(\mem<15><2> ), .B(n1372), .Y(n1706) );
  OAI21X1 U1495 ( .A(n283), .B(n1413), .C(n1706), .Y(n909) );
  NAND2X1 U1496 ( .A(\mem<15><3> ), .B(n1372), .Y(n1707) );
  OAI21X1 U1497 ( .A(n283), .B(n1415), .C(n1707), .Y(n910) );
  NAND2X1 U1498 ( .A(\mem<15><4> ), .B(n1372), .Y(n1708) );
  OAI21X1 U1499 ( .A(n283), .B(n1417), .C(n1708), .Y(n911) );
  NAND2X1 U1500 ( .A(\mem<15><5> ), .B(n1372), .Y(n1709) );
  OAI21X1 U1501 ( .A(n283), .B(n1419), .C(n1709), .Y(n912) );
  NAND2X1 U1502 ( .A(\mem<15><6> ), .B(n1372), .Y(n1710) );
  OAI21X1 U1503 ( .A(n283), .B(n1421), .C(n1710), .Y(n913) );
  NAND2X1 U1504 ( .A(\mem<15><7> ), .B(n1372), .Y(n1711) );
  OAI21X1 U1505 ( .A(n283), .B(n1423), .C(n1711), .Y(n914) );
  NAND2X1 U1506 ( .A(\mem<15><8> ), .B(n1373), .Y(n1712) );
  OAI21X1 U1507 ( .A(n283), .B(n1425), .C(n1712), .Y(n915) );
  NAND2X1 U1508 ( .A(\mem<15><9> ), .B(n1373), .Y(n1713) );
  OAI21X1 U1509 ( .A(n283), .B(n1427), .C(n1713), .Y(n916) );
  NAND2X1 U1510 ( .A(\mem<15><10> ), .B(n1373), .Y(n1714) );
  OAI21X1 U1511 ( .A(n283), .B(n1429), .C(n1714), .Y(n917) );
  NAND2X1 U1512 ( .A(\mem<15><11> ), .B(n1373), .Y(n1715) );
  OAI21X1 U1513 ( .A(n283), .B(n1431), .C(n1715), .Y(n918) );
  NAND2X1 U1514 ( .A(\mem<15><12> ), .B(n1373), .Y(n1716) );
  OAI21X1 U1515 ( .A(n283), .B(n1433), .C(n1716), .Y(n919) );
  NAND2X1 U1516 ( .A(\mem<15><13> ), .B(n1373), .Y(n1717) );
  OAI21X1 U1517 ( .A(n283), .B(n37), .C(n1717), .Y(n920) );
  NAND2X1 U1518 ( .A(\mem<15><14> ), .B(n1373), .Y(n1718) );
  OAI21X1 U1519 ( .A(n283), .B(n26), .C(n1718), .Y(n921) );
  NAND2X1 U1520 ( .A(\mem<15><15> ), .B(n1373), .Y(n1719) );
  OAI21X1 U1521 ( .A(n283), .B(n16), .C(n1719), .Y(n922) );
  NAND2X1 U1522 ( .A(\mem<14><0> ), .B(n1374), .Y(n1720) );
  OAI21X1 U1523 ( .A(n285), .B(n6), .C(n1720), .Y(n923) );
  NAND2X1 U1524 ( .A(\mem<14><1> ), .B(n1374), .Y(n1721) );
  OAI21X1 U1525 ( .A(n285), .B(n1411), .C(n1721), .Y(n924) );
  NAND2X1 U1526 ( .A(\mem<14><2> ), .B(n1374), .Y(n1722) );
  OAI21X1 U1527 ( .A(n285), .B(n1413), .C(n1722), .Y(n925) );
  NAND2X1 U1528 ( .A(\mem<14><3> ), .B(n1374), .Y(n1723) );
  OAI21X1 U1529 ( .A(n285), .B(n1415), .C(n1723), .Y(n926) );
  NAND2X1 U1530 ( .A(\mem<14><4> ), .B(n1374), .Y(n1724) );
  OAI21X1 U1531 ( .A(n285), .B(n1417), .C(n1724), .Y(n927) );
  NAND2X1 U1532 ( .A(\mem<14><5> ), .B(n1374), .Y(n1725) );
  OAI21X1 U1533 ( .A(n285), .B(n1419), .C(n1725), .Y(n928) );
  NAND2X1 U1534 ( .A(\mem<14><6> ), .B(n1374), .Y(n1726) );
  OAI21X1 U1535 ( .A(n285), .B(n1421), .C(n1726), .Y(n929) );
  NAND2X1 U1536 ( .A(\mem<14><7> ), .B(n1374), .Y(n1727) );
  OAI21X1 U1537 ( .A(n285), .B(n1423), .C(n1727), .Y(n930) );
  NAND2X1 U1538 ( .A(\mem<14><8> ), .B(n1375), .Y(n1728) );
  OAI21X1 U1539 ( .A(n285), .B(n1425), .C(n1728), .Y(n931) );
  NAND2X1 U1540 ( .A(\mem<14><9> ), .B(n1375), .Y(n1729) );
  OAI21X1 U1541 ( .A(n285), .B(n1427), .C(n1729), .Y(n932) );
  NAND2X1 U1542 ( .A(\mem<14><10> ), .B(n1375), .Y(n1730) );
  OAI21X1 U1543 ( .A(n285), .B(n1429), .C(n1730), .Y(n933) );
  NAND2X1 U1544 ( .A(\mem<14><11> ), .B(n1375), .Y(n1731) );
  OAI21X1 U1545 ( .A(n285), .B(n1431), .C(n1731), .Y(n934) );
  NAND2X1 U1546 ( .A(\mem<14><12> ), .B(n1375), .Y(n1732) );
  OAI21X1 U1547 ( .A(n285), .B(n1433), .C(n1732), .Y(n935) );
  NAND2X1 U1548 ( .A(\mem<14><13> ), .B(n1375), .Y(n1733) );
  OAI21X1 U1549 ( .A(n285), .B(n36), .C(n1733), .Y(n936) );
  NAND2X1 U1550 ( .A(\mem<14><14> ), .B(n1375), .Y(n1734) );
  OAI21X1 U1551 ( .A(n285), .B(n29), .C(n1734), .Y(n937) );
  NAND2X1 U1552 ( .A(\mem<14><15> ), .B(n1375), .Y(n1735) );
  OAI21X1 U1553 ( .A(n285), .B(n16), .C(n1735), .Y(n938) );
  NAND2X1 U1554 ( .A(\mem<13><0> ), .B(n1376), .Y(n1736) );
  OAI21X1 U1555 ( .A(n287), .B(n5), .C(n1736), .Y(n939) );
  NAND2X1 U1556 ( .A(\mem<13><1> ), .B(n1376), .Y(n1737) );
  OAI21X1 U1557 ( .A(n287), .B(n1411), .C(n1737), .Y(n940) );
  NAND2X1 U1558 ( .A(\mem<13><2> ), .B(n1376), .Y(n1738) );
  OAI21X1 U1559 ( .A(n287), .B(n1413), .C(n1738), .Y(n941) );
  NAND2X1 U1560 ( .A(\mem<13><3> ), .B(n1376), .Y(n1739) );
  OAI21X1 U1561 ( .A(n287), .B(n1415), .C(n1739), .Y(n942) );
  NAND2X1 U1562 ( .A(\mem<13><4> ), .B(n1376), .Y(n1740) );
  OAI21X1 U1563 ( .A(n287), .B(n1417), .C(n1740), .Y(n943) );
  NAND2X1 U1564 ( .A(\mem<13><5> ), .B(n1376), .Y(n1741) );
  OAI21X1 U1565 ( .A(n287), .B(n1419), .C(n1741), .Y(n944) );
  NAND2X1 U1566 ( .A(\mem<13><6> ), .B(n1376), .Y(n1742) );
  OAI21X1 U1567 ( .A(n287), .B(n1421), .C(n1742), .Y(n945) );
  NAND2X1 U1568 ( .A(\mem<13><7> ), .B(n1376), .Y(n1743) );
  OAI21X1 U1569 ( .A(n287), .B(n1423), .C(n1743), .Y(n946) );
  NAND2X1 U1570 ( .A(\mem<13><8> ), .B(n1377), .Y(n1744) );
  OAI21X1 U1571 ( .A(n287), .B(n1425), .C(n1744), .Y(n947) );
  NAND2X1 U1572 ( .A(\mem<13><9> ), .B(n1377), .Y(n1745) );
  OAI21X1 U1573 ( .A(n287), .B(n1427), .C(n1745), .Y(n948) );
  NAND2X1 U1574 ( .A(\mem<13><10> ), .B(n1377), .Y(n1746) );
  OAI21X1 U1575 ( .A(n287), .B(n1429), .C(n1746), .Y(n949) );
  NAND2X1 U1576 ( .A(\mem<13><11> ), .B(n1377), .Y(n1747) );
  OAI21X1 U1577 ( .A(n287), .B(n1431), .C(n1747), .Y(n950) );
  NAND2X1 U1578 ( .A(\mem<13><12> ), .B(n1377), .Y(n1748) );
  OAI21X1 U1579 ( .A(n287), .B(n1433), .C(n1748), .Y(n951) );
  NAND2X1 U1580 ( .A(\mem<13><13> ), .B(n1377), .Y(n1749) );
  OAI21X1 U1581 ( .A(n287), .B(n39), .C(n1749), .Y(n952) );
  NAND2X1 U1582 ( .A(\mem<13><14> ), .B(n1377), .Y(n1750) );
  OAI21X1 U1583 ( .A(n287), .B(n31), .C(n1750), .Y(n953) );
  NAND2X1 U1584 ( .A(\mem<13><15> ), .B(n1377), .Y(n1751) );
  OAI21X1 U1585 ( .A(n287), .B(n19), .C(n1751), .Y(n954) );
  NAND2X1 U1586 ( .A(\mem<12><0> ), .B(n1378), .Y(n1752) );
  OAI21X1 U1587 ( .A(n289), .B(n4), .C(n1752), .Y(n955) );
  NAND2X1 U1588 ( .A(\mem<12><1> ), .B(n1378), .Y(n1753) );
  OAI21X1 U1589 ( .A(n289), .B(n1411), .C(n1753), .Y(n956) );
  NAND2X1 U1590 ( .A(\mem<12><2> ), .B(n1378), .Y(n1754) );
  OAI21X1 U1591 ( .A(n289), .B(n1413), .C(n1754), .Y(n957) );
  NAND2X1 U1592 ( .A(\mem<12><3> ), .B(n1378), .Y(n1755) );
  OAI21X1 U1593 ( .A(n289), .B(n1415), .C(n1755), .Y(n958) );
  NAND2X1 U1594 ( .A(\mem<12><4> ), .B(n1378), .Y(n1756) );
  OAI21X1 U1595 ( .A(n289), .B(n1417), .C(n1756), .Y(n959) );
  NAND2X1 U1596 ( .A(\mem<12><5> ), .B(n1378), .Y(n1757) );
  OAI21X1 U1597 ( .A(n289), .B(n1419), .C(n1757), .Y(n960) );
  NAND2X1 U1598 ( .A(\mem<12><6> ), .B(n1378), .Y(n1758) );
  OAI21X1 U1599 ( .A(n289), .B(n1421), .C(n1758), .Y(n961) );
  NAND2X1 U1600 ( .A(\mem<12><7> ), .B(n1378), .Y(n1759) );
  OAI21X1 U1601 ( .A(n289), .B(n1423), .C(n1759), .Y(n962) );
  NAND2X1 U1602 ( .A(\mem<12><8> ), .B(n1379), .Y(n1760) );
  OAI21X1 U1603 ( .A(n289), .B(n1425), .C(n1760), .Y(n963) );
  NAND2X1 U1604 ( .A(\mem<12><9> ), .B(n1379), .Y(n1761) );
  OAI21X1 U1605 ( .A(n289), .B(n1427), .C(n1761), .Y(n964) );
  NAND2X1 U1606 ( .A(\mem<12><10> ), .B(n1379), .Y(n1762) );
  OAI21X1 U1607 ( .A(n289), .B(n1429), .C(n1762), .Y(n965) );
  NAND2X1 U1608 ( .A(\mem<12><11> ), .B(n1379), .Y(n1763) );
  OAI21X1 U1609 ( .A(n289), .B(n1431), .C(n1763), .Y(n966) );
  NAND2X1 U1610 ( .A(\mem<12><12> ), .B(n1379), .Y(n1764) );
  OAI21X1 U1611 ( .A(n289), .B(n1433), .C(n1764), .Y(n967) );
  NAND2X1 U1612 ( .A(\mem<12><13> ), .B(n1379), .Y(n1765) );
  OAI21X1 U1613 ( .A(n289), .B(n41), .C(n1765), .Y(n968) );
  NAND2X1 U1614 ( .A(\mem<12><14> ), .B(n1379), .Y(n1766) );
  OAI21X1 U1615 ( .A(n289), .B(n29), .C(n1766), .Y(n969) );
  NAND2X1 U1616 ( .A(\mem<12><15> ), .B(n1379), .Y(n1767) );
  OAI21X1 U1617 ( .A(n289), .B(n21), .C(n1767), .Y(n970) );
  NAND2X1 U1618 ( .A(\mem<11><0> ), .B(n1380), .Y(n1768) );
  OAI21X1 U1619 ( .A(n291), .B(n9), .C(n1768), .Y(n971) );
  NAND2X1 U1620 ( .A(\mem<11><1> ), .B(n1380), .Y(n1769) );
  OAI21X1 U1621 ( .A(n291), .B(n1410), .C(n1769), .Y(n972) );
  NAND2X1 U1622 ( .A(\mem<11><2> ), .B(n1380), .Y(n1770) );
  OAI21X1 U1623 ( .A(n291), .B(n1412), .C(n1770), .Y(n973) );
  NAND2X1 U1624 ( .A(\mem<11><3> ), .B(n1380), .Y(n1771) );
  OAI21X1 U1625 ( .A(n291), .B(n1414), .C(n1771), .Y(n974) );
  NAND2X1 U1626 ( .A(\mem<11><4> ), .B(n1380), .Y(n1772) );
  OAI21X1 U1627 ( .A(n291), .B(n1416), .C(n1772), .Y(n975) );
  NAND2X1 U1628 ( .A(\mem<11><5> ), .B(n1380), .Y(n1773) );
  OAI21X1 U1629 ( .A(n291), .B(n1418), .C(n1773), .Y(n976) );
  NAND2X1 U1630 ( .A(\mem<11><6> ), .B(n1380), .Y(n1774) );
  OAI21X1 U1631 ( .A(n291), .B(n1420), .C(n1774), .Y(n977) );
  NAND2X1 U1632 ( .A(\mem<11><7> ), .B(n1380), .Y(n1775) );
  OAI21X1 U1633 ( .A(n291), .B(n1422), .C(n1775), .Y(n978) );
  NAND2X1 U1634 ( .A(\mem<11><8> ), .B(n1381), .Y(n1776) );
  OAI21X1 U1635 ( .A(n291), .B(n1424), .C(n1776), .Y(n979) );
  NAND2X1 U1636 ( .A(\mem<11><9> ), .B(n1381), .Y(n1777) );
  OAI21X1 U1637 ( .A(n291), .B(n1426), .C(n1777), .Y(n980) );
  NAND2X1 U1638 ( .A(\mem<11><10> ), .B(n1381), .Y(n1778) );
  OAI21X1 U1639 ( .A(n291), .B(n1428), .C(n1778), .Y(n981) );
  NAND2X1 U1640 ( .A(\mem<11><11> ), .B(n1381), .Y(n1779) );
  OAI21X1 U1641 ( .A(n291), .B(n1430), .C(n1779), .Y(n982) );
  NAND2X1 U1642 ( .A(\mem<11><12> ), .B(n1381), .Y(n1780) );
  OAI21X1 U1643 ( .A(n291), .B(n1432), .C(n1780), .Y(n983) );
  NAND2X1 U1644 ( .A(\mem<11><13> ), .B(n1381), .Y(n1781) );
  OAI21X1 U1645 ( .A(n291), .B(n40), .C(n1781), .Y(n984) );
  NAND2X1 U1646 ( .A(\mem<11><14> ), .B(n1381), .Y(n1782) );
  OAI21X1 U1647 ( .A(n291), .B(n24), .C(n1782), .Y(n985) );
  NAND2X1 U1648 ( .A(\mem<11><15> ), .B(n1381), .Y(n1783) );
  OAI21X1 U1649 ( .A(n291), .B(n20), .C(n1783), .Y(n986) );
  NAND2X1 U1650 ( .A(\mem<10><0> ), .B(n1382), .Y(n1784) );
  OAI21X1 U1651 ( .A(n293), .B(n4), .C(n1784), .Y(n987) );
  NAND2X1 U1652 ( .A(\mem<10><1> ), .B(n1382), .Y(n1785) );
  OAI21X1 U1653 ( .A(n293), .B(n1410), .C(n1785), .Y(n988) );
  NAND2X1 U1654 ( .A(\mem<10><2> ), .B(n1382), .Y(n1786) );
  OAI21X1 U1655 ( .A(n293), .B(n1412), .C(n1786), .Y(n989) );
  NAND2X1 U1656 ( .A(\mem<10><3> ), .B(n1382), .Y(n1787) );
  OAI21X1 U1657 ( .A(n293), .B(n1414), .C(n1787), .Y(n990) );
  NAND2X1 U1658 ( .A(\mem<10><4> ), .B(n1382), .Y(n1788) );
  OAI21X1 U1659 ( .A(n293), .B(n1416), .C(n1788), .Y(n991) );
  NAND2X1 U1660 ( .A(\mem<10><5> ), .B(n1382), .Y(n1789) );
  OAI21X1 U1661 ( .A(n293), .B(n1418), .C(n1789), .Y(n992) );
  NAND2X1 U1662 ( .A(\mem<10><6> ), .B(n1382), .Y(n1790) );
  OAI21X1 U1663 ( .A(n293), .B(n1420), .C(n1790), .Y(n993) );
  NAND2X1 U1664 ( .A(\mem<10><7> ), .B(n1382), .Y(n1791) );
  OAI21X1 U1665 ( .A(n293), .B(n1422), .C(n1791), .Y(n994) );
  NAND2X1 U1666 ( .A(\mem<10><8> ), .B(n1383), .Y(n1792) );
  OAI21X1 U1667 ( .A(n293), .B(n1424), .C(n1792), .Y(n995) );
  NAND2X1 U1668 ( .A(\mem<10><9> ), .B(n1383), .Y(n1793) );
  OAI21X1 U1669 ( .A(n293), .B(n1426), .C(n1793), .Y(n996) );
  NAND2X1 U1670 ( .A(\mem<10><10> ), .B(n1383), .Y(n1794) );
  OAI21X1 U1671 ( .A(n293), .B(n1428), .C(n1794), .Y(n997) );
  NAND2X1 U1672 ( .A(\mem<10><11> ), .B(n1383), .Y(n1795) );
  OAI21X1 U1673 ( .A(n293), .B(n1430), .C(n1795), .Y(n998) );
  NAND2X1 U1674 ( .A(\mem<10><12> ), .B(n1383), .Y(n1796) );
  OAI21X1 U1675 ( .A(n293), .B(n1432), .C(n1796), .Y(n999) );
  NAND2X1 U1676 ( .A(\mem<10><13> ), .B(n1383), .Y(n1797) );
  OAI21X1 U1677 ( .A(n293), .B(n34), .C(n1797), .Y(n1000) );
  NAND2X1 U1678 ( .A(\mem<10><14> ), .B(n1383), .Y(n1798) );
  OAI21X1 U1679 ( .A(n293), .B(n32), .C(n1798), .Y(n1001) );
  NAND2X1 U1680 ( .A(\mem<10><15> ), .B(n1383), .Y(n1799) );
  OAI21X1 U1681 ( .A(n293), .B(n14), .C(n1799), .Y(n1002) );
  NAND2X1 U1682 ( .A(\mem<9><0> ), .B(n1384), .Y(n1800) );
  OAI21X1 U1683 ( .A(n295), .B(n8), .C(n1800), .Y(n1003) );
  NAND2X1 U1684 ( .A(\mem<9><1> ), .B(n1384), .Y(n1801) );
  OAI21X1 U1685 ( .A(n295), .B(n1410), .C(n1801), .Y(n1004) );
  NAND2X1 U1686 ( .A(\mem<9><2> ), .B(n1384), .Y(n1802) );
  OAI21X1 U1687 ( .A(n295), .B(n1412), .C(n1802), .Y(n1005) );
  NAND2X1 U1688 ( .A(\mem<9><3> ), .B(n1384), .Y(n1803) );
  OAI21X1 U1689 ( .A(n295), .B(n1414), .C(n1803), .Y(n1006) );
  NAND2X1 U1690 ( .A(\mem<9><4> ), .B(n1384), .Y(n1804) );
  OAI21X1 U1691 ( .A(n295), .B(n1416), .C(n1804), .Y(n1007) );
  NAND2X1 U1692 ( .A(\mem<9><5> ), .B(n1384), .Y(n1805) );
  OAI21X1 U1693 ( .A(n295), .B(n1418), .C(n1805), .Y(n1008) );
  NAND2X1 U1694 ( .A(\mem<9><6> ), .B(n1384), .Y(n1806) );
  OAI21X1 U1695 ( .A(n295), .B(n1420), .C(n1806), .Y(n1009) );
  NAND2X1 U1696 ( .A(\mem<9><7> ), .B(n1384), .Y(n1807) );
  OAI21X1 U1697 ( .A(n295), .B(n1422), .C(n1807), .Y(n1010) );
  NAND2X1 U1698 ( .A(\mem<9><8> ), .B(n1385), .Y(n1808) );
  OAI21X1 U1699 ( .A(n295), .B(n1424), .C(n1808), .Y(n1011) );
  NAND2X1 U1700 ( .A(\mem<9><9> ), .B(n1385), .Y(n1809) );
  OAI21X1 U1701 ( .A(n295), .B(n1426), .C(n1809), .Y(n1012) );
  NAND2X1 U1702 ( .A(\mem<9><10> ), .B(n1385), .Y(n1810) );
  OAI21X1 U1703 ( .A(n295), .B(n1428), .C(n1810), .Y(n1013) );
  NAND2X1 U1704 ( .A(\mem<9><11> ), .B(n1385), .Y(n1811) );
  OAI21X1 U1705 ( .A(n295), .B(n1430), .C(n1811), .Y(n1014) );
  NAND2X1 U1706 ( .A(\mem<9><12> ), .B(n1385), .Y(n1812) );
  OAI21X1 U1707 ( .A(n295), .B(n1432), .C(n1812), .Y(n1015) );
  NAND2X1 U1708 ( .A(\mem<9><13> ), .B(n1385), .Y(n1813) );
  OAI21X1 U1709 ( .A(n295), .B(n42), .C(n1813), .Y(n1016) );
  NAND2X1 U1710 ( .A(\mem<9><14> ), .B(n1385), .Y(n1814) );
  OAI21X1 U1711 ( .A(n295), .B(n33), .C(n1814), .Y(n1017) );
  NAND2X1 U1712 ( .A(\mem<9><15> ), .B(n1385), .Y(n1815) );
  OAI21X1 U1713 ( .A(n295), .B(n22), .C(n1815), .Y(n1018) );
  NAND2X1 U1714 ( .A(\mem<8><0> ), .B(n1387), .Y(n1817) );
  OAI21X1 U1715 ( .A(n1386), .B(n5), .C(n1817), .Y(n1019) );
  NAND2X1 U1716 ( .A(\mem<8><1> ), .B(n1387), .Y(n1818) );
  OAI21X1 U1717 ( .A(n1386), .B(n1410), .C(n1818), .Y(n1020) );
  NAND2X1 U1718 ( .A(\mem<8><2> ), .B(n1387), .Y(n1819) );
  OAI21X1 U1719 ( .A(n1386), .B(n1412), .C(n1819), .Y(n1021) );
  NAND2X1 U1720 ( .A(\mem<8><3> ), .B(n1387), .Y(n1820) );
  OAI21X1 U1721 ( .A(n1386), .B(n1414), .C(n1820), .Y(n1022) );
  NAND2X1 U1722 ( .A(\mem<8><4> ), .B(n1387), .Y(n1821) );
  OAI21X1 U1723 ( .A(n1386), .B(n1416), .C(n1821), .Y(n1023) );
  NAND2X1 U1724 ( .A(\mem<8><5> ), .B(n1387), .Y(n1822) );
  OAI21X1 U1725 ( .A(n1386), .B(n1418), .C(n1822), .Y(n1024) );
  NAND2X1 U1726 ( .A(\mem<8><6> ), .B(n1387), .Y(n1823) );
  OAI21X1 U1727 ( .A(n1386), .B(n1420), .C(n1823), .Y(n1025) );
  NAND2X1 U1728 ( .A(\mem<8><7> ), .B(n1387), .Y(n1824) );
  OAI21X1 U1729 ( .A(n1386), .B(n1422), .C(n1824), .Y(n1026) );
  NAND2X1 U1730 ( .A(\mem<8><8> ), .B(n1388), .Y(n1825) );
  OAI21X1 U1731 ( .A(n1386), .B(n1424), .C(n1825), .Y(n1027) );
  NAND2X1 U1732 ( .A(\mem<8><9> ), .B(n1388), .Y(n1826) );
  OAI21X1 U1733 ( .A(n1386), .B(n1426), .C(n1826), .Y(n1028) );
  NAND2X1 U1734 ( .A(\mem<8><10> ), .B(n1388), .Y(n1827) );
  OAI21X1 U1735 ( .A(n1386), .B(n1428), .C(n1827), .Y(n1029) );
  NAND2X1 U1736 ( .A(\mem<8><11> ), .B(n1388), .Y(n1828) );
  OAI21X1 U1737 ( .A(n1386), .B(n1430), .C(n1828), .Y(n1030) );
  NAND2X1 U1738 ( .A(\mem<8><12> ), .B(n1388), .Y(n1829) );
  OAI21X1 U1739 ( .A(n1386), .B(n1432), .C(n1829), .Y(n1031) );
  NAND2X1 U1740 ( .A(\mem<8><13> ), .B(n1388), .Y(n1830) );
  OAI21X1 U1741 ( .A(n1386), .B(n38), .C(n1830), .Y(n1032) );
  NAND2X1 U1742 ( .A(\mem<8><14> ), .B(n1388), .Y(n1831) );
  OAI21X1 U1743 ( .A(n1386), .B(n28), .C(n1831), .Y(n1033) );
  NAND2X1 U1744 ( .A(\mem<8><15> ), .B(n1388), .Y(n1832) );
  OAI21X1 U1745 ( .A(n1386), .B(n18), .C(n1832), .Y(n1034) );
  NAND3X1 U1746 ( .A(n1440), .B(n214), .C(n1441), .Y(n1833) );
  NAND2X1 U1747 ( .A(\mem<7><0> ), .B(n1389), .Y(n1834) );
  OAI21X1 U1748 ( .A(n297), .B(n13), .C(n1834), .Y(n1035) );
  OAI21X1 U1749 ( .A(n297), .B(n1410), .C(n45), .Y(n1036) );
  OAI21X1 U1750 ( .A(n297), .B(n1412), .C(n47), .Y(n1037) );
  OAI21X1 U1751 ( .A(n297), .B(n1414), .C(n49), .Y(n1038) );
  OAI21X1 U1752 ( .A(n297), .B(n1416), .C(n51), .Y(n1039) );
  OAI21X1 U1753 ( .A(n297), .B(n1418), .C(n53), .Y(n1040) );
  OAI21X1 U1754 ( .A(n297), .B(n1420), .C(n55), .Y(n1041) );
  OAI21X1 U1755 ( .A(n297), .B(n1422), .C(n57), .Y(n1042) );
  NAND2X1 U1756 ( .A(\mem<7><8> ), .B(n1390), .Y(n1835) );
  OAI21X1 U1757 ( .A(n297), .B(n1424), .C(n1835), .Y(n1043) );
  NAND2X1 U1758 ( .A(\mem<7><9> ), .B(n1390), .Y(n1836) );
  OAI21X1 U1759 ( .A(n297), .B(n1426), .C(n1836), .Y(n1044) );
  NAND2X1 U1760 ( .A(\mem<7><10> ), .B(n1390), .Y(n1837) );
  OAI21X1 U1761 ( .A(n297), .B(n1428), .C(n1837), .Y(n1045) );
  NAND2X1 U1762 ( .A(\mem<7><11> ), .B(n1390), .Y(n1838) );
  OAI21X1 U1763 ( .A(n297), .B(n1431), .C(n1838), .Y(n1046) );
  NAND2X1 U1764 ( .A(\mem<7><12> ), .B(n1390), .Y(n1839) );
  OAI21X1 U1765 ( .A(n297), .B(n1432), .C(n1839), .Y(n1047) );
  NAND2X1 U1766 ( .A(\mem<7><13> ), .B(n1390), .Y(n1840) );
  OAI21X1 U1767 ( .A(n297), .B(n43), .C(n1840), .Y(n1048) );
  NAND2X1 U1768 ( .A(\mem<7><14> ), .B(n1390), .Y(n1841) );
  OAI21X1 U1769 ( .A(n297), .B(n26), .C(n1841), .Y(n1049) );
  NAND2X1 U1770 ( .A(\mem<7><15> ), .B(n1390), .Y(n1842) );
  OAI21X1 U1771 ( .A(n297), .B(n23), .C(n1842), .Y(n1050) );
  NAND2X1 U1772 ( .A(\mem<6><0> ), .B(n1391), .Y(n1843) );
  OAI21X1 U1773 ( .A(n299), .B(n12), .C(n1843), .Y(n1051) );
  OAI21X1 U1774 ( .A(n299), .B(n1410), .C(n59), .Y(n1052) );
  OAI21X1 U1775 ( .A(n299), .B(n1412), .C(n61), .Y(n1053) );
  OAI21X1 U1776 ( .A(n299), .B(n1414), .C(n63), .Y(n1054) );
  OAI21X1 U1777 ( .A(n299), .B(n1416), .C(n65), .Y(n1055) );
  OAI21X1 U1778 ( .A(n299), .B(n1418), .C(n67), .Y(n1056) );
  OAI21X1 U1779 ( .A(n299), .B(n1420), .C(n69), .Y(n1057) );
  OAI21X1 U1780 ( .A(n299), .B(n1422), .C(n71), .Y(n1058) );
  NAND2X1 U1781 ( .A(\mem<6><8> ), .B(n1392), .Y(n1844) );
  OAI21X1 U1782 ( .A(n299), .B(n1424), .C(n1844), .Y(n1059) );
  NAND2X1 U1783 ( .A(\mem<6><9> ), .B(n1392), .Y(n1845) );
  OAI21X1 U1784 ( .A(n299), .B(n1426), .C(n1845), .Y(n1060) );
  NAND2X1 U1785 ( .A(\mem<6><10> ), .B(n1392), .Y(n1846) );
  OAI21X1 U1786 ( .A(n299), .B(n1428), .C(n1846), .Y(n1061) );
  NAND2X1 U1787 ( .A(\mem<6><11> ), .B(n1392), .Y(n1847) );
  OAI21X1 U1788 ( .A(n299), .B(n1430), .C(n1847), .Y(n1062) );
  NAND2X1 U1789 ( .A(\mem<6><12> ), .B(n1392), .Y(n1848) );
  OAI21X1 U1790 ( .A(n299), .B(n1432), .C(n1848), .Y(n1063) );
  NAND2X1 U1791 ( .A(\mem<6><13> ), .B(n1392), .Y(n1849) );
  OAI21X1 U1792 ( .A(n299), .B(n34), .C(n1849), .Y(n1064) );
  NAND2X1 U1793 ( .A(\mem<6><14> ), .B(n1392), .Y(n1850) );
  OAI21X1 U1794 ( .A(n299), .B(n26), .C(n1850), .Y(n1065) );
  NAND2X1 U1795 ( .A(\mem<6><15> ), .B(n1392), .Y(n1851) );
  OAI21X1 U1796 ( .A(n299), .B(n16), .C(n1851), .Y(n1066) );
  NAND2X1 U1797 ( .A(\mem<5><0> ), .B(n1393), .Y(n1853) );
  OAI21X1 U1798 ( .A(n301), .B(n11), .C(n1853), .Y(n1067) );
  OAI21X1 U1799 ( .A(n301), .B(n1410), .C(n73), .Y(n1068) );
  OAI21X1 U1800 ( .A(n301), .B(n1412), .C(n75), .Y(n1069) );
  OAI21X1 U1801 ( .A(n301), .B(n1414), .C(n77), .Y(n1070) );
  OAI21X1 U1802 ( .A(n301), .B(n1416), .C(n79), .Y(n1071) );
  OAI21X1 U1803 ( .A(n301), .B(n1418), .C(n81), .Y(n1072) );
  OAI21X1 U1804 ( .A(n301), .B(n1420), .C(n83), .Y(n1073) );
  OAI21X1 U1805 ( .A(n301), .B(n1422), .C(n85), .Y(n1074) );
  NAND2X1 U1806 ( .A(\mem<5><8> ), .B(n1394), .Y(n1854) );
  OAI21X1 U1807 ( .A(n301), .B(n1424), .C(n1854), .Y(n1075) );
  NAND2X1 U1808 ( .A(\mem<5><9> ), .B(n1394), .Y(n1855) );
  OAI21X1 U1809 ( .A(n301), .B(n1426), .C(n1855), .Y(n1076) );
  NAND2X1 U1810 ( .A(\mem<5><10> ), .B(n1394), .Y(n1856) );
  OAI21X1 U1811 ( .A(n301), .B(n1428), .C(n1856), .Y(n1077) );
  NAND2X1 U1812 ( .A(\mem<5><11> ), .B(n1394), .Y(n1857) );
  OAI21X1 U1813 ( .A(n301), .B(n1430), .C(n1857), .Y(n1078) );
  NAND2X1 U1814 ( .A(\mem<5><12> ), .B(n1394), .Y(n1858) );
  OAI21X1 U1815 ( .A(n301), .B(n1432), .C(n1858), .Y(n1079) );
  NAND2X1 U1816 ( .A(\mem<5><13> ), .B(n1394), .Y(n1859) );
  OAI21X1 U1817 ( .A(n301), .B(n36), .C(n1859), .Y(n1080) );
  NAND2X1 U1818 ( .A(\mem<5><14> ), .B(n1394), .Y(n1860) );
  OAI21X1 U1819 ( .A(n301), .B(n24), .C(n1860), .Y(n1081) );
  NAND2X1 U1820 ( .A(\mem<5><15> ), .B(n1394), .Y(n1861) );
  OAI21X1 U1821 ( .A(n301), .B(n14), .C(n1861), .Y(n1082) );
  NAND2X1 U1822 ( .A(\mem<4><0> ), .B(n1395), .Y(n1863) );
  OAI21X1 U1823 ( .A(n303), .B(n12), .C(n1863), .Y(n1083) );
  OAI21X1 U1824 ( .A(n303), .B(n1410), .C(n87), .Y(n1084) );
  OAI21X1 U1825 ( .A(n303), .B(n1412), .C(n89), .Y(n1085) );
  OAI21X1 U1826 ( .A(n303), .B(n1414), .C(n91), .Y(n1086) );
  OAI21X1 U1827 ( .A(n303), .B(n1416), .C(n93), .Y(n1087) );
  OAI21X1 U1828 ( .A(n303), .B(n1418), .C(n95), .Y(n1088) );
  OAI21X1 U1829 ( .A(n303), .B(n1420), .C(n97), .Y(n1089) );
  OAI21X1 U1830 ( .A(n303), .B(n1422), .C(n99), .Y(n1090) );
  NAND2X1 U1831 ( .A(\mem<4><8> ), .B(n1396), .Y(n1864) );
  OAI21X1 U1832 ( .A(n303), .B(n1424), .C(n1864), .Y(n1091) );
  NAND2X1 U1833 ( .A(\mem<4><9> ), .B(n1396), .Y(n1865) );
  OAI21X1 U1834 ( .A(n303), .B(n1426), .C(n1865), .Y(n1092) );
  NAND2X1 U1835 ( .A(\mem<4><10> ), .B(n1396), .Y(n1866) );
  OAI21X1 U1836 ( .A(n303), .B(n1428), .C(n1866), .Y(n1093) );
  NAND2X1 U1837 ( .A(\mem<4><11> ), .B(n1396), .Y(n1867) );
  OAI21X1 U1838 ( .A(n303), .B(n1430), .C(n1867), .Y(n1094) );
  NAND2X1 U1839 ( .A(\mem<4><12> ), .B(n1396), .Y(n1868) );
  OAI21X1 U1840 ( .A(n303), .B(n1432), .C(n1868), .Y(n1095) );
  NAND2X1 U1841 ( .A(\mem<4><13> ), .B(n1396), .Y(n1869) );
  OAI21X1 U1842 ( .A(n303), .B(n37), .C(n1869), .Y(n1096) );
  NAND2X1 U1843 ( .A(\mem<4><14> ), .B(n1396), .Y(n1870) );
  OAI21X1 U1844 ( .A(n303), .B(n27), .C(n1870), .Y(n1097) );
  NAND2X1 U1845 ( .A(\mem<4><15> ), .B(n1396), .Y(n1871) );
  OAI21X1 U1846 ( .A(n303), .B(n17), .C(n1871), .Y(n1098) );
  NAND2X1 U1847 ( .A(\mem<3><0> ), .B(n1397), .Y(n1873) );
  OAI21X1 U1848 ( .A(n305), .B(n11), .C(n1873), .Y(n1099) );
  OAI21X1 U1849 ( .A(n305), .B(n1410), .C(n101), .Y(n1100) );
  OAI21X1 U1850 ( .A(n305), .B(n1412), .C(n103), .Y(n1101) );
  OAI21X1 U1851 ( .A(n305), .B(n1414), .C(n105), .Y(n1102) );
  OAI21X1 U1852 ( .A(n305), .B(n1416), .C(n107), .Y(n1103) );
  OAI21X1 U1853 ( .A(n305), .B(n1418), .C(n109), .Y(n1104) );
  OAI21X1 U1854 ( .A(n305), .B(n1420), .C(n111), .Y(n1105) );
  OAI21X1 U1855 ( .A(n305), .B(n1422), .C(n113), .Y(n1106) );
  NAND2X1 U1856 ( .A(\mem<3><8> ), .B(n1398), .Y(n1874) );
  OAI21X1 U1857 ( .A(n305), .B(n1424), .C(n1874), .Y(n1107) );
  NAND2X1 U1858 ( .A(\mem<3><9> ), .B(n1398), .Y(n1875) );
  OAI21X1 U1859 ( .A(n305), .B(n1426), .C(n1875), .Y(n1108) );
  NAND2X1 U1860 ( .A(\mem<3><10> ), .B(n1398), .Y(n1876) );
  OAI21X1 U1861 ( .A(n305), .B(n1428), .C(n1876), .Y(n1109) );
  NAND2X1 U1862 ( .A(\mem<3><11> ), .B(n1398), .Y(n1877) );
  OAI21X1 U1863 ( .A(n305), .B(n1430), .C(n1877), .Y(n1110) );
  NAND2X1 U1864 ( .A(\mem<3><12> ), .B(n1398), .Y(n1878) );
  OAI21X1 U1865 ( .A(n305), .B(n1432), .C(n1878), .Y(n1111) );
  NAND2X1 U1866 ( .A(\mem<3><13> ), .B(n1398), .Y(n1879) );
  OAI21X1 U1867 ( .A(n305), .B(n37), .C(n1879), .Y(n1112) );
  NAND2X1 U1868 ( .A(\mem<3><14> ), .B(n1398), .Y(n1880) );
  OAI21X1 U1869 ( .A(n305), .B(n30), .C(n1880), .Y(n1113) );
  NAND2X1 U1870 ( .A(\mem<3><15> ), .B(n1398), .Y(n1881) );
  OAI21X1 U1871 ( .A(n305), .B(n17), .C(n1881), .Y(n1114) );
  NAND2X1 U1872 ( .A(\mem<2><0> ), .B(n1399), .Y(n1883) );
  OAI21X1 U1873 ( .A(n307), .B(n10), .C(n1883), .Y(n1115) );
  OAI21X1 U1874 ( .A(n307), .B(n1410), .C(n115), .Y(n1116) );
  OAI21X1 U1875 ( .A(n307), .B(n1412), .C(n117), .Y(n1117) );
  OAI21X1 U1876 ( .A(n307), .B(n1414), .C(n119), .Y(n1118) );
  OAI21X1 U1877 ( .A(n307), .B(n1416), .C(n121), .Y(n1119) );
  OAI21X1 U1878 ( .A(n307), .B(n1418), .C(n123), .Y(n1120) );
  OAI21X1 U1879 ( .A(n307), .B(n1420), .C(n125), .Y(n1121) );
  OAI21X1 U1880 ( .A(n307), .B(n1422), .C(n127), .Y(n1122) );
  NAND2X1 U1881 ( .A(\mem<2><8> ), .B(n1400), .Y(n1884) );
  OAI21X1 U1882 ( .A(n307), .B(n1424), .C(n1884), .Y(n1123) );
  NAND2X1 U1883 ( .A(\mem<2><9> ), .B(n1400), .Y(n1885) );
  OAI21X1 U1884 ( .A(n307), .B(n1426), .C(n1885), .Y(n1124) );
  NAND2X1 U1885 ( .A(\mem<2><10> ), .B(n1400), .Y(n1886) );
  OAI21X1 U1886 ( .A(n307), .B(n1428), .C(n1886), .Y(n1125) );
  NAND2X1 U1887 ( .A(\mem<2><11> ), .B(n1400), .Y(n1887) );
  OAI21X1 U1888 ( .A(n307), .B(n1430), .C(n1887), .Y(n1126) );
  NAND2X1 U1889 ( .A(\mem<2><12> ), .B(n1400), .Y(n1888) );
  OAI21X1 U1890 ( .A(n307), .B(n1432), .C(n1888), .Y(n1127) );
  NAND2X1 U1891 ( .A(\mem<2><13> ), .B(n1400), .Y(n1889) );
  OAI21X1 U1892 ( .A(n307), .B(n38), .C(n1889), .Y(n1128) );
  NAND2X1 U1893 ( .A(\mem<2><14> ), .B(n1400), .Y(n1890) );
  OAI21X1 U1894 ( .A(n307), .B(n30), .C(n1890), .Y(n1129) );
  NAND2X1 U1895 ( .A(\mem<2><15> ), .B(n1400), .Y(n1891) );
  OAI21X1 U1896 ( .A(n307), .B(n18), .C(n1891), .Y(n1130) );
  NAND2X1 U1897 ( .A(\mem<1><0> ), .B(n1401), .Y(n1893) );
  OAI21X1 U1898 ( .A(n309), .B(n9), .C(n1893), .Y(n1131) );
  OAI21X1 U1899 ( .A(n309), .B(n1410), .C(n129), .Y(n1132) );
  OAI21X1 U1900 ( .A(n309), .B(n1412), .C(n131), .Y(n1133) );
  OAI21X1 U1901 ( .A(n309), .B(n1414), .C(n133), .Y(n1134) );
  OAI21X1 U1902 ( .A(n309), .B(n1416), .C(n135), .Y(n1135) );
  OAI21X1 U1903 ( .A(n309), .B(n1418), .C(n137), .Y(n1136) );
  OAI21X1 U1904 ( .A(n309), .B(n1420), .C(n139), .Y(n1137) );
  OAI21X1 U1905 ( .A(n309), .B(n1422), .C(n141), .Y(n1138) );
  NAND2X1 U1906 ( .A(\mem<1><8> ), .B(n1402), .Y(n1894) );
  OAI21X1 U1907 ( .A(n309), .B(n1424), .C(n1894), .Y(n1139) );
  NAND2X1 U1908 ( .A(\mem<1><9> ), .B(n1402), .Y(n1895) );
  OAI21X1 U1909 ( .A(n309), .B(n1426), .C(n1895), .Y(n1140) );
  NAND2X1 U1910 ( .A(\mem<1><10> ), .B(n1402), .Y(n1896) );
  OAI21X1 U1911 ( .A(n309), .B(n1428), .C(n1896), .Y(n1141) );
  NAND2X1 U1912 ( .A(\mem<1><11> ), .B(n1402), .Y(n1897) );
  OAI21X1 U1913 ( .A(n309), .B(n1430), .C(n1897), .Y(n1142) );
  NAND2X1 U1914 ( .A(\mem<1><12> ), .B(n1402), .Y(n1898) );
  OAI21X1 U1915 ( .A(n309), .B(n1432), .C(n1898), .Y(n1143) );
  NAND2X1 U1916 ( .A(\mem<1><13> ), .B(n1402), .Y(n1899) );
  OAI21X1 U1917 ( .A(n309), .B(n40), .C(n1899), .Y(n1144) );
  NAND2X1 U1918 ( .A(\mem<1><14> ), .B(n1402), .Y(n1900) );
  OAI21X1 U1919 ( .A(n309), .B(n27), .C(n1900), .Y(n1145) );
  NAND2X1 U1920 ( .A(\mem<1><15> ), .B(n1402), .Y(n1901) );
  OAI21X1 U1921 ( .A(n309), .B(n20), .C(n1901), .Y(n1146) );
  NAND2X1 U1922 ( .A(\mem<0><0> ), .B(n1404), .Y(n1905) );
  OAI21X1 U1923 ( .A(n1403), .B(n8), .C(n1905), .Y(n1147) );
  NAND2X1 U1924 ( .A(\mem<0><1> ), .B(n1404), .Y(n1906) );
  OAI21X1 U1925 ( .A(n1403), .B(n1410), .C(n1906), .Y(n1148) );
  NAND2X1 U1926 ( .A(\mem<0><2> ), .B(n1404), .Y(n1907) );
  OAI21X1 U1927 ( .A(n1403), .B(n1412), .C(n1907), .Y(n1149) );
  NAND2X1 U1928 ( .A(\mem<0><3> ), .B(n1404), .Y(n1908) );
  OAI21X1 U1929 ( .A(n1403), .B(n1414), .C(n1908), .Y(n1150) );
  NAND2X1 U1930 ( .A(\mem<0><4> ), .B(n1404), .Y(n1909) );
  OAI21X1 U1931 ( .A(n1403), .B(n1416), .C(n1909), .Y(n1151) );
  NAND2X1 U1932 ( .A(\mem<0><5> ), .B(n1404), .Y(n1910) );
  OAI21X1 U1933 ( .A(n1403), .B(n1418), .C(n1910), .Y(n1152) );
  NAND2X1 U1934 ( .A(\mem<0><6> ), .B(n1404), .Y(n1911) );
  OAI21X1 U1935 ( .A(n1403), .B(n1420), .C(n1911), .Y(n1153) );
  NAND2X1 U1936 ( .A(\mem<0><7> ), .B(n1404), .Y(n1912) );
  OAI21X1 U1937 ( .A(n1403), .B(n1422), .C(n1912), .Y(n1154) );
  NAND2X1 U1938 ( .A(\mem<0><8> ), .B(n1405), .Y(n1913) );
  OAI21X1 U1939 ( .A(n1403), .B(n1424), .C(n1913), .Y(n1155) );
  NAND2X1 U1940 ( .A(\mem<0><9> ), .B(n1405), .Y(n1914) );
  OAI21X1 U1941 ( .A(n1403), .B(n1426), .C(n1914), .Y(n1156) );
  NAND2X1 U1942 ( .A(\mem<0><10> ), .B(n1405), .Y(n1915) );
  OAI21X1 U1943 ( .A(n1403), .B(n1428), .C(n1915), .Y(n1157) );
  NAND2X1 U1944 ( .A(\mem<0><11> ), .B(n1405), .Y(n1916) );
  OAI21X1 U1945 ( .A(n1403), .B(n1430), .C(n1916), .Y(n1158) );
  NAND2X1 U1946 ( .A(\mem<0><12> ), .B(n1405), .Y(n1917) );
  OAI21X1 U1947 ( .A(n1403), .B(n1432), .C(n1917), .Y(n1159) );
  NAND2X1 U1948 ( .A(\mem<0><13> ), .B(n1405), .Y(n1918) );
  OAI21X1 U1949 ( .A(n1403), .B(n39), .C(n1918), .Y(n1160) );
  NAND2X1 U1950 ( .A(\mem<0><14> ), .B(n1405), .Y(n1919) );
  OAI21X1 U1951 ( .A(n1403), .B(n29), .C(n1919), .Y(n1161) );
  NAND2X1 U1952 ( .A(\mem<0><15> ), .B(n1405), .Y(n1920) );
  OAI21X1 U1953 ( .A(n1403), .B(n19), .C(n1920), .Y(n1162) );
endmodule


module memc_Size16_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2160), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2161), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2162), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2163), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2164), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2165), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2166), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2167), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2168), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2169), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2170), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2171), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2172), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2173), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2174), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2175), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2176), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2177), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2178), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2179), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2180), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2181), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2182), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2183), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2184), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2185), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2186), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2187), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2188), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2189), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2190), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2191), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2192), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2193), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2194), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2195), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2196), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2197), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2198), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2199), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2200), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2201), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2202), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2203), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2204), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2205), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2206), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2207), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2208), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2209), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2210), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2211), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2212), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2213), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2214), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2215), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2216), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2217), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2218), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2219), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2220), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2221), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2222), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2223), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2224), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2225), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2226), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2227), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2228), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2229), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2230), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2231), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2232), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2233), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2234), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2235), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2236), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2237), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2238), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2239), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2240), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2241), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2242), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2243), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2244), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2245), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2246), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2247), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2248), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2249), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2250), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2251), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2252), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2253), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2254), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2255), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2256), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2257), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2258), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2259), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2260), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2261), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2262), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2263), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2264), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2265), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2266), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2267), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2268), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2269), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2270), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2271), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2272), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2273), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2274), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2275), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2276), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2277), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2278), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2279), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2280), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2281), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2282), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2283), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2284), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2285), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2286), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2287), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2288), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2289), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2290), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2291), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2292), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2293), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2294), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2295), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2296), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2297), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2298), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2299), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2300), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2301), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2302), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2303), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2304), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2305), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2306), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2307), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2308), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2309), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2310), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2311), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2312), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2313), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2314), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2315), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2316), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2317), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2318), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2319), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2320), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2321), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2322), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2323), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2324), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2325), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2326), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2327), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2328), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2329), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2330), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2331), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2332), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2333), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2334), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2335), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2336), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2337), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2338), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2339), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2340), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2341), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2342), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2343), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2344), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2345), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2346), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2347), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2348), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2349), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2350), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2351), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2352), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2353), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2354), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2355), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2356), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2357), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2358), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2359), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2360), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2361), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2362), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2363), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2364), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2365), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2366), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2367), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2368), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2369), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2370), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2371), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2372), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2373), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2374), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2375), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2376), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2377), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2378), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2379), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2380), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2381), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2382), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2383), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2384), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2385), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2386), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2387), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2388), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2389), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2390), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2391), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2392), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2393), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2394), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2395), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2396), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2397), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2398), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2399), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2400), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2401), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2402), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2403), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2404), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2405), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2406), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2407), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2408), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2409), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2410), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2411), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2412), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2413), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2414), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2415), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2416), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2417), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2418), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2419), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2420), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2421), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2422), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2423), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2424), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2425), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2426), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2427), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2428), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2429), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2430), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2431), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2432), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2433), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2434), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2435), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2436), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2437), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2438), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2439), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2440), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2441), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2442), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2443), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2444), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2445), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2446), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2447), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2448), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2449), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2450), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2451), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2452), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2453), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2454), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2455), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2456), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2457), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2458), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2459), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2460), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2461), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2462), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2463), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2464), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2465), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2466), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2467), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2468), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2469), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2470), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2471), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2472), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2473), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2474), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2475), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2476), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2477), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2478), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2479), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2480), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2481), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2482), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2483), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2484), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2485), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2486), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2487), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2488), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2489), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2490), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2491), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2492), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2493), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2494), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2495), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2496), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2497), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2498), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2499), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2500), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2501), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2502), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2503), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2504), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2505), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2506), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2507), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2508), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2509), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2510), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2511), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2512), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2513), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2514), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2515), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2516), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2517), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2518), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2519), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2520), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2521), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2522), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2523), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2524), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2525), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2526), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2527), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2528), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2529), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2530), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2531), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2532), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2533), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2534), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2535), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2536), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2537), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2538), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2539), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2540), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2541), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2542), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2543), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2544), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2545), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2546), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2547), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2548), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2549), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2550), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2551), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2552), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2553), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2554), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2555), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2556), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2557), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2558), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2559), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2560), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2561), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2562), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2563), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2564), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2565), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2566), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2567), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2568), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2569), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2570), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2571), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2572), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2573), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2574), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2575), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2576), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2577), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2578), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2579), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2580), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2581), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2582), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2583), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2584), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2585), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2586), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2587), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2588), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2589), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2590), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2591), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2592), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2593), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2594), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2595), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2596), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2597), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2598), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2599), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2600), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2601), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2602), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2603), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2604), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2605), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2606), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2607), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2608), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2609), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2610), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2611), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2612), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2613), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2614), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2615), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2616), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2617), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2618), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2619), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2620), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2621), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2622), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2623), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2624), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2625), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2626), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2627), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2628), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2629), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2630), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2631), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2632), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2633), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2634), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2635), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2636), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2637), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2638), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2639), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2640), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2641), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2642), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2643), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2644), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2645), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2646), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2647), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2648), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2649), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2650), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2651), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2652), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2653), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2654), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2655), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2656), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2657), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2658), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2659), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2660), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2661), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2662), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2663), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2664), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2665), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2666), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2667), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2668), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2669), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2670), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2671), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2672) );
  INVX2 U2 ( .A(n1946), .Y(n1862) );
  INVX4 U3 ( .A(n1862), .Y(n1843) );
  INVX2 U4 ( .A(n1843), .Y(n1848) );
  INVX1 U5 ( .A(n1843), .Y(n1856) );
  INVX2 U6 ( .A(n1843), .Y(n1853) );
  INVX1 U7 ( .A(n1843), .Y(n1852) );
  INVX2 U8 ( .A(n1843), .Y(n1855) );
  INVX1 U9 ( .A(n1843), .Y(n1851) );
  INVX1 U10 ( .A(n1862), .Y(n1842) );
  INVX1 U11 ( .A(n1841), .Y(n1861) );
  INVX2 U12 ( .A(n1843), .Y(n1850) );
  INVX2 U13 ( .A(n1843), .Y(n1849) );
  INVX1 U14 ( .A(n1841), .Y(n1860) );
  INVX2 U15 ( .A(n1843), .Y(n1846) );
  INVX1 U16 ( .A(n1810), .Y(N25) );
  INVX1 U17 ( .A(n1945), .Y(n1841) );
  INVX1 U18 ( .A(n1829), .Y(n1830) );
  INVX1 U19 ( .A(n1829), .Y(n1831) );
  INVX1 U20 ( .A(n1829), .Y(n1832) );
  INVX2 U21 ( .A(n1829), .Y(n1839) );
  INVX1 U22 ( .A(n1951), .Y(n1822) );
  INVX1 U23 ( .A(n1951), .Y(n1821) );
  INVX1 U24 ( .A(n1951), .Y(n1820) );
  INVX1 U25 ( .A(n1803), .Y(N32) );
  INVX1 U26 ( .A(n1804), .Y(N31) );
  INVX1 U27 ( .A(n1805), .Y(N30) );
  INVX1 U28 ( .A(n1806), .Y(N29) );
  INVX1 U29 ( .A(n1807), .Y(N28) );
  INVX1 U30 ( .A(n1808), .Y(N27) );
  INVX1 U31 ( .A(n1809), .Y(N26) );
  INVX1 U32 ( .A(n1811), .Y(N24) );
  INVX1 U33 ( .A(n1812), .Y(N23) );
  INVX1 U34 ( .A(n1813), .Y(N22) );
  INVX1 U35 ( .A(n1814), .Y(N21) );
  INVX1 U36 ( .A(n1815), .Y(N20) );
  INVX1 U37 ( .A(n1816), .Y(N19) );
  INVX1 U38 ( .A(n1817), .Y(N18) );
  INVX1 U39 ( .A(n1818), .Y(N17) );
  INVX1 U40 ( .A(n1947), .Y(n1828) );
  INVX1 U41 ( .A(n1949), .Y(n1827) );
  INVX1 U42 ( .A(n1949), .Y(n1825) );
  INVX1 U43 ( .A(n1949), .Y(n1826) );
  INVX1 U44 ( .A(N14), .Y(n1952) );
  INVX1 U45 ( .A(n1949), .Y(n1824) );
  INVX1 U46 ( .A(n1949), .Y(n1823) );
  INVX1 U47 ( .A(n1952), .Y(n1819) );
  INVX1 U48 ( .A(rst), .Y(n1944) );
  INVX1 U49 ( .A(n1947), .Y(n1829) );
  INVX1 U50 ( .A(n1239), .Y(n1863) );
  INVX1 U51 ( .A(n1240), .Y(n1870) );
  INVX1 U52 ( .A(n1241), .Y(n1887) );
  INVX1 U53 ( .A(n1242), .Y(n1904) );
  INVX2 U54 ( .A(n2), .Y(n1) );
  INVX2 U55 ( .A(n2), .Y(n3) );
  OR2X2 U56 ( .A(write), .B(rst), .Y(n2) );
  AND2X2 U57 ( .A(write), .B(n1944), .Y(n4) );
  AND2X2 U58 ( .A(\data_in<0> ), .B(n1909), .Y(n5) );
  AND2X2 U59 ( .A(n1907), .B(n1243), .Y(n6) );
  AND2X2 U60 ( .A(\data_in<1> ), .B(n1909), .Y(n7) );
  AND2X2 U61 ( .A(\data_in<2> ), .B(n1909), .Y(n8) );
  AND2X2 U62 ( .A(\data_in<3> ), .B(n1909), .Y(n9) );
  AND2X2 U63 ( .A(\data_in<4> ), .B(n1909), .Y(n10) );
  AND2X2 U64 ( .A(\data_in<5> ), .B(n1909), .Y(n11) );
  AND2X2 U65 ( .A(\data_in<6> ), .B(n1909), .Y(n12) );
  AND2X2 U66 ( .A(\data_in<7> ), .B(n1909), .Y(n13) );
  AND2X2 U67 ( .A(\data_in<8> ), .B(n1909), .Y(n14) );
  AND2X2 U68 ( .A(\data_in<9> ), .B(n1909), .Y(n15) );
  AND2X2 U69 ( .A(\data_in<10> ), .B(n1909), .Y(n16) );
  AND2X2 U70 ( .A(\data_in<11> ), .B(n1908), .Y(n17) );
  AND2X2 U71 ( .A(\data_in<12> ), .B(n1908), .Y(n18) );
  AND2X2 U72 ( .A(\data_in<13> ), .B(n1908), .Y(n19) );
  AND2X2 U73 ( .A(\data_in<14> ), .B(n1908), .Y(n20) );
  AND2X2 U74 ( .A(\data_in<15> ), .B(n1908), .Y(n21) );
  AND2X2 U75 ( .A(n1907), .B(n1247), .Y(n22) );
  AND2X2 U76 ( .A(n1907), .B(n1251), .Y(n23) );
  AND2X2 U77 ( .A(n1907), .B(n1255), .Y(n24) );
  AND2X2 U78 ( .A(n1907), .B(n1259), .Y(n25) );
  AND2X2 U79 ( .A(n1907), .B(n1263), .Y(n26) );
  AND2X2 U80 ( .A(n1907), .B(n1267), .Y(n27) );
  AND2X2 U81 ( .A(n1907), .B(n1239), .Y(n28) );
  AND2X2 U82 ( .A(n1907), .B(n1273), .Y(n29) );
  AND2X2 U83 ( .A(n1907), .B(n1277), .Y(n30) );
  AND2X2 U84 ( .A(n1907), .B(n1281), .Y(n31) );
  AND2X2 U85 ( .A(n1907), .B(n1285), .Y(n32) );
  AND2X2 U86 ( .A(n1908), .B(n1289), .Y(n33) );
  INVX1 U87 ( .A(n33), .Y(n34) );
  AND2X2 U88 ( .A(n1909), .B(n1291), .Y(n35) );
  INVX1 U89 ( .A(n35), .Y(n36) );
  AND2X2 U90 ( .A(n1908), .B(n1293), .Y(n37) );
  INVX1 U91 ( .A(n37), .Y(n38) );
  AND2X2 U92 ( .A(n1909), .B(n1240), .Y(n39) );
  INVX1 U93 ( .A(n39), .Y(n40) );
  AND2X2 U94 ( .A(n1909), .B(n1295), .Y(n41) );
  INVX1 U95 ( .A(n41), .Y(n42) );
  AND2X2 U96 ( .A(n1909), .B(n1297), .Y(n43) );
  INVX1 U97 ( .A(n43), .Y(n44) );
  AND2X2 U98 ( .A(n1908), .B(n1299), .Y(n45) );
  INVX1 U99 ( .A(n45), .Y(n46) );
  AND2X2 U100 ( .A(n1909), .B(n1301), .Y(n47) );
  INVX1 U101 ( .A(n47), .Y(n48) );
  AND2X2 U102 ( .A(n1908), .B(n1303), .Y(n49) );
  INVX1 U103 ( .A(n49), .Y(n50) );
  AND2X2 U104 ( .A(n1909), .B(n1305), .Y(n51) );
  INVX1 U105 ( .A(n51), .Y(n52) );
  AND2X2 U106 ( .A(n1908), .B(n1307), .Y(n53) );
  INVX1 U107 ( .A(n53), .Y(n54) );
  AND2X2 U108 ( .A(n1908), .B(n1241), .Y(n55) );
  INVX1 U109 ( .A(n55), .Y(n56) );
  AND2X2 U110 ( .A(n1908), .B(n1309), .Y(n57) );
  INVX1 U111 ( .A(n57), .Y(n58) );
  AND2X2 U112 ( .A(n1908), .B(n1311), .Y(n59) );
  INVX1 U113 ( .A(n59), .Y(n60) );
  AND2X2 U114 ( .A(n1908), .B(n1313), .Y(n61) );
  INVX1 U115 ( .A(n61), .Y(n62) );
  AND2X2 U116 ( .A(n1908), .B(n1315), .Y(n63) );
  INVX1 U117 ( .A(n63), .Y(n64) );
  AND2X2 U118 ( .A(n1908), .B(n1317), .Y(n65) );
  INVX1 U119 ( .A(n65), .Y(n66) );
  AND2X2 U120 ( .A(n1908), .B(n1319), .Y(n67) );
  INVX1 U121 ( .A(n67), .Y(n68) );
  AND2X2 U122 ( .A(n1908), .B(n1321), .Y(n69) );
  INVX1 U123 ( .A(n69), .Y(n70) );
  AND2X2 U124 ( .A(n1909), .B(n1242), .Y(n71) );
  INVX1 U125 ( .A(n71), .Y(n72) );
  AND2X2 U126 ( .A(\mem<19><0> ), .B(n1864), .Y(n73) );
  INVX1 U127 ( .A(n73), .Y(n74) );
  AND2X2 U128 ( .A(\mem<19><1> ), .B(n1864), .Y(n75) );
  INVX1 U129 ( .A(n75), .Y(n76) );
  AND2X2 U130 ( .A(\mem<19><2> ), .B(n1864), .Y(n77) );
  INVX1 U131 ( .A(n77), .Y(n78) );
  AND2X2 U132 ( .A(\mem<19><3> ), .B(n1864), .Y(n79) );
  INVX1 U133 ( .A(n79), .Y(n80) );
  AND2X2 U134 ( .A(\mem<19><4> ), .B(n1864), .Y(n81) );
  INVX1 U135 ( .A(n81), .Y(n82) );
  AND2X2 U136 ( .A(\mem<19><5> ), .B(n1864), .Y(n83) );
  INVX1 U137 ( .A(n83), .Y(n84) );
  AND2X2 U138 ( .A(\mem<19><6> ), .B(n1864), .Y(n85) );
  INVX1 U139 ( .A(n85), .Y(n86) );
  AND2X2 U140 ( .A(\mem<19><7> ), .B(n1864), .Y(n87) );
  INVX1 U141 ( .A(n87), .Y(n88) );
  AND2X2 U142 ( .A(\mem<19><8> ), .B(n1865), .Y(n89) );
  INVX1 U143 ( .A(n89), .Y(n90) );
  AND2X2 U144 ( .A(\mem<19><9> ), .B(n1865), .Y(n91) );
  INVX1 U145 ( .A(n91), .Y(n92) );
  AND2X2 U146 ( .A(\mem<19><10> ), .B(n1865), .Y(n93) );
  INVX1 U147 ( .A(n93), .Y(n94) );
  AND2X2 U148 ( .A(\mem<19><11> ), .B(n1865), .Y(n95) );
  INVX1 U149 ( .A(n95), .Y(n96) );
  AND2X2 U150 ( .A(\mem<19><12> ), .B(n1865), .Y(n97) );
  INVX1 U151 ( .A(n97), .Y(n98) );
  AND2X2 U152 ( .A(\mem<19><13> ), .B(n1865), .Y(n99) );
  INVX1 U153 ( .A(n99), .Y(n100) );
  AND2X2 U154 ( .A(\mem<19><14> ), .B(n1865), .Y(n101) );
  INVX1 U155 ( .A(n101), .Y(n102) );
  AND2X2 U156 ( .A(\mem<19><15> ), .B(n1865), .Y(n103) );
  INVX1 U157 ( .A(n103), .Y(n104) );
  AND2X2 U158 ( .A(\mem<18><0> ), .B(n1866), .Y(n105) );
  INVX1 U159 ( .A(n105), .Y(n106) );
  AND2X2 U160 ( .A(\mem<18><1> ), .B(n1866), .Y(n107) );
  INVX1 U161 ( .A(n107), .Y(n108) );
  AND2X2 U162 ( .A(\mem<18><2> ), .B(n1866), .Y(n109) );
  INVX1 U163 ( .A(n109), .Y(n110) );
  AND2X2 U164 ( .A(\mem<18><3> ), .B(n1866), .Y(n111) );
  INVX1 U165 ( .A(n111), .Y(n112) );
  AND2X2 U166 ( .A(\mem<18><4> ), .B(n1866), .Y(n113) );
  INVX1 U167 ( .A(n113), .Y(n114) );
  AND2X2 U168 ( .A(\mem<18><5> ), .B(n1866), .Y(n115) );
  INVX1 U169 ( .A(n115), .Y(n116) );
  AND2X2 U170 ( .A(\mem<18><6> ), .B(n1866), .Y(n117) );
  INVX1 U171 ( .A(n117), .Y(n118) );
  AND2X2 U172 ( .A(\mem<18><7> ), .B(n1866), .Y(n119) );
  INVX1 U173 ( .A(n119), .Y(n120) );
  AND2X2 U174 ( .A(\mem<18><8> ), .B(n1867), .Y(n121) );
  INVX1 U175 ( .A(n121), .Y(n122) );
  AND2X2 U176 ( .A(\mem<18><9> ), .B(n1867), .Y(n123) );
  INVX1 U177 ( .A(n123), .Y(n124) );
  AND2X2 U178 ( .A(\mem<18><10> ), .B(n1867), .Y(n125) );
  INVX1 U179 ( .A(n125), .Y(n126) );
  AND2X2 U180 ( .A(\mem<18><11> ), .B(n1867), .Y(n127) );
  INVX1 U181 ( .A(n127), .Y(n128) );
  AND2X2 U182 ( .A(\mem<18><12> ), .B(n1867), .Y(n129) );
  INVX1 U183 ( .A(n129), .Y(n130) );
  AND2X2 U184 ( .A(\mem<18><13> ), .B(n1867), .Y(n131) );
  INVX1 U185 ( .A(n131), .Y(n132) );
  AND2X2 U186 ( .A(\mem<18><14> ), .B(n1867), .Y(n133) );
  INVX1 U187 ( .A(n133), .Y(n134) );
  AND2X2 U188 ( .A(\mem<18><15> ), .B(n1867), .Y(n135) );
  INVX1 U189 ( .A(n135), .Y(n136) );
  AND2X2 U190 ( .A(\mem<17><0> ), .B(n1868), .Y(n137) );
  INVX1 U191 ( .A(n137), .Y(n138) );
  AND2X2 U192 ( .A(\mem<17><1> ), .B(n1868), .Y(n139) );
  INVX1 U193 ( .A(n139), .Y(n140) );
  AND2X2 U194 ( .A(\mem<17><2> ), .B(n1868), .Y(n141) );
  INVX1 U195 ( .A(n141), .Y(n142) );
  AND2X2 U196 ( .A(\mem<17><3> ), .B(n1868), .Y(n143) );
  INVX1 U197 ( .A(n143), .Y(n144) );
  AND2X2 U198 ( .A(\mem<17><4> ), .B(n1868), .Y(n145) );
  INVX1 U199 ( .A(n145), .Y(n146) );
  AND2X2 U200 ( .A(\mem<17><5> ), .B(n1868), .Y(n147) );
  INVX1 U201 ( .A(n147), .Y(n148) );
  AND2X2 U202 ( .A(\mem<17><6> ), .B(n1868), .Y(n149) );
  INVX1 U203 ( .A(n149), .Y(n150) );
  AND2X2 U204 ( .A(\mem<17><7> ), .B(n1868), .Y(n151) );
  INVX1 U205 ( .A(n151), .Y(n152) );
  AND2X2 U206 ( .A(\mem<17><8> ), .B(n1869), .Y(n153) );
  INVX1 U207 ( .A(n153), .Y(n154) );
  AND2X2 U208 ( .A(\mem<17><9> ), .B(n1869), .Y(n155) );
  INVX1 U209 ( .A(n155), .Y(n156) );
  AND2X2 U210 ( .A(\mem<17><10> ), .B(n1869), .Y(n157) );
  INVX1 U211 ( .A(n157), .Y(n158) );
  AND2X2 U212 ( .A(\mem<17><11> ), .B(n1869), .Y(n159) );
  INVX1 U213 ( .A(n159), .Y(n160) );
  AND2X2 U214 ( .A(\mem<17><12> ), .B(n1869), .Y(n161) );
  INVX1 U215 ( .A(n161), .Y(n162) );
  AND2X2 U216 ( .A(\mem<17><13> ), .B(n1869), .Y(n163) );
  INVX1 U217 ( .A(n163), .Y(n164) );
  AND2X2 U218 ( .A(\mem<17><14> ), .B(n1869), .Y(n165) );
  INVX1 U219 ( .A(n165), .Y(n166) );
  AND2X2 U220 ( .A(\mem<17><15> ), .B(n1869), .Y(n167) );
  INVX1 U221 ( .A(n167), .Y(n168) );
  AND2X2 U222 ( .A(\mem<16><0> ), .B(n1871), .Y(n169) );
  INVX1 U223 ( .A(n169), .Y(n170) );
  AND2X2 U224 ( .A(\mem<16><1> ), .B(n1871), .Y(n171) );
  INVX1 U225 ( .A(n171), .Y(n172) );
  AND2X2 U226 ( .A(\mem<16><2> ), .B(n1871), .Y(n173) );
  INVX1 U227 ( .A(n173), .Y(n174) );
  AND2X2 U228 ( .A(\mem<16><3> ), .B(n1871), .Y(n175) );
  INVX1 U229 ( .A(n175), .Y(n176) );
  AND2X2 U230 ( .A(\mem<16><4> ), .B(n1871), .Y(n177) );
  INVX1 U231 ( .A(n177), .Y(n178) );
  AND2X2 U232 ( .A(\mem<16><5> ), .B(n1871), .Y(n179) );
  INVX1 U233 ( .A(n179), .Y(n180) );
  AND2X2 U234 ( .A(\mem<16><6> ), .B(n1871), .Y(n181) );
  INVX1 U235 ( .A(n181), .Y(n182) );
  AND2X2 U236 ( .A(\mem<16><7> ), .B(n1871), .Y(n183) );
  INVX1 U237 ( .A(n183), .Y(n184) );
  AND2X2 U238 ( .A(\mem<16><8> ), .B(n1872), .Y(n185) );
  INVX1 U239 ( .A(n185), .Y(n186) );
  AND2X2 U240 ( .A(\mem<16><9> ), .B(n1872), .Y(n187) );
  INVX1 U241 ( .A(n187), .Y(n188) );
  AND2X2 U242 ( .A(\mem<16><10> ), .B(n1872), .Y(n189) );
  INVX1 U243 ( .A(n189), .Y(n190) );
  AND2X2 U244 ( .A(\mem<16><11> ), .B(n1872), .Y(n191) );
  INVX1 U245 ( .A(n191), .Y(n192) );
  AND2X2 U246 ( .A(\mem<16><12> ), .B(n1872), .Y(n193) );
  INVX1 U247 ( .A(n193), .Y(n194) );
  AND2X2 U248 ( .A(\mem<16><13> ), .B(n1872), .Y(n195) );
  INVX1 U249 ( .A(n195), .Y(n196) );
  AND2X2 U250 ( .A(\mem<16><14> ), .B(n1872), .Y(n197) );
  INVX1 U251 ( .A(n197), .Y(n198) );
  AND2X2 U252 ( .A(\mem<16><15> ), .B(n1872), .Y(n199) );
  INVX1 U253 ( .A(n199), .Y(n200) );
  AND2X2 U254 ( .A(\mem<15><0> ), .B(n1873), .Y(n201) );
  INVX1 U255 ( .A(n201), .Y(n202) );
  AND2X2 U256 ( .A(\mem<15><1> ), .B(n1873), .Y(n203) );
  INVX1 U257 ( .A(n203), .Y(n204) );
  AND2X2 U258 ( .A(\mem<15><2> ), .B(n1873), .Y(n205) );
  INVX1 U259 ( .A(n205), .Y(n206) );
  AND2X2 U260 ( .A(\mem<15><3> ), .B(n1873), .Y(n207) );
  INVX1 U261 ( .A(n207), .Y(n208) );
  AND2X2 U262 ( .A(\mem<15><4> ), .B(n1873), .Y(n209) );
  INVX1 U263 ( .A(n209), .Y(n210) );
  AND2X2 U264 ( .A(\mem<15><5> ), .B(n1873), .Y(n211) );
  INVX1 U265 ( .A(n211), .Y(n212) );
  AND2X2 U266 ( .A(\mem<15><6> ), .B(n1873), .Y(n213) );
  INVX1 U267 ( .A(n213), .Y(n215) );
  AND2X2 U268 ( .A(\mem<15><7> ), .B(n1873), .Y(n216) );
  INVX1 U269 ( .A(n216), .Y(n217) );
  AND2X2 U270 ( .A(\mem<15><8> ), .B(n1874), .Y(n218) );
  INVX1 U271 ( .A(n218), .Y(n219) );
  AND2X2 U272 ( .A(\mem<15><9> ), .B(n1874), .Y(n220) );
  INVX1 U273 ( .A(n220), .Y(n221) );
  AND2X2 U274 ( .A(\mem<15><10> ), .B(n1874), .Y(n222) );
  INVX1 U275 ( .A(n222), .Y(n223) );
  AND2X2 U276 ( .A(\mem<15><11> ), .B(n1874), .Y(n224) );
  INVX1 U277 ( .A(n224), .Y(n225) );
  AND2X2 U278 ( .A(\mem<15><12> ), .B(n1874), .Y(n226) );
  INVX1 U279 ( .A(n226), .Y(n227) );
  AND2X2 U280 ( .A(\mem<15><13> ), .B(n1874), .Y(n228) );
  INVX1 U281 ( .A(n228), .Y(n229) );
  AND2X2 U282 ( .A(\mem<15><14> ), .B(n1874), .Y(n230) );
  INVX1 U283 ( .A(n230), .Y(n231) );
  AND2X2 U284 ( .A(\mem<15><15> ), .B(n1874), .Y(n232) );
  INVX1 U285 ( .A(n232), .Y(n233) );
  AND2X2 U286 ( .A(\mem<14><0> ), .B(n1875), .Y(n234) );
  INVX1 U287 ( .A(n234), .Y(n235) );
  AND2X2 U288 ( .A(\mem<14><1> ), .B(n1875), .Y(n236) );
  INVX1 U289 ( .A(n236), .Y(n237) );
  AND2X2 U290 ( .A(\mem<14><2> ), .B(n1875), .Y(n238) );
  INVX1 U291 ( .A(n238), .Y(n239) );
  AND2X2 U292 ( .A(\mem<14><3> ), .B(n1875), .Y(n240) );
  INVX1 U293 ( .A(n240), .Y(n241) );
  AND2X2 U294 ( .A(\mem<14><4> ), .B(n1875), .Y(n242) );
  INVX1 U295 ( .A(n242), .Y(n243) );
  AND2X2 U296 ( .A(\mem<14><5> ), .B(n1875), .Y(n244) );
  INVX1 U297 ( .A(n244), .Y(n245) );
  AND2X2 U298 ( .A(\mem<14><6> ), .B(n1875), .Y(n246) );
  INVX1 U299 ( .A(n246), .Y(n247) );
  AND2X2 U300 ( .A(\mem<14><7> ), .B(n1875), .Y(n248) );
  INVX1 U301 ( .A(n248), .Y(n249) );
  AND2X2 U302 ( .A(\mem<14><8> ), .B(n1876), .Y(n250) );
  INVX1 U303 ( .A(n250), .Y(n251) );
  AND2X2 U304 ( .A(\mem<14><9> ), .B(n1876), .Y(n252) );
  INVX1 U305 ( .A(n252), .Y(n253) );
  AND2X2 U306 ( .A(\mem<14><10> ), .B(n1876), .Y(n254) );
  INVX1 U307 ( .A(n254), .Y(n255) );
  AND2X2 U308 ( .A(\mem<14><11> ), .B(n1876), .Y(n256) );
  INVX1 U309 ( .A(n256), .Y(n257) );
  AND2X2 U310 ( .A(\mem<14><12> ), .B(n1876), .Y(n258) );
  INVX1 U311 ( .A(n258), .Y(n259) );
  AND2X2 U312 ( .A(\mem<14><13> ), .B(n1876), .Y(n260) );
  INVX1 U313 ( .A(n260), .Y(n261) );
  AND2X2 U314 ( .A(\mem<14><14> ), .B(n1876), .Y(n262) );
  INVX1 U315 ( .A(n262), .Y(n263) );
  AND2X2 U316 ( .A(\mem<14><15> ), .B(n1876), .Y(n264) );
  INVX1 U317 ( .A(n264), .Y(n265) );
  AND2X2 U318 ( .A(\mem<13><0> ), .B(n1877), .Y(n266) );
  INVX1 U319 ( .A(n266), .Y(n267) );
  AND2X2 U320 ( .A(\mem<13><1> ), .B(n1877), .Y(n268) );
  INVX1 U321 ( .A(n268), .Y(n269) );
  AND2X2 U322 ( .A(\mem<13><2> ), .B(n1877), .Y(n270) );
  INVX1 U323 ( .A(n270), .Y(n271) );
  AND2X2 U324 ( .A(\mem<13><3> ), .B(n1877), .Y(n272) );
  INVX1 U325 ( .A(n272), .Y(n273) );
  AND2X2 U326 ( .A(\mem<13><4> ), .B(n1877), .Y(n274) );
  INVX1 U327 ( .A(n274), .Y(n275) );
  AND2X2 U328 ( .A(\mem<13><5> ), .B(n1877), .Y(n276) );
  INVX1 U329 ( .A(n276), .Y(n277) );
  AND2X2 U330 ( .A(\mem<13><6> ), .B(n1877), .Y(n278) );
  INVX1 U331 ( .A(n278), .Y(n279) );
  AND2X2 U332 ( .A(\mem<13><7> ), .B(n1877), .Y(n280) );
  INVX1 U333 ( .A(n280), .Y(n281) );
  AND2X2 U334 ( .A(\mem<13><8> ), .B(n1878), .Y(n282) );
  INVX1 U335 ( .A(n282), .Y(n283) );
  AND2X2 U336 ( .A(\mem<13><9> ), .B(n1878), .Y(n284) );
  INVX1 U337 ( .A(n284), .Y(n285) );
  AND2X2 U338 ( .A(\mem<13><10> ), .B(n1878), .Y(n286) );
  INVX1 U339 ( .A(n286), .Y(n287) );
  AND2X2 U340 ( .A(\mem<13><11> ), .B(n1878), .Y(n288) );
  INVX1 U341 ( .A(n288), .Y(n289) );
  AND2X2 U342 ( .A(\mem<13><12> ), .B(n1878), .Y(n290) );
  INVX1 U343 ( .A(n290), .Y(n291) );
  AND2X2 U344 ( .A(\mem<13><13> ), .B(n1878), .Y(n292) );
  INVX1 U345 ( .A(n292), .Y(n293) );
  AND2X2 U346 ( .A(\mem<13><14> ), .B(n1878), .Y(n294) );
  INVX1 U347 ( .A(n294), .Y(n295) );
  AND2X2 U348 ( .A(\mem<13><15> ), .B(n1878), .Y(n296) );
  INVX1 U349 ( .A(n296), .Y(n297) );
  AND2X2 U350 ( .A(\mem<12><0> ), .B(n1879), .Y(n298) );
  INVX1 U351 ( .A(n298), .Y(n299) );
  AND2X2 U352 ( .A(\mem<12><1> ), .B(n1879), .Y(n300) );
  INVX1 U353 ( .A(n300), .Y(n301) );
  AND2X2 U354 ( .A(\mem<12><2> ), .B(n1879), .Y(n302) );
  INVX1 U355 ( .A(n302), .Y(n303) );
  AND2X2 U356 ( .A(\mem<12><3> ), .B(n1879), .Y(n304) );
  INVX1 U357 ( .A(n304), .Y(n305) );
  AND2X2 U358 ( .A(\mem<12><4> ), .B(n1879), .Y(n306) );
  INVX1 U359 ( .A(n306), .Y(n307) );
  AND2X2 U360 ( .A(\mem<12><5> ), .B(n1879), .Y(n308) );
  INVX1 U361 ( .A(n308), .Y(n309) );
  AND2X2 U362 ( .A(\mem<12><6> ), .B(n1879), .Y(n310) );
  INVX1 U363 ( .A(n310), .Y(n311) );
  AND2X2 U364 ( .A(\mem<12><7> ), .B(n1879), .Y(n312) );
  INVX1 U365 ( .A(n312), .Y(n313) );
  AND2X2 U366 ( .A(\mem<12><8> ), .B(n1880), .Y(n314) );
  INVX1 U367 ( .A(n314), .Y(n315) );
  AND2X2 U368 ( .A(\mem<12><9> ), .B(n1880), .Y(n316) );
  INVX1 U369 ( .A(n316), .Y(n317) );
  AND2X2 U370 ( .A(\mem<12><10> ), .B(n1880), .Y(n318) );
  INVX1 U371 ( .A(n318), .Y(n319) );
  AND2X2 U372 ( .A(\mem<12><11> ), .B(n1880), .Y(n320) );
  INVX1 U373 ( .A(n320), .Y(n321) );
  AND2X2 U374 ( .A(\mem<12><12> ), .B(n1880), .Y(n322) );
  INVX1 U375 ( .A(n322), .Y(n323) );
  AND2X2 U376 ( .A(\mem<12><13> ), .B(n1880), .Y(n324) );
  INVX1 U377 ( .A(n324), .Y(n325) );
  AND2X2 U378 ( .A(\mem<12><14> ), .B(n1880), .Y(n326) );
  INVX1 U379 ( .A(n326), .Y(n327) );
  AND2X2 U380 ( .A(\mem<12><15> ), .B(n1880), .Y(n328) );
  INVX1 U381 ( .A(n328), .Y(n329) );
  AND2X2 U382 ( .A(\mem<11><0> ), .B(n1881), .Y(n330) );
  INVX1 U383 ( .A(n330), .Y(n331) );
  AND2X2 U384 ( .A(\mem<11><1> ), .B(n1881), .Y(n332) );
  INVX1 U385 ( .A(n332), .Y(n333) );
  AND2X2 U386 ( .A(\mem<11><2> ), .B(n1881), .Y(n334) );
  INVX1 U387 ( .A(n334), .Y(n335) );
  AND2X2 U388 ( .A(\mem<11><3> ), .B(n1881), .Y(n336) );
  INVX1 U389 ( .A(n336), .Y(n337) );
  AND2X2 U390 ( .A(\mem<11><4> ), .B(n1881), .Y(n338) );
  INVX1 U391 ( .A(n338), .Y(n339) );
  AND2X2 U392 ( .A(\mem<11><5> ), .B(n1881), .Y(n340) );
  INVX1 U393 ( .A(n340), .Y(n341) );
  AND2X2 U394 ( .A(\mem<11><6> ), .B(n1881), .Y(n342) );
  INVX1 U395 ( .A(n342), .Y(n343) );
  AND2X2 U396 ( .A(\mem<11><7> ), .B(n1881), .Y(n344) );
  INVX1 U397 ( .A(n344), .Y(n345) );
  AND2X2 U398 ( .A(\mem<11><8> ), .B(n1882), .Y(n346) );
  INVX1 U399 ( .A(n346), .Y(n347) );
  AND2X2 U400 ( .A(\mem<11><9> ), .B(n1882), .Y(n348) );
  INVX1 U401 ( .A(n348), .Y(n349) );
  AND2X2 U402 ( .A(\mem<11><10> ), .B(n1882), .Y(n350) );
  INVX1 U403 ( .A(n350), .Y(n351) );
  AND2X2 U404 ( .A(\mem<11><11> ), .B(n1882), .Y(n352) );
  INVX1 U405 ( .A(n352), .Y(n353) );
  AND2X2 U406 ( .A(\mem<11><12> ), .B(n1882), .Y(n354) );
  INVX1 U407 ( .A(n354), .Y(n355) );
  AND2X2 U408 ( .A(\mem<11><13> ), .B(n1882), .Y(n356) );
  INVX1 U409 ( .A(n356), .Y(n357) );
  AND2X2 U410 ( .A(\mem<11><14> ), .B(n1882), .Y(n358) );
  INVX1 U411 ( .A(n358), .Y(n359) );
  AND2X2 U412 ( .A(\mem<11><15> ), .B(n1882), .Y(n360) );
  INVX1 U413 ( .A(n360), .Y(n361) );
  AND2X2 U414 ( .A(\mem<10><0> ), .B(n1883), .Y(n362) );
  INVX1 U415 ( .A(n362), .Y(n363) );
  AND2X2 U416 ( .A(\mem<10><1> ), .B(n1883), .Y(n364) );
  INVX1 U417 ( .A(n364), .Y(n365) );
  AND2X2 U418 ( .A(\mem<10><2> ), .B(n1883), .Y(n366) );
  INVX1 U419 ( .A(n366), .Y(n367) );
  AND2X2 U420 ( .A(\mem<10><3> ), .B(n1883), .Y(n368) );
  INVX1 U421 ( .A(n368), .Y(n369) );
  AND2X2 U422 ( .A(\mem<10><4> ), .B(n1883), .Y(n370) );
  INVX1 U423 ( .A(n370), .Y(n371) );
  AND2X2 U424 ( .A(\mem<10><5> ), .B(n1883), .Y(n372) );
  INVX1 U425 ( .A(n372), .Y(n373) );
  AND2X2 U426 ( .A(\mem<10><6> ), .B(n1883), .Y(n374) );
  INVX1 U427 ( .A(n374), .Y(n375) );
  AND2X2 U428 ( .A(\mem<10><7> ), .B(n1883), .Y(n376) );
  INVX1 U429 ( .A(n376), .Y(n377) );
  AND2X2 U430 ( .A(\mem<10><8> ), .B(n1884), .Y(n378) );
  INVX1 U431 ( .A(n378), .Y(n379) );
  AND2X2 U432 ( .A(\mem<10><9> ), .B(n1884), .Y(n380) );
  INVX1 U433 ( .A(n380), .Y(n381) );
  AND2X2 U434 ( .A(\mem<10><10> ), .B(n1884), .Y(n382) );
  INVX1 U435 ( .A(n382), .Y(n383) );
  AND2X2 U436 ( .A(\mem<10><11> ), .B(n1884), .Y(n384) );
  INVX1 U437 ( .A(n384), .Y(n385) );
  AND2X2 U438 ( .A(\mem<10><12> ), .B(n1884), .Y(n386) );
  INVX1 U439 ( .A(n386), .Y(n387) );
  AND2X2 U440 ( .A(\mem<10><13> ), .B(n1884), .Y(n388) );
  INVX1 U441 ( .A(n388), .Y(n389) );
  AND2X2 U442 ( .A(\mem<10><14> ), .B(n1884), .Y(n390) );
  INVX1 U443 ( .A(n390), .Y(n391) );
  AND2X2 U444 ( .A(\mem<10><15> ), .B(n1884), .Y(n392) );
  INVX1 U445 ( .A(n392), .Y(n393) );
  AND2X2 U446 ( .A(\mem<9><0> ), .B(n1885), .Y(n394) );
  INVX1 U447 ( .A(n394), .Y(n395) );
  AND2X2 U448 ( .A(\mem<9><1> ), .B(n1885), .Y(n396) );
  INVX1 U449 ( .A(n396), .Y(n397) );
  AND2X2 U450 ( .A(\mem<9><2> ), .B(n1885), .Y(n398) );
  INVX1 U451 ( .A(n398), .Y(n399) );
  AND2X2 U452 ( .A(\mem<9><3> ), .B(n1885), .Y(n400) );
  INVX1 U453 ( .A(n400), .Y(n401) );
  AND2X2 U454 ( .A(\mem<9><4> ), .B(n1885), .Y(n402) );
  INVX1 U455 ( .A(n402), .Y(n403) );
  AND2X2 U456 ( .A(\mem<9><5> ), .B(n1885), .Y(n404) );
  INVX1 U457 ( .A(n404), .Y(n405) );
  AND2X2 U458 ( .A(\mem<9><6> ), .B(n1885), .Y(n406) );
  INVX1 U459 ( .A(n406), .Y(n407) );
  AND2X2 U460 ( .A(\mem<9><7> ), .B(n1885), .Y(n408) );
  INVX1 U461 ( .A(n408), .Y(n409) );
  AND2X2 U462 ( .A(\mem<9><8> ), .B(n1886), .Y(n410) );
  INVX1 U463 ( .A(n410), .Y(n411) );
  AND2X2 U464 ( .A(\mem<9><9> ), .B(n1886), .Y(n412) );
  INVX1 U465 ( .A(n412), .Y(n413) );
  AND2X2 U466 ( .A(\mem<9><10> ), .B(n1886), .Y(n414) );
  INVX1 U467 ( .A(n414), .Y(n415) );
  AND2X2 U468 ( .A(\mem<9><11> ), .B(n1886), .Y(n416) );
  INVX1 U469 ( .A(n416), .Y(n417) );
  AND2X2 U470 ( .A(\mem<9><12> ), .B(n1886), .Y(n418) );
  INVX1 U471 ( .A(n418), .Y(n419) );
  AND2X2 U472 ( .A(\mem<9><13> ), .B(n1886), .Y(n420) );
  INVX1 U473 ( .A(n420), .Y(n421) );
  AND2X2 U474 ( .A(\mem<9><14> ), .B(n1886), .Y(n422) );
  INVX1 U475 ( .A(n422), .Y(n423) );
  AND2X2 U476 ( .A(\mem<9><15> ), .B(n1886), .Y(n424) );
  INVX1 U477 ( .A(n424), .Y(n425) );
  AND2X2 U478 ( .A(\mem<8><0> ), .B(n1888), .Y(n426) );
  INVX1 U479 ( .A(n426), .Y(n427) );
  AND2X2 U480 ( .A(\mem<8><1> ), .B(n1888), .Y(n428) );
  INVX1 U481 ( .A(n428), .Y(n429) );
  AND2X2 U482 ( .A(\mem<8><2> ), .B(n1888), .Y(n430) );
  INVX1 U483 ( .A(n430), .Y(n431) );
  AND2X2 U484 ( .A(\mem<8><3> ), .B(n1888), .Y(n432) );
  INVX1 U485 ( .A(n432), .Y(n433) );
  AND2X2 U486 ( .A(\mem<8><4> ), .B(n1888), .Y(n434) );
  INVX1 U487 ( .A(n434), .Y(n435) );
  AND2X2 U488 ( .A(\mem<8><5> ), .B(n1888), .Y(n436) );
  INVX1 U489 ( .A(n436), .Y(n437) );
  AND2X2 U490 ( .A(\mem<8><6> ), .B(n1888), .Y(n438) );
  INVX1 U491 ( .A(n438), .Y(n439) );
  AND2X2 U492 ( .A(\mem<8><7> ), .B(n1888), .Y(n440) );
  INVX1 U493 ( .A(n440), .Y(n441) );
  AND2X2 U494 ( .A(\mem<8><8> ), .B(n1889), .Y(n442) );
  INVX1 U495 ( .A(n442), .Y(n443) );
  AND2X2 U496 ( .A(\mem<8><9> ), .B(n1889), .Y(n444) );
  INVX1 U497 ( .A(n444), .Y(n445) );
  AND2X2 U498 ( .A(\mem<8><10> ), .B(n1889), .Y(n446) );
  INVX1 U499 ( .A(n446), .Y(n447) );
  AND2X2 U500 ( .A(\mem<8><11> ), .B(n1889), .Y(n448) );
  INVX1 U501 ( .A(n448), .Y(n449) );
  AND2X2 U502 ( .A(\mem<8><12> ), .B(n1889), .Y(n450) );
  INVX1 U503 ( .A(n450), .Y(n451) );
  AND2X2 U504 ( .A(\mem<8><13> ), .B(n1889), .Y(n452) );
  INVX1 U505 ( .A(n452), .Y(n453) );
  AND2X2 U506 ( .A(\mem<8><14> ), .B(n1889), .Y(n454) );
  INVX1 U507 ( .A(n454), .Y(n455) );
  AND2X2 U508 ( .A(\mem<8><15> ), .B(n1889), .Y(n456) );
  INVX1 U509 ( .A(n456), .Y(n457) );
  AND2X2 U510 ( .A(\mem<7><0> ), .B(n1890), .Y(n458) );
  INVX1 U511 ( .A(n458), .Y(n459) );
  AND2X2 U512 ( .A(\mem<7><1> ), .B(n1890), .Y(n460) );
  INVX1 U513 ( .A(n460), .Y(n461) );
  AND2X2 U514 ( .A(\mem<7><2> ), .B(n1890), .Y(n462) );
  INVX1 U515 ( .A(n462), .Y(n463) );
  AND2X2 U516 ( .A(\mem<7><3> ), .B(n1890), .Y(n464) );
  INVX1 U517 ( .A(n464), .Y(n465) );
  AND2X2 U518 ( .A(\mem<7><4> ), .B(n1890), .Y(n466) );
  INVX1 U519 ( .A(n466), .Y(n467) );
  AND2X2 U520 ( .A(\mem<7><5> ), .B(n1890), .Y(n468) );
  INVX1 U521 ( .A(n468), .Y(n469) );
  AND2X2 U522 ( .A(\mem<7><6> ), .B(n1890), .Y(n470) );
  INVX1 U523 ( .A(n470), .Y(n471) );
  AND2X2 U524 ( .A(\mem<7><7> ), .B(n1890), .Y(n472) );
  INVX1 U525 ( .A(n472), .Y(n473) );
  AND2X2 U526 ( .A(\mem<7><8> ), .B(n1891), .Y(n474) );
  INVX1 U527 ( .A(n474), .Y(n475) );
  AND2X2 U528 ( .A(\mem<7><9> ), .B(n1891), .Y(n476) );
  INVX1 U529 ( .A(n476), .Y(n477) );
  AND2X2 U530 ( .A(\mem<7><10> ), .B(n1891), .Y(n478) );
  INVX1 U531 ( .A(n478), .Y(n479) );
  AND2X2 U532 ( .A(\mem<7><11> ), .B(n1891), .Y(n480) );
  INVX1 U533 ( .A(n480), .Y(n481) );
  AND2X2 U534 ( .A(\mem<7><12> ), .B(n1891), .Y(n482) );
  INVX1 U535 ( .A(n482), .Y(n483) );
  AND2X2 U536 ( .A(\mem<7><13> ), .B(n1891), .Y(n484) );
  INVX1 U537 ( .A(n484), .Y(n485) );
  AND2X2 U538 ( .A(\mem<7><14> ), .B(n1891), .Y(n486) );
  INVX1 U539 ( .A(n486), .Y(n487) );
  AND2X2 U540 ( .A(\mem<7><15> ), .B(n1891), .Y(n488) );
  INVX1 U541 ( .A(n488), .Y(n489) );
  AND2X2 U542 ( .A(\mem<6><0> ), .B(n1892), .Y(n490) );
  INVX1 U543 ( .A(n490), .Y(n491) );
  AND2X2 U544 ( .A(\mem<6><1> ), .B(n1892), .Y(n492) );
  INVX1 U545 ( .A(n492), .Y(n493) );
  AND2X2 U546 ( .A(\mem<6><2> ), .B(n1892), .Y(n494) );
  INVX1 U547 ( .A(n494), .Y(n495) );
  AND2X2 U548 ( .A(\mem<6><3> ), .B(n1892), .Y(n496) );
  INVX1 U549 ( .A(n496), .Y(n497) );
  AND2X2 U550 ( .A(\mem<6><4> ), .B(n1892), .Y(n498) );
  INVX1 U551 ( .A(n498), .Y(n499) );
  AND2X2 U552 ( .A(\mem<6><5> ), .B(n1892), .Y(n500) );
  INVX1 U553 ( .A(n500), .Y(n501) );
  AND2X2 U554 ( .A(\mem<6><6> ), .B(n1892), .Y(n502) );
  INVX1 U555 ( .A(n502), .Y(n503) );
  AND2X2 U556 ( .A(\mem<6><7> ), .B(n1892), .Y(n504) );
  INVX1 U557 ( .A(n504), .Y(n505) );
  AND2X2 U558 ( .A(\mem<6><8> ), .B(n1893), .Y(n506) );
  INVX1 U559 ( .A(n506), .Y(n507) );
  AND2X2 U560 ( .A(\mem<6><9> ), .B(n1893), .Y(n508) );
  INVX1 U561 ( .A(n508), .Y(n509) );
  AND2X2 U562 ( .A(\mem<6><10> ), .B(n1893), .Y(n510) );
  INVX1 U563 ( .A(n510), .Y(n511) );
  AND2X2 U564 ( .A(\mem<6><11> ), .B(n1893), .Y(n512) );
  INVX1 U565 ( .A(n512), .Y(n513) );
  AND2X2 U566 ( .A(\mem<6><12> ), .B(n1893), .Y(n514) );
  INVX1 U567 ( .A(n514), .Y(n515) );
  AND2X2 U568 ( .A(\mem<6><13> ), .B(n1893), .Y(n516) );
  INVX1 U569 ( .A(n516), .Y(n517) );
  AND2X2 U570 ( .A(\mem<6><14> ), .B(n1893), .Y(n518) );
  INVX1 U571 ( .A(n518), .Y(n519) );
  AND2X2 U572 ( .A(\mem<6><15> ), .B(n1893), .Y(n520) );
  INVX1 U573 ( .A(n520), .Y(n521) );
  AND2X2 U574 ( .A(\mem<5><0> ), .B(n1894), .Y(n522) );
  INVX1 U575 ( .A(n522), .Y(n523) );
  AND2X2 U576 ( .A(\mem<5><1> ), .B(n1894), .Y(n524) );
  INVX1 U577 ( .A(n524), .Y(n525) );
  AND2X2 U578 ( .A(\mem<5><2> ), .B(n1894), .Y(n526) );
  INVX1 U579 ( .A(n526), .Y(n527) );
  AND2X2 U580 ( .A(\mem<5><3> ), .B(n1894), .Y(n528) );
  INVX1 U581 ( .A(n528), .Y(n529) );
  AND2X2 U582 ( .A(\mem<5><4> ), .B(n1894), .Y(n530) );
  INVX1 U583 ( .A(n530), .Y(n531) );
  AND2X2 U584 ( .A(\mem<5><5> ), .B(n1894), .Y(n532) );
  INVX1 U585 ( .A(n532), .Y(n533) );
  AND2X2 U586 ( .A(\mem<5><6> ), .B(n1894), .Y(n534) );
  INVX1 U587 ( .A(n534), .Y(n535) );
  AND2X2 U588 ( .A(\mem<5><7> ), .B(n1894), .Y(n536) );
  INVX1 U589 ( .A(n536), .Y(n537) );
  AND2X2 U590 ( .A(\mem<5><8> ), .B(n1895), .Y(n538) );
  INVX1 U591 ( .A(n538), .Y(n539) );
  AND2X2 U592 ( .A(\mem<5><9> ), .B(n1895), .Y(n540) );
  INVX1 U593 ( .A(n540), .Y(n541) );
  AND2X2 U594 ( .A(\mem<5><10> ), .B(n1895), .Y(n542) );
  INVX1 U595 ( .A(n542), .Y(n543) );
  AND2X2 U596 ( .A(\mem<5><11> ), .B(n1895), .Y(n544) );
  INVX1 U597 ( .A(n544), .Y(n545) );
  AND2X2 U598 ( .A(\mem<5><12> ), .B(n1895), .Y(n546) );
  INVX1 U599 ( .A(n546), .Y(n547) );
  AND2X2 U600 ( .A(\mem<5><13> ), .B(n1895), .Y(n548) );
  INVX1 U601 ( .A(n548), .Y(n549) );
  AND2X2 U602 ( .A(\mem<5><14> ), .B(n1895), .Y(n550) );
  INVX1 U603 ( .A(n550), .Y(n551) );
  AND2X2 U604 ( .A(\mem<5><15> ), .B(n1895), .Y(n552) );
  INVX1 U605 ( .A(n552), .Y(n553) );
  AND2X2 U606 ( .A(\mem<4><0> ), .B(n1896), .Y(n554) );
  INVX1 U607 ( .A(n554), .Y(n555) );
  AND2X2 U608 ( .A(\mem<4><1> ), .B(n1896), .Y(n556) );
  INVX1 U609 ( .A(n556), .Y(n557) );
  AND2X2 U610 ( .A(\mem<4><2> ), .B(n1896), .Y(n558) );
  INVX1 U611 ( .A(n558), .Y(n559) );
  AND2X2 U612 ( .A(\mem<4><3> ), .B(n1896), .Y(n560) );
  INVX1 U613 ( .A(n560), .Y(n561) );
  AND2X2 U614 ( .A(\mem<4><4> ), .B(n1896), .Y(n562) );
  INVX1 U615 ( .A(n562), .Y(n563) );
  AND2X2 U616 ( .A(\mem<4><5> ), .B(n1896), .Y(n564) );
  INVX1 U617 ( .A(n564), .Y(n565) );
  AND2X2 U618 ( .A(\mem<4><6> ), .B(n1896), .Y(n566) );
  INVX1 U619 ( .A(n566), .Y(n567) );
  AND2X2 U620 ( .A(\mem<4><7> ), .B(n1896), .Y(n568) );
  INVX1 U621 ( .A(n568), .Y(n569) );
  AND2X2 U622 ( .A(\mem<4><8> ), .B(n1897), .Y(n570) );
  INVX1 U623 ( .A(n570), .Y(n571) );
  AND2X2 U624 ( .A(\mem<4><9> ), .B(n1897), .Y(n572) );
  INVX1 U625 ( .A(n572), .Y(n573) );
  AND2X2 U626 ( .A(\mem<4><10> ), .B(n1897), .Y(n574) );
  INVX1 U627 ( .A(n574), .Y(n575) );
  AND2X2 U628 ( .A(\mem<4><11> ), .B(n1897), .Y(n576) );
  INVX1 U629 ( .A(n576), .Y(n577) );
  AND2X2 U630 ( .A(\mem<4><12> ), .B(n1897), .Y(n578) );
  INVX1 U631 ( .A(n578), .Y(n579) );
  AND2X2 U632 ( .A(\mem<4><13> ), .B(n1897), .Y(n580) );
  INVX1 U633 ( .A(n580), .Y(n581) );
  AND2X2 U634 ( .A(\mem<4><14> ), .B(n1897), .Y(n582) );
  INVX1 U635 ( .A(n582), .Y(n583) );
  AND2X2 U636 ( .A(\mem<4><15> ), .B(n1897), .Y(n584) );
  INVX1 U637 ( .A(n584), .Y(n585) );
  AND2X2 U638 ( .A(\mem<3><0> ), .B(n1898), .Y(n586) );
  INVX1 U639 ( .A(n586), .Y(n587) );
  AND2X2 U640 ( .A(\mem<3><1> ), .B(n1898), .Y(n588) );
  INVX1 U641 ( .A(n588), .Y(n589) );
  AND2X2 U642 ( .A(\mem<3><2> ), .B(n1898), .Y(n590) );
  INVX1 U643 ( .A(n590), .Y(n591) );
  AND2X2 U644 ( .A(\mem<3><3> ), .B(n1898), .Y(n592) );
  INVX1 U645 ( .A(n592), .Y(n593) );
  AND2X2 U646 ( .A(\mem<3><4> ), .B(n1898), .Y(n594) );
  INVX1 U647 ( .A(n594), .Y(n595) );
  AND2X2 U648 ( .A(\mem<3><5> ), .B(n1898), .Y(n596) );
  INVX1 U649 ( .A(n596), .Y(n597) );
  AND2X2 U650 ( .A(\mem<3><6> ), .B(n1898), .Y(n598) );
  INVX1 U651 ( .A(n598), .Y(n599) );
  AND2X2 U652 ( .A(\mem<3><7> ), .B(n1898), .Y(n600) );
  INVX1 U653 ( .A(n600), .Y(n601) );
  AND2X2 U654 ( .A(\mem<3><8> ), .B(n1899), .Y(n602) );
  INVX1 U655 ( .A(n602), .Y(n603) );
  AND2X2 U656 ( .A(\mem<3><9> ), .B(n1899), .Y(n604) );
  INVX1 U657 ( .A(n604), .Y(n605) );
  AND2X2 U658 ( .A(\mem<3><10> ), .B(n1899), .Y(n606) );
  INVX1 U659 ( .A(n606), .Y(n607) );
  AND2X2 U660 ( .A(\mem<3><11> ), .B(n1899), .Y(n608) );
  INVX1 U661 ( .A(n608), .Y(n609) );
  AND2X2 U662 ( .A(\mem<3><12> ), .B(n1899), .Y(n610) );
  INVX1 U663 ( .A(n610), .Y(n611) );
  AND2X2 U664 ( .A(\mem<3><13> ), .B(n1899), .Y(n612) );
  INVX1 U665 ( .A(n612), .Y(n613) );
  AND2X2 U666 ( .A(\mem<3><14> ), .B(n1899), .Y(n614) );
  INVX1 U667 ( .A(n614), .Y(n615) );
  AND2X2 U668 ( .A(\mem<3><15> ), .B(n1899), .Y(n616) );
  INVX1 U669 ( .A(n616), .Y(n617) );
  AND2X2 U670 ( .A(\mem<2><0> ), .B(n1900), .Y(n618) );
  INVX1 U671 ( .A(n618), .Y(n619) );
  AND2X2 U672 ( .A(\mem<2><1> ), .B(n1900), .Y(n620) );
  INVX1 U673 ( .A(n620), .Y(n621) );
  AND2X2 U674 ( .A(\mem<2><2> ), .B(n1900), .Y(n622) );
  INVX1 U675 ( .A(n622), .Y(n623) );
  AND2X2 U676 ( .A(\mem<2><3> ), .B(n1900), .Y(n624) );
  INVX1 U677 ( .A(n624), .Y(n625) );
  AND2X2 U678 ( .A(\mem<2><4> ), .B(n1900), .Y(n626) );
  INVX1 U679 ( .A(n626), .Y(n627) );
  AND2X2 U680 ( .A(\mem<2><5> ), .B(n1900), .Y(n628) );
  INVX1 U681 ( .A(n628), .Y(n629) );
  AND2X2 U682 ( .A(\mem<2><6> ), .B(n1900), .Y(n630) );
  INVX1 U683 ( .A(n630), .Y(n631) );
  AND2X2 U684 ( .A(\mem<2><7> ), .B(n1900), .Y(n632) );
  INVX1 U685 ( .A(n632), .Y(n633) );
  AND2X2 U686 ( .A(\mem<2><8> ), .B(n1901), .Y(n634) );
  INVX1 U687 ( .A(n634), .Y(n635) );
  AND2X2 U688 ( .A(\mem<2><9> ), .B(n1901), .Y(n636) );
  INVX1 U689 ( .A(n636), .Y(n637) );
  AND2X2 U690 ( .A(\mem<2><10> ), .B(n1901), .Y(n638) );
  INVX1 U691 ( .A(n638), .Y(n639) );
  AND2X2 U692 ( .A(\mem<2><11> ), .B(n1901), .Y(n640) );
  INVX1 U693 ( .A(n640), .Y(n641) );
  AND2X2 U694 ( .A(\mem<2><12> ), .B(n1901), .Y(n642) );
  INVX1 U695 ( .A(n642), .Y(n643) );
  AND2X2 U696 ( .A(\mem<2><13> ), .B(n1901), .Y(n644) );
  INVX1 U697 ( .A(n644), .Y(n645) );
  AND2X2 U698 ( .A(\mem<2><14> ), .B(n1901), .Y(n646) );
  INVX1 U699 ( .A(n646), .Y(n647) );
  AND2X2 U700 ( .A(\mem<2><15> ), .B(n1901), .Y(n648) );
  INVX1 U701 ( .A(n648), .Y(n649) );
  AND2X2 U702 ( .A(\mem<1><0> ), .B(n1902), .Y(n650) );
  INVX1 U703 ( .A(n650), .Y(n1163) );
  AND2X2 U704 ( .A(\mem<1><1> ), .B(n1902), .Y(n1164) );
  INVX1 U705 ( .A(n1164), .Y(n1165) );
  AND2X2 U706 ( .A(\mem<1><2> ), .B(n1902), .Y(n1166) );
  INVX1 U707 ( .A(n1166), .Y(n1167) );
  AND2X2 U708 ( .A(\mem<1><3> ), .B(n1902), .Y(n1168) );
  INVX1 U709 ( .A(n1168), .Y(n1169) );
  AND2X2 U710 ( .A(\mem<1><4> ), .B(n1902), .Y(n1170) );
  INVX1 U711 ( .A(n1170), .Y(n1171) );
  AND2X2 U712 ( .A(\mem<1><5> ), .B(n1902), .Y(n1172) );
  INVX1 U713 ( .A(n1172), .Y(n1173) );
  AND2X2 U714 ( .A(\mem<1><6> ), .B(n1902), .Y(n1174) );
  INVX1 U715 ( .A(n1174), .Y(n1175) );
  AND2X2 U716 ( .A(\mem<1><7> ), .B(n1902), .Y(n1176) );
  INVX1 U717 ( .A(n1176), .Y(n1177) );
  AND2X2 U718 ( .A(\mem<1><8> ), .B(n1903), .Y(n1178) );
  INVX1 U719 ( .A(n1178), .Y(n1179) );
  AND2X2 U720 ( .A(\mem<1><9> ), .B(n1903), .Y(n1180) );
  INVX1 U721 ( .A(n1180), .Y(n1181) );
  AND2X2 U722 ( .A(\mem<1><10> ), .B(n1903), .Y(n1182) );
  INVX1 U723 ( .A(n1182), .Y(n1183) );
  AND2X2 U724 ( .A(\mem<1><11> ), .B(n1903), .Y(n1184) );
  INVX1 U725 ( .A(n1184), .Y(n1185) );
  AND2X2 U726 ( .A(\mem<1><12> ), .B(n1903), .Y(n1186) );
  INVX1 U727 ( .A(n1186), .Y(n1187) );
  AND2X2 U728 ( .A(\mem<1><13> ), .B(n1903), .Y(n1188) );
  INVX1 U729 ( .A(n1188), .Y(n1189) );
  AND2X2 U730 ( .A(\mem<1><14> ), .B(n1903), .Y(n1190) );
  INVX1 U731 ( .A(n1190), .Y(n1191) );
  AND2X2 U732 ( .A(\mem<1><15> ), .B(n1903), .Y(n1192) );
  INVX1 U733 ( .A(n1192), .Y(n1193) );
  AND2X2 U734 ( .A(\mem<0><0> ), .B(n1905), .Y(n1194) );
  INVX1 U735 ( .A(n1194), .Y(n1195) );
  AND2X2 U736 ( .A(\mem<0><1> ), .B(n1905), .Y(n1196) );
  INVX1 U737 ( .A(n1196), .Y(n1197) );
  AND2X2 U738 ( .A(\mem<0><2> ), .B(n1905), .Y(n1198) );
  INVX1 U739 ( .A(n1198), .Y(n1199) );
  AND2X2 U740 ( .A(\mem<0><3> ), .B(n1905), .Y(n1200) );
  INVX1 U741 ( .A(n1200), .Y(n1201) );
  AND2X2 U742 ( .A(\mem<0><4> ), .B(n1905), .Y(n1202) );
  INVX1 U743 ( .A(n1202), .Y(n1203) );
  AND2X2 U744 ( .A(\mem<0><5> ), .B(n1905), .Y(n1204) );
  INVX1 U745 ( .A(n1204), .Y(n1205) );
  AND2X2 U746 ( .A(\mem<0><6> ), .B(n1905), .Y(n1206) );
  INVX1 U747 ( .A(n1206), .Y(n1207) );
  AND2X2 U748 ( .A(\mem<0><7> ), .B(n1905), .Y(n1208) );
  INVX1 U749 ( .A(n1208), .Y(n1209) );
  AND2X2 U750 ( .A(\mem<0><8> ), .B(n1906), .Y(n1210) );
  INVX1 U751 ( .A(n1210), .Y(n1211) );
  AND2X2 U752 ( .A(\mem<0><9> ), .B(n1906), .Y(n1212) );
  INVX1 U753 ( .A(n1212), .Y(n1213) );
  AND2X2 U754 ( .A(\mem<0><10> ), .B(n1906), .Y(n1214) );
  INVX1 U755 ( .A(n1214), .Y(n1215) );
  AND2X2 U756 ( .A(\mem<0><11> ), .B(n1906), .Y(n1216) );
  INVX1 U757 ( .A(n1216), .Y(n1217) );
  AND2X2 U758 ( .A(\mem<0><12> ), .B(n1906), .Y(n1218) );
  INVX1 U759 ( .A(n1218), .Y(n1219) );
  AND2X2 U760 ( .A(\mem<0><13> ), .B(n1906), .Y(n1220) );
  INVX1 U761 ( .A(n1220), .Y(n1221) );
  AND2X2 U762 ( .A(\mem<0><14> ), .B(n1906), .Y(n1222) );
  INVX1 U763 ( .A(n1222), .Y(n1223) );
  AND2X2 U764 ( .A(\mem<0><15> ), .B(n1906), .Y(n1224) );
  INVX1 U765 ( .A(n1224), .Y(n1225) );
  INVX1 U766 ( .A(n1948), .Y(n1947) );
  INVX1 U767 ( .A(n1946), .Y(n1945) );
  INVX1 U768 ( .A(n1951), .Y(n1950) );
  INVX1 U769 ( .A(N13), .Y(n1951) );
  AND2X1 U770 ( .A(n1825), .B(n1947), .Y(n1226) );
  AND2X1 U771 ( .A(n2672), .B(N14), .Y(n1227) );
  INVX2 U772 ( .A(n1911), .Y(n1907) );
  BUFX2 U773 ( .A(n34), .Y(n1864) );
  BUFX2 U774 ( .A(n34), .Y(n1865) );
  BUFX2 U775 ( .A(n36), .Y(n1866) );
  BUFX2 U776 ( .A(n36), .Y(n1867) );
  BUFX2 U777 ( .A(n38), .Y(n1868) );
  BUFX2 U778 ( .A(n38), .Y(n1869) );
  BUFX2 U779 ( .A(n40), .Y(n1871) );
  BUFX2 U780 ( .A(n40), .Y(n1872) );
  BUFX2 U781 ( .A(n42), .Y(n1873) );
  BUFX2 U782 ( .A(n42), .Y(n1874) );
  BUFX2 U783 ( .A(n44), .Y(n1875) );
  BUFX2 U784 ( .A(n44), .Y(n1876) );
  BUFX2 U785 ( .A(n46), .Y(n1877) );
  BUFX2 U786 ( .A(n46), .Y(n1878) );
  BUFX2 U787 ( .A(n48), .Y(n1879) );
  BUFX2 U788 ( .A(n48), .Y(n1880) );
  BUFX2 U789 ( .A(n50), .Y(n1881) );
  BUFX2 U790 ( .A(n50), .Y(n1882) );
  BUFX2 U791 ( .A(n52), .Y(n1883) );
  BUFX2 U792 ( .A(n52), .Y(n1884) );
  BUFX2 U793 ( .A(n54), .Y(n1885) );
  BUFX2 U794 ( .A(n54), .Y(n1886) );
  BUFX2 U795 ( .A(n56), .Y(n1888) );
  BUFX2 U796 ( .A(n56), .Y(n1889) );
  BUFX2 U797 ( .A(n58), .Y(n1890) );
  BUFX2 U798 ( .A(n58), .Y(n1891) );
  BUFX2 U799 ( .A(n60), .Y(n1892) );
  BUFX2 U800 ( .A(n60), .Y(n1893) );
  BUFX2 U801 ( .A(n62), .Y(n1894) );
  BUFX2 U802 ( .A(n62), .Y(n1895) );
  BUFX2 U803 ( .A(n64), .Y(n1896) );
  BUFX2 U804 ( .A(n64), .Y(n1897) );
  BUFX2 U805 ( .A(n66), .Y(n1898) );
  BUFX2 U806 ( .A(n66), .Y(n1899) );
  BUFX2 U807 ( .A(n68), .Y(n1900) );
  BUFX2 U808 ( .A(n68), .Y(n1901) );
  BUFX2 U809 ( .A(n70), .Y(n1902) );
  BUFX2 U810 ( .A(n70), .Y(n1903) );
  BUFX2 U811 ( .A(n72), .Y(n1905) );
  BUFX2 U812 ( .A(n72), .Y(n1906) );
  BUFX2 U813 ( .A(n1985), .Y(n1228) );
  INVX1 U814 ( .A(n1228), .Y(n2153) );
  BUFX2 U815 ( .A(n2002), .Y(n1229) );
  INVX1 U816 ( .A(n1229), .Y(n2154) );
  BUFX2 U817 ( .A(n2019), .Y(n1230) );
  INVX1 U818 ( .A(n1230), .Y(n2155) );
  BUFX2 U819 ( .A(n2036), .Y(n1231) );
  INVX1 U820 ( .A(n1231), .Y(n2156) );
  BUFX2 U821 ( .A(n2053), .Y(n1232) );
  INVX1 U822 ( .A(n1232), .Y(n2157) );
  BUFX2 U823 ( .A(n2150), .Y(n1233) );
  INVX1 U824 ( .A(n1233), .Y(n2151) );
  BUFX2 U825 ( .A(n2152), .Y(n1234) );
  INVX1 U826 ( .A(n1234), .Y(n2158) );
  AND2X1 U827 ( .A(n1945), .B(n1226), .Y(n1235) );
  AND2X1 U828 ( .A(n1950), .B(n1227), .Y(n1236) );
  INVX1 U829 ( .A(n4), .Y(n1911) );
  INVX4 U830 ( .A(n4), .Y(n1910) );
  AND2X1 U831 ( .A(n1946), .B(n1226), .Y(n1237) );
  AND2X1 U832 ( .A(n1951), .B(n1227), .Y(n1238) );
  AND2X1 U833 ( .A(n1236), .B(n2159), .Y(n1239) );
  AND2X1 U834 ( .A(n2159), .B(n1238), .Y(n1240) );
  AND2X1 U835 ( .A(n2159), .B(n2151), .Y(n1241) );
  AND2X1 U836 ( .A(n2159), .B(n2158), .Y(n1242) );
  AND2X1 U837 ( .A(n1235), .B(n1236), .Y(n1243) );
  INVX1 U838 ( .A(n1243), .Y(n1244) );
  INVX1 U839 ( .A(n6), .Y(n1245) );
  INVX1 U840 ( .A(n6), .Y(n1246) );
  AND2X1 U841 ( .A(n1236), .B(n1237), .Y(n1247) );
  INVX1 U842 ( .A(n1247), .Y(n1248) );
  INVX1 U843 ( .A(n22), .Y(n1249) );
  INVX1 U844 ( .A(n22), .Y(n1250) );
  AND2X1 U845 ( .A(n1236), .B(n2153), .Y(n1251) );
  INVX1 U846 ( .A(n1251), .Y(n1252) );
  INVX1 U847 ( .A(n23), .Y(n1253) );
  INVX1 U848 ( .A(n23), .Y(n1254) );
  AND2X1 U849 ( .A(n1236), .B(n2154), .Y(n1255) );
  INVX1 U850 ( .A(n1255), .Y(n1256) );
  INVX1 U851 ( .A(n24), .Y(n1257) );
  INVX1 U852 ( .A(n24), .Y(n1258) );
  AND2X1 U853 ( .A(n1236), .B(n2155), .Y(n1259) );
  INVX1 U854 ( .A(n1259), .Y(n1260) );
  INVX1 U855 ( .A(n25), .Y(n1261) );
  INVX1 U856 ( .A(n25), .Y(n1262) );
  AND2X1 U857 ( .A(n1236), .B(n2156), .Y(n1263) );
  INVX1 U858 ( .A(n1263), .Y(n1264) );
  INVX1 U859 ( .A(n26), .Y(n1265) );
  INVX1 U860 ( .A(n26), .Y(n1266) );
  AND2X1 U861 ( .A(n1236), .B(n2157), .Y(n1267) );
  INVX1 U862 ( .A(n1267), .Y(n1268) );
  INVX1 U863 ( .A(n27), .Y(n1269) );
  INVX1 U864 ( .A(n27), .Y(n1270) );
  INVX1 U865 ( .A(n28), .Y(n1271) );
  INVX1 U866 ( .A(n28), .Y(n1272) );
  AND2X1 U867 ( .A(n1235), .B(n1238), .Y(n1273) );
  INVX1 U868 ( .A(n1273), .Y(n1274) );
  INVX1 U869 ( .A(n29), .Y(n1275) );
  INVX1 U870 ( .A(n29), .Y(n1276) );
  AND2X1 U871 ( .A(n1237), .B(n1238), .Y(n1277) );
  INVX1 U872 ( .A(n1277), .Y(n1278) );
  INVX1 U873 ( .A(n30), .Y(n1279) );
  INVX1 U874 ( .A(n30), .Y(n1280) );
  AND2X1 U875 ( .A(n2153), .B(n1238), .Y(n1281) );
  INVX1 U876 ( .A(n1281), .Y(n1282) );
  INVX1 U877 ( .A(n31), .Y(n1283) );
  INVX1 U878 ( .A(n31), .Y(n1284) );
  AND2X1 U879 ( .A(n2154), .B(n1238), .Y(n1285) );
  INVX1 U880 ( .A(n1285), .Y(n1286) );
  INVX1 U881 ( .A(n32), .Y(n1287) );
  INVX1 U882 ( .A(n32), .Y(n1288) );
  AND2X1 U883 ( .A(n2155), .B(n1238), .Y(n1289) );
  INVX1 U884 ( .A(n1289), .Y(n1290) );
  AND2X1 U885 ( .A(n2156), .B(n1238), .Y(n1291) );
  INVX1 U886 ( .A(n1291), .Y(n1292) );
  AND2X1 U887 ( .A(n2157), .B(n1238), .Y(n1293) );
  INVX1 U888 ( .A(n1293), .Y(n1294) );
  AND2X1 U889 ( .A(n1235), .B(n2151), .Y(n1295) );
  INVX1 U890 ( .A(n1295), .Y(n1296) );
  AND2X1 U891 ( .A(n1237), .B(n2151), .Y(n1297) );
  INVX1 U892 ( .A(n1297), .Y(n1298) );
  AND2X1 U893 ( .A(n2153), .B(n2151), .Y(n1299) );
  INVX1 U894 ( .A(n1299), .Y(n1300) );
  AND2X1 U895 ( .A(n2154), .B(n2151), .Y(n1301) );
  INVX1 U896 ( .A(n1301), .Y(n1302) );
  AND2X1 U897 ( .A(n2155), .B(n2151), .Y(n1303) );
  INVX1 U898 ( .A(n1303), .Y(n1304) );
  AND2X1 U899 ( .A(n2156), .B(n2151), .Y(n1305) );
  INVX1 U900 ( .A(n1305), .Y(n1306) );
  AND2X1 U901 ( .A(n2157), .B(n2151), .Y(n1307) );
  INVX1 U902 ( .A(n1307), .Y(n1308) );
  AND2X1 U903 ( .A(n1235), .B(n2158), .Y(n1309) );
  INVX1 U904 ( .A(n1309), .Y(n1310) );
  AND2X1 U905 ( .A(n1237), .B(n2158), .Y(n1311) );
  INVX1 U906 ( .A(n1311), .Y(n1312) );
  AND2X1 U907 ( .A(n2153), .B(n2158), .Y(n1313) );
  INVX1 U908 ( .A(n1313), .Y(n1314) );
  AND2X1 U909 ( .A(n2154), .B(n2158), .Y(n1315) );
  INVX1 U910 ( .A(n1315), .Y(n1316) );
  AND2X1 U911 ( .A(n2155), .B(n2158), .Y(n1317) );
  INVX1 U912 ( .A(n1317), .Y(n1318) );
  AND2X1 U913 ( .A(n2156), .B(n2158), .Y(n1319) );
  INVX1 U914 ( .A(n1319), .Y(n1320) );
  AND2X1 U915 ( .A(n2157), .B(n2158), .Y(n1321) );
  INVX1 U916 ( .A(n1321), .Y(n1322) );
  MUX2X1 U917 ( .B(n1324), .A(n1325), .S(n1830), .Y(n1323) );
  MUX2X1 U918 ( .B(n1327), .A(n1328), .S(n1830), .Y(n1326) );
  MUX2X1 U919 ( .B(n1330), .A(n1331), .S(n1830), .Y(n1329) );
  MUX2X1 U920 ( .B(n1333), .A(n1334), .S(n1830), .Y(n1332) );
  MUX2X1 U921 ( .B(n1336), .A(n1337), .S(n1822), .Y(n1335) );
  MUX2X1 U922 ( .B(n1339), .A(n1340), .S(n1830), .Y(n1338) );
  MUX2X1 U923 ( .B(n1342), .A(n1343), .S(n1830), .Y(n1341) );
  MUX2X1 U924 ( .B(n1345), .A(n1346), .S(n1830), .Y(n1344) );
  MUX2X1 U925 ( .B(n1348), .A(n1349), .S(n1830), .Y(n1347) );
  MUX2X1 U926 ( .B(n1351), .A(n1352), .S(n1822), .Y(n1350) );
  MUX2X1 U927 ( .B(n1354), .A(n1355), .S(n1831), .Y(n1353) );
  MUX2X1 U928 ( .B(n1357), .A(n1358), .S(n1831), .Y(n1356) );
  MUX2X1 U929 ( .B(n1360), .A(n1361), .S(n1831), .Y(n1359) );
  MUX2X1 U930 ( .B(n1363), .A(n1364), .S(n1831), .Y(n1362) );
  MUX2X1 U931 ( .B(n1366), .A(n1367), .S(n1822), .Y(n1365) );
  MUX2X1 U932 ( .B(n1369), .A(n1370), .S(n1831), .Y(n1368) );
  MUX2X1 U933 ( .B(n1372), .A(n1373), .S(n1831), .Y(n1371) );
  MUX2X1 U934 ( .B(n1375), .A(n1376), .S(n1831), .Y(n1374) );
  MUX2X1 U935 ( .B(n1378), .A(n1379), .S(n1831), .Y(n1377) );
  MUX2X1 U936 ( .B(n1381), .A(n1382), .S(n1822), .Y(n1380) );
  MUX2X1 U937 ( .B(n1384), .A(n1385), .S(n1831), .Y(n1383) );
  MUX2X1 U938 ( .B(n1387), .A(n1388), .S(n1831), .Y(n1386) );
  MUX2X1 U939 ( .B(n1390), .A(n1391), .S(n1831), .Y(n1389) );
  MUX2X1 U940 ( .B(n1393), .A(n1394), .S(n1831), .Y(n1392) );
  MUX2X1 U941 ( .B(n1396), .A(n1397), .S(n1822), .Y(n1395) );
  MUX2X1 U942 ( .B(n1399), .A(n1400), .S(n1832), .Y(n1398) );
  MUX2X1 U943 ( .B(n1402), .A(n1403), .S(n1832), .Y(n1401) );
  MUX2X1 U944 ( .B(n1405), .A(n1406), .S(n1832), .Y(n1404) );
  MUX2X1 U945 ( .B(n1408), .A(n1409), .S(n1832), .Y(n1407) );
  MUX2X1 U946 ( .B(n1411), .A(n1412), .S(n1822), .Y(n1410) );
  MUX2X1 U947 ( .B(n1414), .A(n1415), .S(n1832), .Y(n1413) );
  MUX2X1 U948 ( .B(n1417), .A(n1418), .S(n1832), .Y(n1416) );
  MUX2X1 U949 ( .B(n1420), .A(n1421), .S(n1832), .Y(n1419) );
  MUX2X1 U950 ( .B(n1423), .A(n1424), .S(n1832), .Y(n1422) );
  MUX2X1 U951 ( .B(n1426), .A(n1427), .S(n1822), .Y(n1425) );
  MUX2X1 U952 ( .B(n1429), .A(n1430), .S(n1832), .Y(n1428) );
  MUX2X1 U953 ( .B(n1432), .A(n1433), .S(n1832), .Y(n1431) );
  MUX2X1 U954 ( .B(n1435), .A(n1436), .S(n1832), .Y(n1434) );
  MUX2X1 U955 ( .B(n1438), .A(n1439), .S(n1832), .Y(n1437) );
  MUX2X1 U956 ( .B(n1441), .A(n1442), .S(n1822), .Y(n1440) );
  MUX2X1 U957 ( .B(n1444), .A(n1445), .S(n1833), .Y(n1443) );
  MUX2X1 U958 ( .B(n1447), .A(n1448), .S(n1833), .Y(n1446) );
  MUX2X1 U959 ( .B(n1450), .A(n1451), .S(n1833), .Y(n1449) );
  MUX2X1 U960 ( .B(n1453), .A(n1454), .S(n1833), .Y(n1452) );
  MUX2X1 U961 ( .B(n1456), .A(n1457), .S(n1822), .Y(n1455) );
  MUX2X1 U962 ( .B(n1459), .A(n1460), .S(n1833), .Y(n1458) );
  MUX2X1 U963 ( .B(n1462), .A(n1463), .S(n1833), .Y(n1461) );
  MUX2X1 U964 ( .B(n1465), .A(n1466), .S(n1833), .Y(n1464) );
  MUX2X1 U965 ( .B(n1468), .A(n1469), .S(n1833), .Y(n1467) );
  MUX2X1 U966 ( .B(n1471), .A(n1472), .S(n1822), .Y(n1470) );
  MUX2X1 U967 ( .B(n1474), .A(n1475), .S(n1833), .Y(n1473) );
  MUX2X1 U968 ( .B(n1477), .A(n1478), .S(n1833), .Y(n1476) );
  MUX2X1 U969 ( .B(n1480), .A(n1481), .S(n1833), .Y(n1479) );
  MUX2X1 U970 ( .B(n1483), .A(n1484), .S(n1833), .Y(n1482) );
  MUX2X1 U971 ( .B(n1486), .A(n1487), .S(n1822), .Y(n1485) );
  MUX2X1 U972 ( .B(n1489), .A(n1490), .S(n1834), .Y(n1488) );
  MUX2X1 U973 ( .B(n1492), .A(n1493), .S(n1834), .Y(n1491) );
  MUX2X1 U974 ( .B(n1495), .A(n1496), .S(n1834), .Y(n1494) );
  MUX2X1 U975 ( .B(n1498), .A(n1499), .S(n1834), .Y(n1497) );
  MUX2X1 U976 ( .B(n1501), .A(n1502), .S(n1822), .Y(n1500) );
  MUX2X1 U977 ( .B(n1504), .A(n1505), .S(n1834), .Y(n1503) );
  MUX2X1 U978 ( .B(n1507), .A(n1508), .S(n1834), .Y(n1506) );
  MUX2X1 U979 ( .B(n1510), .A(n1511), .S(n1834), .Y(n1509) );
  MUX2X1 U980 ( .B(n1513), .A(n1514), .S(n1834), .Y(n1512) );
  MUX2X1 U981 ( .B(n1516), .A(n1517), .S(n1821), .Y(n1515) );
  MUX2X1 U982 ( .B(n1519), .A(n1520), .S(n1834), .Y(n1518) );
  MUX2X1 U983 ( .B(n1522), .A(n1523), .S(n1834), .Y(n1521) );
  MUX2X1 U984 ( .B(n1525), .A(n1526), .S(n1834), .Y(n1524) );
  MUX2X1 U985 ( .B(n1528), .A(n1529), .S(n1834), .Y(n1527) );
  MUX2X1 U986 ( .B(n1531), .A(n1532), .S(n1821), .Y(n1530) );
  MUX2X1 U987 ( .B(n1534), .A(n1535), .S(n1835), .Y(n1533) );
  MUX2X1 U988 ( .B(n1537), .A(n1538), .S(n1835), .Y(n1536) );
  MUX2X1 U989 ( .B(n1540), .A(n1541), .S(n1835), .Y(n1539) );
  MUX2X1 U990 ( .B(n1543), .A(n1544), .S(n1835), .Y(n1542) );
  MUX2X1 U991 ( .B(n1546), .A(n1547), .S(n1821), .Y(n1545) );
  MUX2X1 U992 ( .B(n1549), .A(n1550), .S(n1835), .Y(n1548) );
  MUX2X1 U993 ( .B(n1552), .A(n1553), .S(n1835), .Y(n1551) );
  MUX2X1 U994 ( .B(n1555), .A(n1556), .S(n1835), .Y(n1554) );
  MUX2X1 U995 ( .B(n1558), .A(n1559), .S(n1835), .Y(n1557) );
  MUX2X1 U996 ( .B(n1561), .A(n1562), .S(n1821), .Y(n1560) );
  MUX2X1 U997 ( .B(n1564), .A(n1565), .S(n1835), .Y(n1563) );
  MUX2X1 U998 ( .B(n1567), .A(n1568), .S(n1835), .Y(n1566) );
  MUX2X1 U999 ( .B(n1570), .A(n1571), .S(n1835), .Y(n1569) );
  MUX2X1 U1000 ( .B(n1573), .A(n1574), .S(n1835), .Y(n1572) );
  MUX2X1 U1001 ( .B(n1576), .A(n1577), .S(n1821), .Y(n1575) );
  MUX2X1 U1002 ( .B(n1579), .A(n1580), .S(n1836), .Y(n1578) );
  MUX2X1 U1003 ( .B(n1582), .A(n1583), .S(n1836), .Y(n1581) );
  MUX2X1 U1004 ( .B(n1585), .A(n1586), .S(n1836), .Y(n1584) );
  MUX2X1 U1005 ( .B(n1588), .A(n1589), .S(n1836), .Y(n1587) );
  MUX2X1 U1006 ( .B(n1591), .A(n1592), .S(n1821), .Y(n1590) );
  MUX2X1 U1007 ( .B(n1594), .A(n1595), .S(n1836), .Y(n1593) );
  MUX2X1 U1008 ( .B(n1597), .A(n1598), .S(n1836), .Y(n1596) );
  MUX2X1 U1009 ( .B(n1600), .A(n1601), .S(n1836), .Y(n1599) );
  MUX2X1 U1010 ( .B(n1603), .A(n1604), .S(n1836), .Y(n1602) );
  MUX2X1 U1011 ( .B(n1606), .A(n1607), .S(n1821), .Y(n1605) );
  MUX2X1 U1012 ( .B(n1609), .A(n1610), .S(n1836), .Y(n1608) );
  MUX2X1 U1013 ( .B(n1612), .A(n1613), .S(n1836), .Y(n1611) );
  MUX2X1 U1014 ( .B(n1615), .A(n1616), .S(n1836), .Y(n1614) );
  MUX2X1 U1015 ( .B(n1618), .A(n1619), .S(n1836), .Y(n1617) );
  MUX2X1 U1016 ( .B(n1621), .A(n1622), .S(n1821), .Y(n1620) );
  MUX2X1 U1017 ( .B(n1624), .A(n1625), .S(n1837), .Y(n1623) );
  MUX2X1 U1018 ( .B(n1627), .A(n1628), .S(n1837), .Y(n1626) );
  MUX2X1 U1019 ( .B(n1630), .A(n1631), .S(n1837), .Y(n1629) );
  MUX2X1 U1020 ( .B(n1633), .A(n1634), .S(n1837), .Y(n1632) );
  MUX2X1 U1021 ( .B(n1636), .A(n1637), .S(n1821), .Y(n1635) );
  MUX2X1 U1022 ( .B(n1639), .A(n1640), .S(n1837), .Y(n1638) );
  MUX2X1 U1023 ( .B(n1642), .A(n1643), .S(n1837), .Y(n1641) );
  MUX2X1 U1024 ( .B(n1645), .A(n1646), .S(n1837), .Y(n1644) );
  MUX2X1 U1025 ( .B(n1648), .A(n1649), .S(n1837), .Y(n1647) );
  MUX2X1 U1026 ( .B(n1651), .A(n1652), .S(n1821), .Y(n1650) );
  MUX2X1 U1027 ( .B(n1654), .A(n1655), .S(n1837), .Y(n1653) );
  MUX2X1 U1028 ( .B(n1657), .A(n1658), .S(n1837), .Y(n1656) );
  MUX2X1 U1029 ( .B(n1660), .A(n1661), .S(n1837), .Y(n1659) );
  MUX2X1 U1030 ( .B(n1663), .A(n1664), .S(n1837), .Y(n1662) );
  MUX2X1 U1031 ( .B(n1666), .A(n1667), .S(n1821), .Y(n1665) );
  MUX2X1 U1032 ( .B(n1669), .A(n1670), .S(n1838), .Y(n1668) );
  MUX2X1 U1033 ( .B(n1672), .A(n1673), .S(n1838), .Y(n1671) );
  MUX2X1 U1034 ( .B(n1675), .A(n1676), .S(n1838), .Y(n1674) );
  MUX2X1 U1035 ( .B(n1678), .A(n1679), .S(n1838), .Y(n1677) );
  MUX2X1 U1036 ( .B(n1681), .A(n1682), .S(n1821), .Y(n1680) );
  MUX2X1 U1037 ( .B(n1684), .A(n1685), .S(n1838), .Y(n1683) );
  MUX2X1 U1038 ( .B(n1687), .A(n1688), .S(n1838), .Y(n1686) );
  MUX2X1 U1039 ( .B(n1690), .A(n1691), .S(n1838), .Y(n1689) );
  MUX2X1 U1040 ( .B(n1693), .A(n1694), .S(n1838), .Y(n1692) );
  MUX2X1 U1041 ( .B(n1696), .A(n1697), .S(n1820), .Y(n1695) );
  MUX2X1 U1042 ( .B(n1699), .A(n1700), .S(n1838), .Y(n1698) );
  MUX2X1 U1043 ( .B(n1702), .A(n1703), .S(n1838), .Y(n1701) );
  MUX2X1 U1044 ( .B(n1705), .A(n1706), .S(n1838), .Y(n1704) );
  MUX2X1 U1045 ( .B(n1708), .A(n1709), .S(n1838), .Y(n1707) );
  MUX2X1 U1046 ( .B(n1711), .A(n1712), .S(n1820), .Y(n1710) );
  MUX2X1 U1047 ( .B(n1714), .A(n1715), .S(n1839), .Y(n1713) );
  MUX2X1 U1048 ( .B(n1717), .A(n1718), .S(n1839), .Y(n1716) );
  MUX2X1 U1049 ( .B(n1720), .A(n1721), .S(n1839), .Y(n1719) );
  MUX2X1 U1050 ( .B(n1723), .A(n1724), .S(n1839), .Y(n1722) );
  MUX2X1 U1051 ( .B(n1726), .A(n1727), .S(n1820), .Y(n1725) );
  MUX2X1 U1052 ( .B(n1729), .A(n1730), .S(n1839), .Y(n1728) );
  MUX2X1 U1053 ( .B(n1732), .A(n1733), .S(n1839), .Y(n1731) );
  MUX2X1 U1054 ( .B(n1735), .A(n1736), .S(n1839), .Y(n1734) );
  MUX2X1 U1055 ( .B(n1738), .A(n1739), .S(n1839), .Y(n1737) );
  MUX2X1 U1056 ( .B(n1741), .A(n1742), .S(n1820), .Y(n1740) );
  MUX2X1 U1057 ( .B(n1744), .A(n1745), .S(n1839), .Y(n1743) );
  MUX2X1 U1058 ( .B(n1747), .A(n1748), .S(n1839), .Y(n1746) );
  MUX2X1 U1059 ( .B(n1750), .A(n1751), .S(n1839), .Y(n1749) );
  MUX2X1 U1060 ( .B(n1753), .A(n1754), .S(n1839), .Y(n1752) );
  MUX2X1 U1061 ( .B(n1756), .A(n1757), .S(n1820), .Y(n1755) );
  MUX2X1 U1062 ( .B(n1759), .A(n1760), .S(n1840), .Y(n1758) );
  MUX2X1 U1063 ( .B(n1762), .A(n1763), .S(n1840), .Y(n1761) );
  MUX2X1 U1064 ( .B(n1765), .A(n1766), .S(n1840), .Y(n1764) );
  MUX2X1 U1065 ( .B(n1768), .A(n1769), .S(n1840), .Y(n1767) );
  MUX2X1 U1066 ( .B(n1771), .A(n1772), .S(n1820), .Y(n1770) );
  MUX2X1 U1067 ( .B(n1774), .A(n1775), .S(n1840), .Y(n1773) );
  MUX2X1 U1068 ( .B(n1777), .A(n1778), .S(n1840), .Y(n1776) );
  MUX2X1 U1069 ( .B(n1780), .A(n1781), .S(n1840), .Y(n1779) );
  MUX2X1 U1070 ( .B(n1783), .A(n1784), .S(n1840), .Y(n1782) );
  MUX2X1 U1071 ( .B(n1786), .A(n1787), .S(n1820), .Y(n1785) );
  MUX2X1 U1072 ( .B(n1789), .A(n1790), .S(n1840), .Y(n1788) );
  MUX2X1 U1073 ( .B(n1792), .A(n1793), .S(n1840), .Y(n1791) );
  MUX2X1 U1074 ( .B(n1795), .A(n1796), .S(n1840), .Y(n1794) );
  MUX2X1 U1075 ( .B(n1798), .A(n1799), .S(n1840), .Y(n1797) );
  MUX2X1 U1076 ( .B(n1801), .A(n1802), .S(n1820), .Y(n1800) );
  MUX2X1 U1077 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1851), .Y(n1325) );
  MUX2X1 U1078 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1855), .Y(n1324) );
  MUX2X1 U1079 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1855), .Y(n1328) );
  MUX2X1 U1080 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1855), .Y(n1327) );
  MUX2X1 U1081 ( .B(n1326), .A(n1323), .S(n1827), .Y(n1337) );
  MUX2X1 U1082 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1844), .Y(n1331) );
  MUX2X1 U1083 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1844), .Y(n1330) );
  MUX2X1 U1084 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1844), .Y(n1334) );
  MUX2X1 U1085 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1844), .Y(n1333) );
  MUX2X1 U1086 ( .B(n1332), .A(n1329), .S(n1827), .Y(n1336) );
  MUX2X1 U1087 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1844), .Y(n1340) );
  MUX2X1 U1088 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1844), .Y(n1339) );
  MUX2X1 U1089 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1844), .Y(n1343) );
  MUX2X1 U1090 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1844), .Y(n1342) );
  MUX2X1 U1091 ( .B(n1341), .A(n1338), .S(n1827), .Y(n1352) );
  MUX2X1 U1092 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1844), .Y(n1346) );
  MUX2X1 U1093 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1844), .Y(n1345) );
  MUX2X1 U1094 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1844), .Y(n1349) );
  MUX2X1 U1095 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1844), .Y(n1348) );
  MUX2X1 U1096 ( .B(n1347), .A(n1344), .S(n1827), .Y(n1351) );
  MUX2X1 U1097 ( .B(n1350), .A(n1335), .S(n1819), .Y(n1803) );
  MUX2X1 U1098 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1845), .Y(n1355) );
  MUX2X1 U1099 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1845), .Y(n1354) );
  MUX2X1 U1100 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1845), .Y(n1358) );
  MUX2X1 U1101 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1845), .Y(n1357) );
  MUX2X1 U1102 ( .B(n1356), .A(n1353), .S(n1827), .Y(n1367) );
  MUX2X1 U1103 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1845), .Y(n1361) );
  MUX2X1 U1104 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1845), .Y(n1360) );
  MUX2X1 U1105 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1845), .Y(n1364) );
  MUX2X1 U1106 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1845), .Y(n1363) );
  MUX2X1 U1107 ( .B(n1362), .A(n1359), .S(n1827), .Y(n1366) );
  MUX2X1 U1108 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1845), .Y(n1370) );
  MUX2X1 U1109 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1845), .Y(n1369) );
  MUX2X1 U1110 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1845), .Y(n1373) );
  MUX2X1 U1111 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1845), .Y(n1372) );
  MUX2X1 U1112 ( .B(n1371), .A(n1368), .S(n1827), .Y(n1382) );
  MUX2X1 U1113 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1846), .Y(n1376) );
  MUX2X1 U1114 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1846), .Y(n1375) );
  MUX2X1 U1115 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1846), .Y(n1379) );
  MUX2X1 U1116 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1846), .Y(n1378) );
  MUX2X1 U1117 ( .B(n1377), .A(n1374), .S(n1827), .Y(n1381) );
  MUX2X1 U1118 ( .B(n1380), .A(n1365), .S(n1819), .Y(n1804) );
  MUX2X1 U1119 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1846), .Y(n1385) );
  MUX2X1 U1120 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1846), .Y(n1384) );
  MUX2X1 U1121 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1846), .Y(n1388) );
  MUX2X1 U1122 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1846), .Y(n1387) );
  MUX2X1 U1123 ( .B(n1386), .A(n1383), .S(n1827), .Y(n1397) );
  MUX2X1 U1124 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1846), .Y(n1391) );
  MUX2X1 U1125 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1846), .Y(n1390) );
  MUX2X1 U1126 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1846), .Y(n1394) );
  MUX2X1 U1127 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1846), .Y(n1393) );
  MUX2X1 U1128 ( .B(n1392), .A(n1389), .S(n1827), .Y(n1396) );
  MUX2X1 U1129 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1847), .Y(n1400) );
  MUX2X1 U1130 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1847), .Y(n1399) );
  MUX2X1 U1131 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1847), .Y(n1403) );
  MUX2X1 U1132 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1847), .Y(n1402) );
  MUX2X1 U1133 ( .B(n1401), .A(n1398), .S(n1827), .Y(n1412) );
  MUX2X1 U1134 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1847), .Y(n1406) );
  MUX2X1 U1135 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1847), .Y(n1405) );
  MUX2X1 U1136 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1847), .Y(n1409) );
  MUX2X1 U1137 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1847), .Y(n1408) );
  MUX2X1 U1138 ( .B(n1407), .A(n1404), .S(n1827), .Y(n1411) );
  MUX2X1 U1139 ( .B(n1410), .A(n1395), .S(n1819), .Y(n1805) );
  MUX2X1 U1140 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1847), .Y(n1415) );
  MUX2X1 U1141 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1847), .Y(n1414) );
  MUX2X1 U1142 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1847), .Y(n1418) );
  MUX2X1 U1143 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1847), .Y(n1417) );
  MUX2X1 U1144 ( .B(n1416), .A(n1413), .S(n1826), .Y(n1427) );
  MUX2X1 U1145 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1853), .Y(n1421) );
  MUX2X1 U1146 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1856), .Y(n1420) );
  MUX2X1 U1147 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1853), .Y(n1424) );
  MUX2X1 U1148 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1848), .Y(n1423) );
  MUX2X1 U1149 ( .B(n1422), .A(n1419), .S(n1826), .Y(n1426) );
  MUX2X1 U1150 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1853), .Y(n1430) );
  MUX2X1 U1151 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1848), .Y(n1429) );
  MUX2X1 U1152 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1848), .Y(n1433) );
  MUX2X1 U1153 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1848), .Y(n1432) );
  MUX2X1 U1154 ( .B(n1431), .A(n1428), .S(n1826), .Y(n1442) );
  MUX2X1 U1155 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1854), .Y(n1436) );
  MUX2X1 U1156 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1854), .Y(n1435) );
  MUX2X1 U1157 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1848), .Y(n1439) );
  MUX2X1 U1158 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1848), .Y(n1438) );
  MUX2X1 U1159 ( .B(n1437), .A(n1434), .S(n1826), .Y(n1441) );
  MUX2X1 U1160 ( .B(n1440), .A(n1425), .S(n1819), .Y(n1806) );
  MUX2X1 U1161 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1848), .Y(n1445) );
  MUX2X1 U1162 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1848), .Y(n1444) );
  MUX2X1 U1163 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1848), .Y(n1448) );
  MUX2X1 U1164 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1848), .Y(n1447) );
  MUX2X1 U1165 ( .B(n1446), .A(n1443), .S(n1826), .Y(n1457) );
  MUX2X1 U1166 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1848), .Y(n1451) );
  MUX2X1 U1167 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1848), .Y(n1450) );
  MUX2X1 U1168 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1848), .Y(n1454) );
  MUX2X1 U1169 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1848), .Y(n1453) );
  MUX2X1 U1170 ( .B(n1452), .A(n1449), .S(n1826), .Y(n1456) );
  MUX2X1 U1171 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1848), .Y(n1460) );
  MUX2X1 U1172 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1848), .Y(n1459) );
  MUX2X1 U1173 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1848), .Y(n1463) );
  MUX2X1 U1174 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1848), .Y(n1462) );
  MUX2X1 U1175 ( .B(n1461), .A(n1458), .S(n1826), .Y(n1472) );
  MUX2X1 U1177 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1849), .Y(n1466) );
  MUX2X1 U1178 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1849), .Y(n1465) );
  MUX2X1 U1179 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1849), .Y(n1469) );
  MUX2X1 U1180 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1849), .Y(n1468) );
  MUX2X1 U1181 ( .B(n1467), .A(n1464), .S(n1826), .Y(n1471) );
  MUX2X1 U1182 ( .B(n1470), .A(n1455), .S(n1819), .Y(n1807) );
  MUX2X1 U1183 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1849), .Y(n1475) );
  MUX2X1 U1184 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1849), .Y(n1474) );
  MUX2X1 U1185 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1849), .Y(n1478) );
  MUX2X1 U1186 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1849), .Y(n1477) );
  MUX2X1 U1187 ( .B(n1476), .A(n1473), .S(n1826), .Y(n1487) );
  MUX2X1 U1188 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1849), .Y(n1481) );
  MUX2X1 U1189 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1849), .Y(n1480) );
  MUX2X1 U1190 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1849), .Y(n1484) );
  MUX2X1 U1191 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1849), .Y(n1483) );
  MUX2X1 U1192 ( .B(n1482), .A(n1479), .S(n1826), .Y(n1486) );
  MUX2X1 U1193 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1850), .Y(n1490) );
  MUX2X1 U1194 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1850), .Y(n1489) );
  MUX2X1 U1195 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1850), .Y(n1493) );
  MUX2X1 U1196 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1850), .Y(n1492) );
  MUX2X1 U1197 ( .B(n1491), .A(n1488), .S(n1826), .Y(n1502) );
  MUX2X1 U1198 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1850), .Y(n1496) );
  MUX2X1 U1199 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1850), .Y(n1495) );
  MUX2X1 U1200 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1850), .Y(n1499) );
  MUX2X1 U1201 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1850), .Y(n1498) );
  MUX2X1 U1202 ( .B(n1497), .A(n1494), .S(n1826), .Y(n1501) );
  MUX2X1 U1203 ( .B(n1500), .A(n1485), .S(n1819), .Y(n1808) );
  MUX2X1 U1204 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1850), .Y(n1505) );
  MUX2X1 U1205 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1850), .Y(n1504) );
  MUX2X1 U1206 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1850), .Y(n1508) );
  MUX2X1 U1207 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1850), .Y(n1507) );
  MUX2X1 U1208 ( .B(n1506), .A(n1503), .S(n1825), .Y(n1517) );
  MUX2X1 U1209 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1851), .Y(n1511) );
  MUX2X1 U1210 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1851), .Y(n1510) );
  MUX2X1 U1211 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1851), .Y(n1514) );
  MUX2X1 U1212 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1851), .Y(n1513) );
  MUX2X1 U1213 ( .B(n1512), .A(n1509), .S(n1825), .Y(n1516) );
  MUX2X1 U1214 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1851), .Y(n1520) );
  MUX2X1 U1215 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1851), .Y(n1519) );
  MUX2X1 U1216 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1851), .Y(n1523) );
  MUX2X1 U1217 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1851), .Y(n1522) );
  MUX2X1 U1218 ( .B(n1521), .A(n1518), .S(n1825), .Y(n1532) );
  MUX2X1 U1219 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1851), .Y(n1526) );
  MUX2X1 U1220 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1851), .Y(n1525) );
  MUX2X1 U1221 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1851), .Y(n1529) );
  MUX2X1 U1222 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1851), .Y(n1528) );
  MUX2X1 U1223 ( .B(n1527), .A(n1524), .S(n1825), .Y(n1531) );
  MUX2X1 U1224 ( .B(n1530), .A(n1515), .S(n1819), .Y(n1809) );
  MUX2X1 U1225 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1852), .Y(n1535) );
  MUX2X1 U1226 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1852), .Y(n1534) );
  MUX2X1 U1227 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1852), .Y(n1538) );
  MUX2X1 U1228 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1852), .Y(n1537) );
  MUX2X1 U1229 ( .B(n1536), .A(n1533), .S(n1825), .Y(n1547) );
  MUX2X1 U1230 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1852), .Y(n1541) );
  MUX2X1 U1231 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1852), .Y(n1540) );
  MUX2X1 U1232 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1852), .Y(n1544) );
  MUX2X1 U1233 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1852), .Y(n1543) );
  MUX2X1 U1234 ( .B(n1542), .A(n1539), .S(n1825), .Y(n1546) );
  MUX2X1 U1235 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1852), .Y(n1550) );
  MUX2X1 U1236 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1852), .Y(n1549) );
  MUX2X1 U1237 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1852), .Y(n1553) );
  MUX2X1 U1238 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1852), .Y(n1552) );
  MUX2X1 U1239 ( .B(n1551), .A(n1548), .S(n1825), .Y(n1562) );
  MUX2X1 U1240 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1853), .Y(n1556) );
  MUX2X1 U1241 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1853), .Y(n1555) );
  MUX2X1 U1242 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1853), .Y(n1559) );
  MUX2X1 U1243 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1853), .Y(n1558) );
  MUX2X1 U1244 ( .B(n1557), .A(n1554), .S(n1825), .Y(n1561) );
  MUX2X1 U1245 ( .B(n1560), .A(n1545), .S(n1819), .Y(n1810) );
  MUX2X1 U1246 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1853), .Y(n1565) );
  MUX2X1 U1247 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1853), .Y(n1564) );
  MUX2X1 U1248 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1853), .Y(n1568) );
  MUX2X1 U1249 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1853), .Y(n1567) );
  MUX2X1 U1250 ( .B(n1566), .A(n1563), .S(n1825), .Y(n1577) );
  MUX2X1 U1251 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1853), .Y(n1571) );
  MUX2X1 U1252 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1853), .Y(n1570) );
  MUX2X1 U1253 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1853), .Y(n1574) );
  MUX2X1 U1254 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1853), .Y(n1573) );
  MUX2X1 U1255 ( .B(n1572), .A(n1569), .S(n1825), .Y(n1576) );
  MUX2X1 U1256 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1854), .Y(n1580) );
  MUX2X1 U1257 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1854), .Y(n1579) );
  MUX2X1 U1258 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1854), .Y(n1583) );
  MUX2X1 U1259 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1854), .Y(n1582) );
  MUX2X1 U1260 ( .B(n1581), .A(n1578), .S(n1825), .Y(n1592) );
  MUX2X1 U1261 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1854), .Y(n1586) );
  MUX2X1 U1262 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1854), .Y(n1585) );
  MUX2X1 U1263 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1854), .Y(n1589) );
  MUX2X1 U1264 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1854), .Y(n1588) );
  MUX2X1 U1265 ( .B(n1587), .A(n1584), .S(n1825), .Y(n1591) );
  MUX2X1 U1266 ( .B(n1590), .A(n1575), .S(n1819), .Y(n1811) );
  MUX2X1 U1267 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1854), .Y(n1595) );
  MUX2X1 U1268 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1854), .Y(n1594) );
  MUX2X1 U1269 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1854), .Y(n1598) );
  MUX2X1 U1270 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1854), .Y(n1597) );
  MUX2X1 U1271 ( .B(n1596), .A(n1593), .S(n1824), .Y(n1607) );
  MUX2X1 U1272 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1855), .Y(n1601) );
  MUX2X1 U1273 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1855), .Y(n1600) );
  MUX2X1 U1274 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1855), .Y(n1604) );
  MUX2X1 U1275 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1855), .Y(n1603) );
  MUX2X1 U1276 ( .B(n1602), .A(n1599), .S(n1824), .Y(n1606) );
  MUX2X1 U1277 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1855), .Y(n1610) );
  MUX2X1 U1278 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1855), .Y(n1609) );
  MUX2X1 U1279 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1855), .Y(n1613) );
  MUX2X1 U1280 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1855), .Y(n1612) );
  MUX2X1 U1281 ( .B(n1611), .A(n1608), .S(n1824), .Y(n1622) );
  MUX2X1 U1282 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1855), .Y(n1616) );
  MUX2X1 U1283 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1855), .Y(n1615) );
  MUX2X1 U1284 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1855), .Y(n1619) );
  MUX2X1 U1285 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1855), .Y(n1618) );
  MUX2X1 U1286 ( .B(n1617), .A(n1614), .S(n1824), .Y(n1621) );
  MUX2X1 U1287 ( .B(n1620), .A(n1605), .S(n1819), .Y(n1812) );
  MUX2X1 U1288 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1856), .Y(n1625) );
  MUX2X1 U1289 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1856), .Y(n1624) );
  MUX2X1 U1290 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1856), .Y(n1628) );
  MUX2X1 U1291 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1856), .Y(n1627) );
  MUX2X1 U1292 ( .B(n1626), .A(n1623), .S(n1824), .Y(n1637) );
  MUX2X1 U1293 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1856), .Y(n1631) );
  MUX2X1 U1294 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1856), .Y(n1630) );
  MUX2X1 U1295 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1856), .Y(n1634) );
  MUX2X1 U1296 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1856), .Y(n1633) );
  MUX2X1 U1297 ( .B(n1632), .A(n1629), .S(n1824), .Y(n1636) );
  MUX2X1 U1298 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1856), .Y(n1640) );
  MUX2X1 U1299 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1856), .Y(n1639) );
  MUX2X1 U1300 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1856), .Y(n1643) );
  MUX2X1 U1301 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1856), .Y(n1642) );
  MUX2X1 U1302 ( .B(n1641), .A(n1638), .S(n1824), .Y(n1652) );
  MUX2X1 U1303 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1857), .Y(n1646) );
  MUX2X1 U1304 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1857), .Y(n1645) );
  MUX2X1 U1305 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1857), .Y(n1649) );
  MUX2X1 U1306 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1857), .Y(n1648) );
  MUX2X1 U1307 ( .B(n1647), .A(n1644), .S(n1824), .Y(n1651) );
  MUX2X1 U1308 ( .B(n1650), .A(n1635), .S(n1819), .Y(n1813) );
  MUX2X1 U1309 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1857), .Y(n1655) );
  MUX2X1 U1310 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1857), .Y(n1654) );
  MUX2X1 U1311 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1857), .Y(n1658) );
  MUX2X1 U1312 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1857), .Y(n1657) );
  MUX2X1 U1313 ( .B(n1656), .A(n1653), .S(n1824), .Y(n1667) );
  MUX2X1 U1314 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1857), .Y(n1661) );
  MUX2X1 U1315 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1857), .Y(n1660) );
  MUX2X1 U1316 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1857), .Y(n1664) );
  MUX2X1 U1317 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1857), .Y(n1663) );
  MUX2X1 U1318 ( .B(n1662), .A(n1659), .S(n1824), .Y(n1666) );
  MUX2X1 U1319 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1858), .Y(n1670) );
  MUX2X1 U1320 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1858), .Y(n1669) );
  MUX2X1 U1321 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1858), .Y(n1673) );
  MUX2X1 U1322 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1858), .Y(n1672) );
  MUX2X1 U1323 ( .B(n1671), .A(n1668), .S(n1824), .Y(n1682) );
  MUX2X1 U1324 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1858), .Y(n1676) );
  MUX2X1 U1325 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1858), .Y(n1675) );
  MUX2X1 U1326 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1858), .Y(n1679) );
  MUX2X1 U1327 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1858), .Y(n1678) );
  MUX2X1 U1328 ( .B(n1677), .A(n1674), .S(n1824), .Y(n1681) );
  MUX2X1 U1329 ( .B(n1680), .A(n1665), .S(n1819), .Y(n1814) );
  MUX2X1 U1330 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1858), .Y(n1685) );
  MUX2X1 U1331 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1858), .Y(n1684) );
  MUX2X1 U1332 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1858), .Y(n1688) );
  MUX2X1 U1333 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1858), .Y(n1687) );
  MUX2X1 U1334 ( .B(n1686), .A(n1683), .S(n1823), .Y(n1697) );
  MUX2X1 U1335 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1859), .Y(n1691) );
  MUX2X1 U1336 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1859), .Y(n1690) );
  MUX2X1 U1337 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1859), .Y(n1694) );
  MUX2X1 U1338 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1859), .Y(n1693) );
  MUX2X1 U1339 ( .B(n1692), .A(n1689), .S(n1823), .Y(n1696) );
  MUX2X1 U1340 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1859), .Y(n1700) );
  MUX2X1 U1341 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1859), .Y(n1699) );
  MUX2X1 U1342 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1859), .Y(n1703) );
  MUX2X1 U1343 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1859), .Y(n1702) );
  MUX2X1 U1344 ( .B(n1701), .A(n1698), .S(n1823), .Y(n1712) );
  MUX2X1 U1345 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1859), .Y(n1706) );
  MUX2X1 U1346 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1859), .Y(n1705) );
  MUX2X1 U1347 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1859), .Y(n1709) );
  MUX2X1 U1348 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1859), .Y(n1708) );
  MUX2X1 U1349 ( .B(n1707), .A(n1704), .S(n1823), .Y(n1711) );
  MUX2X1 U1350 ( .B(n1710), .A(n1695), .S(n1819), .Y(n1815) );
  MUX2X1 U1351 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1848), .Y(n1715) );
  MUX2X1 U1352 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1847), .Y(n1714) );
  MUX2X1 U1353 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1853), .Y(n1718) );
  MUX2X1 U1354 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1849), .Y(n1717) );
  MUX2X1 U1355 ( .B(n1716), .A(n1713), .S(n1823), .Y(n1727) );
  MUX2X1 U1356 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1860), .Y(n1721) );
  MUX2X1 U1357 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1849), .Y(n1720) );
  MUX2X1 U1358 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1848), .Y(n1724) );
  MUX2X1 U1359 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1849), .Y(n1723) );
  MUX2X1 U1360 ( .B(n1722), .A(n1719), .S(n1823), .Y(n1726) );
  MUX2X1 U1361 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1850), .Y(n1730) );
  MUX2X1 U1362 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1847), .Y(n1729) );
  MUX2X1 U1363 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1862), .Y(n1733) );
  MUX2X1 U1364 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1846), .Y(n1732) );
  MUX2X1 U1365 ( .B(n1731), .A(n1728), .S(n1823), .Y(n1742) );
  MUX2X1 U1366 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1861), .Y(n1736) );
  MUX2X1 U1367 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1848), .Y(n1735) );
  MUX2X1 U1368 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1848), .Y(n1739) );
  MUX2X1 U1369 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1847), .Y(n1738) );
  MUX2X1 U1370 ( .B(n1737), .A(n1734), .S(n1823), .Y(n1741) );
  MUX2X1 U1371 ( .B(n1740), .A(n1725), .S(n1819), .Y(n1816) );
  MUX2X1 U1372 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1848), .Y(n1745) );
  MUX2X1 U1373 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1849), .Y(n1744) );
  MUX2X1 U1374 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1850), .Y(n1748) );
  MUX2X1 U1375 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1850), .Y(n1747) );
  MUX2X1 U1376 ( .B(n1746), .A(n1743), .S(n1823), .Y(n1757) );
  MUX2X1 U1377 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1850), .Y(n1751) );
  MUX2X1 U1378 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1847), .Y(n1750) );
  MUX2X1 U1379 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1849), .Y(n1754) );
  MUX2X1 U1380 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1849), .Y(n1753) );
  MUX2X1 U1381 ( .B(n1752), .A(n1749), .S(n1823), .Y(n1756) );
  MUX2X1 U1382 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1860), .Y(n1760) );
  MUX2X1 U1383 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1860), .Y(n1759) );
  MUX2X1 U1384 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1860), .Y(n1763) );
  MUX2X1 U1385 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1860), .Y(n1762) );
  MUX2X1 U1386 ( .B(n1761), .A(n1758), .S(n1823), .Y(n1772) );
  MUX2X1 U1387 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1860), .Y(n1766) );
  MUX2X1 U1388 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1860), .Y(n1765) );
  MUX2X1 U1389 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1860), .Y(n1769) );
  MUX2X1 U1390 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1860), .Y(n1768) );
  MUX2X1 U1391 ( .B(n1767), .A(n1764), .S(n1823), .Y(n1771) );
  MUX2X1 U1392 ( .B(n1770), .A(n1755), .S(n1819), .Y(n1817) );
  MUX2X1 U1393 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1860), .Y(n1775) );
  MUX2X1 U1394 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1860), .Y(n1774) );
  MUX2X1 U1395 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1860), .Y(n1778) );
  MUX2X1 U1396 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1860), .Y(n1777) );
  MUX2X1 U1397 ( .B(n1776), .A(n1773), .S(n1823), .Y(n1787) );
  MUX2X1 U1398 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1861), .Y(n1781) );
  MUX2X1 U1399 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1861), .Y(n1780) );
  MUX2X1 U1400 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1861), .Y(n1784) );
  MUX2X1 U1401 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1861), .Y(n1783) );
  MUX2X1 U1402 ( .B(n1782), .A(n1779), .S(n1823), .Y(n1786) );
  MUX2X1 U1403 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1861), .Y(n1790) );
  MUX2X1 U1404 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1861), .Y(n1789) );
  MUX2X1 U1405 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1861), .Y(n1793) );
  MUX2X1 U1406 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1861), .Y(n1792) );
  MUX2X1 U1407 ( .B(n1791), .A(n1788), .S(n1824), .Y(n1802) );
  MUX2X1 U1408 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1861), .Y(n1796) );
  MUX2X1 U1409 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1861), .Y(n1795) );
  MUX2X1 U1410 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1861), .Y(n1799) );
  MUX2X1 U1411 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1861), .Y(n1798) );
  MUX2X1 U1412 ( .B(n1797), .A(n1794), .S(n1823), .Y(n1801) );
  MUX2X1 U1413 ( .B(n1800), .A(n1785), .S(n1819), .Y(n1818) );
  INVX8 U1414 ( .A(n1828), .Y(n1833) );
  INVX8 U1415 ( .A(n1828), .Y(n1834) );
  INVX8 U1416 ( .A(n1828), .Y(n1835) );
  INVX8 U1417 ( .A(n1828), .Y(n1836) );
  INVX8 U1418 ( .A(n1828), .Y(n1837) );
  INVX8 U1419 ( .A(n1828), .Y(n1838) );
  INVX8 U1420 ( .A(n1828), .Y(n1840) );
  INVX8 U1421 ( .A(n1842), .Y(n1844) );
  INVX8 U1422 ( .A(n1842), .Y(n1845) );
  INVX8 U1423 ( .A(n1843), .Y(n1847) );
  INVX8 U1424 ( .A(n1842), .Y(n1854) );
  INVX8 U1425 ( .A(n1842), .Y(n1857) );
  INVX8 U1426 ( .A(n1842), .Y(n1858) );
  INVX8 U1427 ( .A(n1842), .Y(n1859) );
  INVX1 U1428 ( .A(N12), .Y(n1949) );
  INVX1 U1429 ( .A(N11), .Y(n1948) );
  INVX1 U1430 ( .A(N10), .Y(n1946) );
  INVX8 U1431 ( .A(n1910), .Y(n1908) );
  INVX8 U1432 ( .A(n1910), .Y(n1909) );
  INVX8 U1433 ( .A(n5), .Y(n1912) );
  INVX8 U1434 ( .A(n5), .Y(n1913) );
  INVX8 U1435 ( .A(n7), .Y(n1914) );
  INVX8 U1436 ( .A(n7), .Y(n1915) );
  INVX8 U1437 ( .A(n8), .Y(n1916) );
  INVX8 U1438 ( .A(n8), .Y(n1917) );
  INVX8 U1439 ( .A(n9), .Y(n1918) );
  INVX8 U1440 ( .A(n9), .Y(n1919) );
  INVX8 U1441 ( .A(n10), .Y(n1920) );
  INVX8 U1442 ( .A(n10), .Y(n1921) );
  INVX8 U1443 ( .A(n11), .Y(n1922) );
  INVX8 U1444 ( .A(n11), .Y(n1923) );
  INVX8 U1445 ( .A(n12), .Y(n1924) );
  INVX8 U1446 ( .A(n12), .Y(n1925) );
  INVX8 U1447 ( .A(n13), .Y(n1926) );
  INVX8 U1448 ( .A(n13), .Y(n1927) );
  INVX8 U1449 ( .A(n14), .Y(n1928) );
  INVX8 U1450 ( .A(n14), .Y(n1929) );
  INVX8 U1451 ( .A(n15), .Y(n1930) );
  INVX8 U1452 ( .A(n15), .Y(n1931) );
  INVX8 U1453 ( .A(n16), .Y(n1932) );
  INVX8 U1454 ( .A(n16), .Y(n1933) );
  INVX8 U1455 ( .A(n17), .Y(n1934) );
  INVX8 U1456 ( .A(n17), .Y(n1935) );
  INVX8 U1457 ( .A(n18), .Y(n1936) );
  INVX8 U1458 ( .A(n18), .Y(n1937) );
  INVX8 U1459 ( .A(n19), .Y(n1938) );
  INVX8 U1460 ( .A(n19), .Y(n1939) );
  INVX8 U1461 ( .A(n20), .Y(n1940) );
  INVX8 U1462 ( .A(n20), .Y(n1941) );
  INVX8 U1463 ( .A(n21), .Y(n1942) );
  INVX8 U1464 ( .A(n21), .Y(n1943) );
  AND2X2 U1465 ( .A(N32), .B(n1), .Y(\data_out<0> ) );
  AND2X2 U1466 ( .A(n1), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U1467 ( .A(N30), .B(n1), .Y(\data_out<2> ) );
  AND2X2 U1468 ( .A(N29), .B(n1), .Y(\data_out<3> ) );
  AND2X2 U1469 ( .A(N28), .B(n1), .Y(\data_out<4> ) );
  AND2X2 U1470 ( .A(N27), .B(n3), .Y(\data_out<5> ) );
  AND2X2 U1471 ( .A(N26), .B(n3), .Y(\data_out<6> ) );
  AND2X2 U1472 ( .A(N25), .B(n3), .Y(\data_out<7> ) );
  AND2X2 U1473 ( .A(N24), .B(n1), .Y(\data_out<8> ) );
  AND2X2 U1474 ( .A(N23), .B(n3), .Y(\data_out<9> ) );
  AND2X2 U1475 ( .A(N22), .B(n3), .Y(\data_out<10> ) );
  AND2X2 U1476 ( .A(N21), .B(n3), .Y(\data_out<11> ) );
  AND2X2 U1477 ( .A(N20), .B(n1), .Y(\data_out<12> ) );
  AND2X2 U1478 ( .A(N19), .B(n3), .Y(\data_out<13> ) );
  AND2X2 U1479 ( .A(N18), .B(n3), .Y(\data_out<14> ) );
  AND2X2 U1480 ( .A(n1), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U1481 ( .A(\mem<31><0> ), .B(n1245), .Y(n1953) );
  OAI21X1 U1482 ( .A(n1244), .B(n1912), .C(n1953), .Y(n2671) );
  NAND2X1 U1483 ( .A(\mem<31><1> ), .B(n1245), .Y(n1954) );
  OAI21X1 U1484 ( .A(n1915), .B(n1244), .C(n1954), .Y(n2670) );
  NAND2X1 U1485 ( .A(\mem<31><2> ), .B(n1245), .Y(n1955) );
  OAI21X1 U1486 ( .A(n1917), .B(n1244), .C(n1955), .Y(n2669) );
  NAND2X1 U1487 ( .A(\mem<31><3> ), .B(n1245), .Y(n1956) );
  OAI21X1 U1488 ( .A(n1919), .B(n1244), .C(n1956), .Y(n2668) );
  NAND2X1 U1489 ( .A(\mem<31><4> ), .B(n1245), .Y(n1957) );
  OAI21X1 U1490 ( .A(n1921), .B(n1244), .C(n1957), .Y(n2667) );
  NAND2X1 U1491 ( .A(\mem<31><5> ), .B(n1245), .Y(n1958) );
  OAI21X1 U1492 ( .A(n1923), .B(n1244), .C(n1958), .Y(n2666) );
  NAND2X1 U1493 ( .A(\mem<31><6> ), .B(n1245), .Y(n1959) );
  OAI21X1 U1494 ( .A(n1925), .B(n1244), .C(n1959), .Y(n2665) );
  NAND2X1 U1495 ( .A(\mem<31><7> ), .B(n1245), .Y(n1960) );
  OAI21X1 U1496 ( .A(n1927), .B(n1244), .C(n1960), .Y(n2664) );
  NAND2X1 U1497 ( .A(\mem<31><8> ), .B(n1246), .Y(n1961) );
  OAI21X1 U1498 ( .A(n1929), .B(n1244), .C(n1961), .Y(n2663) );
  NAND2X1 U1499 ( .A(\mem<31><9> ), .B(n1246), .Y(n1962) );
  OAI21X1 U1500 ( .A(n1931), .B(n1244), .C(n1962), .Y(n2662) );
  NAND2X1 U1501 ( .A(\mem<31><10> ), .B(n1246), .Y(n1963) );
  OAI21X1 U1502 ( .A(n1933), .B(n1244), .C(n1963), .Y(n2661) );
  NAND2X1 U1503 ( .A(\mem<31><11> ), .B(n1246), .Y(n1964) );
  OAI21X1 U1504 ( .A(n1935), .B(n1244), .C(n1964), .Y(n2660) );
  NAND2X1 U1505 ( .A(\mem<31><12> ), .B(n1246), .Y(n1965) );
  OAI21X1 U1506 ( .A(n1937), .B(n1244), .C(n1965), .Y(n2659) );
  NAND2X1 U1507 ( .A(\mem<31><13> ), .B(n1246), .Y(n1966) );
  OAI21X1 U1508 ( .A(n1939), .B(n1244), .C(n1966), .Y(n2658) );
  NAND2X1 U1509 ( .A(\mem<31><14> ), .B(n1246), .Y(n1967) );
  OAI21X1 U1510 ( .A(n1941), .B(n1244), .C(n1967), .Y(n2657) );
  NAND2X1 U1511 ( .A(\mem<31><15> ), .B(n1246), .Y(n1968) );
  OAI21X1 U1512 ( .A(n1943), .B(n1244), .C(n1968), .Y(n2656) );
  NAND2X1 U1513 ( .A(\mem<30><0> ), .B(n1250), .Y(n1969) );
  OAI21X1 U1514 ( .A(n1248), .B(n1912), .C(n1969), .Y(n2655) );
  NAND2X1 U1515 ( .A(\mem<30><1> ), .B(n1250), .Y(n1970) );
  OAI21X1 U1516 ( .A(n1248), .B(n1915), .C(n1970), .Y(n2654) );
  NAND2X1 U1517 ( .A(\mem<30><2> ), .B(n1250), .Y(n1971) );
  OAI21X1 U1518 ( .A(n1248), .B(n1917), .C(n1971), .Y(n2653) );
  NAND2X1 U1519 ( .A(\mem<30><3> ), .B(n1250), .Y(n1972) );
  OAI21X1 U1520 ( .A(n1248), .B(n1919), .C(n1972), .Y(n2652) );
  NAND2X1 U1521 ( .A(\mem<30><4> ), .B(n1250), .Y(n1973) );
  OAI21X1 U1522 ( .A(n1248), .B(n1921), .C(n1973), .Y(n2651) );
  NAND2X1 U1523 ( .A(\mem<30><5> ), .B(n1250), .Y(n1974) );
  OAI21X1 U1524 ( .A(n1248), .B(n1923), .C(n1974), .Y(n2650) );
  NAND2X1 U1525 ( .A(\mem<30><6> ), .B(n1250), .Y(n1975) );
  OAI21X1 U1526 ( .A(n1248), .B(n1925), .C(n1975), .Y(n2649) );
  NAND2X1 U1527 ( .A(\mem<30><7> ), .B(n1250), .Y(n1976) );
  OAI21X1 U1528 ( .A(n1248), .B(n1927), .C(n1976), .Y(n2648) );
  NAND2X1 U1529 ( .A(\mem<30><8> ), .B(n1249), .Y(n1977) );
  OAI21X1 U1530 ( .A(n1248), .B(n1928), .C(n1977), .Y(n2647) );
  NAND2X1 U1531 ( .A(\mem<30><9> ), .B(n1249), .Y(n1978) );
  OAI21X1 U1532 ( .A(n1248), .B(n1930), .C(n1978), .Y(n2646) );
  NAND2X1 U1533 ( .A(\mem<30><10> ), .B(n1249), .Y(n1979) );
  OAI21X1 U1534 ( .A(n1248), .B(n1932), .C(n1979), .Y(n2645) );
  NAND2X1 U1535 ( .A(\mem<30><11> ), .B(n1249), .Y(n1980) );
  OAI21X1 U1536 ( .A(n1248), .B(n1934), .C(n1980), .Y(n2644) );
  NAND2X1 U1537 ( .A(\mem<30><12> ), .B(n1249), .Y(n1981) );
  OAI21X1 U1538 ( .A(n1248), .B(n1936), .C(n1981), .Y(n2643) );
  NAND2X1 U1539 ( .A(\mem<30><13> ), .B(n1249), .Y(n1982) );
  OAI21X1 U1540 ( .A(n1248), .B(n1938), .C(n1982), .Y(n2642) );
  NAND2X1 U1541 ( .A(\mem<30><14> ), .B(n1249), .Y(n1983) );
  OAI21X1 U1542 ( .A(n1248), .B(n1940), .C(n1983), .Y(n2641) );
  NAND2X1 U1543 ( .A(\mem<30><15> ), .B(n1249), .Y(n1984) );
  OAI21X1 U1544 ( .A(n1248), .B(n1942), .C(n1984), .Y(n2640) );
  NAND3X1 U1545 ( .A(n1945), .B(n1825), .C(n1948), .Y(n1985) );
  NAND2X1 U1546 ( .A(\mem<29><0> ), .B(n1254), .Y(n1986) );
  OAI21X1 U1547 ( .A(n1252), .B(n1912), .C(n1986), .Y(n2639) );
  NAND2X1 U1548 ( .A(\mem<29><1> ), .B(n1254), .Y(n1987) );
  OAI21X1 U1549 ( .A(n1252), .B(n1914), .C(n1987), .Y(n2638) );
  NAND2X1 U1550 ( .A(\mem<29><2> ), .B(n1254), .Y(n1988) );
  OAI21X1 U1551 ( .A(n1252), .B(n1916), .C(n1988), .Y(n2637) );
  NAND2X1 U1552 ( .A(\mem<29><3> ), .B(n1254), .Y(n1989) );
  OAI21X1 U1553 ( .A(n1252), .B(n1918), .C(n1989), .Y(n2636) );
  NAND2X1 U1554 ( .A(\mem<29><4> ), .B(n1254), .Y(n1990) );
  OAI21X1 U1555 ( .A(n1252), .B(n1920), .C(n1990), .Y(n2635) );
  NAND2X1 U1556 ( .A(\mem<29><5> ), .B(n1254), .Y(n1991) );
  OAI21X1 U1557 ( .A(n1252), .B(n1922), .C(n1991), .Y(n2634) );
  NAND2X1 U1558 ( .A(\mem<29><6> ), .B(n1254), .Y(n1992) );
  OAI21X1 U1559 ( .A(n1252), .B(n1924), .C(n1992), .Y(n2633) );
  NAND2X1 U1560 ( .A(\mem<29><7> ), .B(n1254), .Y(n1993) );
  OAI21X1 U1561 ( .A(n1252), .B(n1926), .C(n1993), .Y(n2632) );
  NAND2X1 U1562 ( .A(\mem<29><8> ), .B(n1253), .Y(n1994) );
  OAI21X1 U1563 ( .A(n1252), .B(n1929), .C(n1994), .Y(n2631) );
  NAND2X1 U1564 ( .A(\mem<29><9> ), .B(n1253), .Y(n1995) );
  OAI21X1 U1565 ( .A(n1252), .B(n1931), .C(n1995), .Y(n2630) );
  NAND2X1 U1566 ( .A(\mem<29><10> ), .B(n1253), .Y(n1996) );
  OAI21X1 U1567 ( .A(n1252), .B(n1933), .C(n1996), .Y(n2629) );
  NAND2X1 U1568 ( .A(\mem<29><11> ), .B(n1253), .Y(n1997) );
  OAI21X1 U1569 ( .A(n1252), .B(n1935), .C(n1997), .Y(n2628) );
  NAND2X1 U1570 ( .A(\mem<29><12> ), .B(n1253), .Y(n1998) );
  OAI21X1 U1571 ( .A(n1252), .B(n1937), .C(n1998), .Y(n2627) );
  NAND2X1 U1572 ( .A(\mem<29><13> ), .B(n1253), .Y(n1999) );
  OAI21X1 U1573 ( .A(n1252), .B(n1939), .C(n1999), .Y(n2626) );
  NAND2X1 U1574 ( .A(\mem<29><14> ), .B(n1253), .Y(n2000) );
  OAI21X1 U1575 ( .A(n1252), .B(n1941), .C(n2000), .Y(n2625) );
  NAND2X1 U1576 ( .A(\mem<29><15> ), .B(n1253), .Y(n2001) );
  OAI21X1 U1577 ( .A(n1252), .B(n1943), .C(n2001), .Y(n2624) );
  NAND3X1 U1578 ( .A(n1826), .B(n1948), .C(n1946), .Y(n2002) );
  NAND2X1 U1579 ( .A(\mem<28><0> ), .B(n1258), .Y(n2003) );
  OAI21X1 U1580 ( .A(n1256), .B(n1912), .C(n2003), .Y(n2623) );
  NAND2X1 U1581 ( .A(\mem<28><1> ), .B(n1258), .Y(n2004) );
  OAI21X1 U1582 ( .A(n1256), .B(n1915), .C(n2004), .Y(n2622) );
  NAND2X1 U1583 ( .A(\mem<28><2> ), .B(n1258), .Y(n2005) );
  OAI21X1 U1584 ( .A(n1256), .B(n1917), .C(n2005), .Y(n2621) );
  NAND2X1 U1585 ( .A(\mem<28><3> ), .B(n1258), .Y(n2006) );
  OAI21X1 U1586 ( .A(n1256), .B(n1919), .C(n2006), .Y(n2620) );
  NAND2X1 U1587 ( .A(\mem<28><4> ), .B(n1258), .Y(n2007) );
  OAI21X1 U1588 ( .A(n1256), .B(n1921), .C(n2007), .Y(n2619) );
  NAND2X1 U1589 ( .A(\mem<28><5> ), .B(n1258), .Y(n2008) );
  OAI21X1 U1590 ( .A(n1256), .B(n1923), .C(n2008), .Y(n2618) );
  NAND2X1 U1591 ( .A(\mem<28><6> ), .B(n1258), .Y(n2009) );
  OAI21X1 U1592 ( .A(n1256), .B(n1925), .C(n2009), .Y(n2617) );
  NAND2X1 U1593 ( .A(\mem<28><7> ), .B(n1258), .Y(n2010) );
  OAI21X1 U1594 ( .A(n1256), .B(n1927), .C(n2010), .Y(n2616) );
  NAND2X1 U1595 ( .A(\mem<28><8> ), .B(n1257), .Y(n2011) );
  OAI21X1 U1596 ( .A(n1256), .B(n1928), .C(n2011), .Y(n2615) );
  NAND2X1 U1597 ( .A(\mem<28><9> ), .B(n1257), .Y(n2012) );
  OAI21X1 U1598 ( .A(n1256), .B(n1930), .C(n2012), .Y(n2614) );
  NAND2X1 U1599 ( .A(\mem<28><10> ), .B(n1257), .Y(n2013) );
  OAI21X1 U1600 ( .A(n1256), .B(n1932), .C(n2013), .Y(n2613) );
  NAND2X1 U1601 ( .A(\mem<28><11> ), .B(n1257), .Y(n2014) );
  OAI21X1 U1602 ( .A(n1256), .B(n1934), .C(n2014), .Y(n2612) );
  NAND2X1 U1603 ( .A(\mem<28><12> ), .B(n1257), .Y(n2015) );
  OAI21X1 U1604 ( .A(n1256), .B(n1936), .C(n2015), .Y(n2611) );
  NAND2X1 U1605 ( .A(\mem<28><13> ), .B(n1257), .Y(n2016) );
  OAI21X1 U1606 ( .A(n1256), .B(n1938), .C(n2016), .Y(n2610) );
  NAND2X1 U1607 ( .A(\mem<28><14> ), .B(n1257), .Y(n2017) );
  OAI21X1 U1608 ( .A(n1256), .B(n1940), .C(n2017), .Y(n2609) );
  NAND2X1 U1609 ( .A(\mem<28><15> ), .B(n1257), .Y(n2018) );
  OAI21X1 U1610 ( .A(n1256), .B(n1942), .C(n2018), .Y(n2608) );
  NAND3X1 U1611 ( .A(n1945), .B(n1947), .C(n1949), .Y(n2019) );
  NAND2X1 U1612 ( .A(\mem<27><0> ), .B(n1262), .Y(n2020) );
  OAI21X1 U1613 ( .A(n1260), .B(n1912), .C(n2020), .Y(n2607) );
  NAND2X1 U1614 ( .A(\mem<27><1> ), .B(n1262), .Y(n2021) );
  OAI21X1 U1615 ( .A(n1260), .B(n1914), .C(n2021), .Y(n2606) );
  NAND2X1 U1616 ( .A(\mem<27><2> ), .B(n1262), .Y(n2022) );
  OAI21X1 U1617 ( .A(n1260), .B(n1916), .C(n2022), .Y(n2605) );
  NAND2X1 U1618 ( .A(\mem<27><3> ), .B(n1262), .Y(n2023) );
  OAI21X1 U1619 ( .A(n1260), .B(n1918), .C(n2023), .Y(n2604) );
  NAND2X1 U1620 ( .A(\mem<27><4> ), .B(n1262), .Y(n2024) );
  OAI21X1 U1621 ( .A(n1260), .B(n1920), .C(n2024), .Y(n2603) );
  NAND2X1 U1622 ( .A(\mem<27><5> ), .B(n1262), .Y(n2025) );
  OAI21X1 U1623 ( .A(n1260), .B(n1922), .C(n2025), .Y(n2602) );
  NAND2X1 U1624 ( .A(\mem<27><6> ), .B(n1262), .Y(n2026) );
  OAI21X1 U1625 ( .A(n1260), .B(n1924), .C(n2026), .Y(n2601) );
  NAND2X1 U1626 ( .A(\mem<27><7> ), .B(n1262), .Y(n2027) );
  OAI21X1 U1627 ( .A(n1260), .B(n1926), .C(n2027), .Y(n2600) );
  NAND2X1 U1628 ( .A(\mem<27><8> ), .B(n1261), .Y(n2028) );
  OAI21X1 U1629 ( .A(n1260), .B(n1929), .C(n2028), .Y(n2599) );
  NAND2X1 U1630 ( .A(\mem<27><9> ), .B(n1261), .Y(n2029) );
  OAI21X1 U1631 ( .A(n1260), .B(n1931), .C(n2029), .Y(n2598) );
  NAND2X1 U1632 ( .A(\mem<27><10> ), .B(n1261), .Y(n2030) );
  OAI21X1 U1633 ( .A(n1260), .B(n1933), .C(n2030), .Y(n2597) );
  NAND2X1 U1634 ( .A(\mem<27><11> ), .B(n1261), .Y(n2031) );
  OAI21X1 U1635 ( .A(n1260), .B(n1935), .C(n2031), .Y(n2596) );
  NAND2X1 U1636 ( .A(\mem<27><12> ), .B(n1261), .Y(n2032) );
  OAI21X1 U1637 ( .A(n1260), .B(n1937), .C(n2032), .Y(n2595) );
  NAND2X1 U1638 ( .A(\mem<27><13> ), .B(n1261), .Y(n2033) );
  OAI21X1 U1639 ( .A(n1260), .B(n1939), .C(n2033), .Y(n2594) );
  NAND2X1 U1640 ( .A(\mem<27><14> ), .B(n1261), .Y(n2034) );
  OAI21X1 U1641 ( .A(n1260), .B(n1941), .C(n2034), .Y(n2593) );
  NAND2X1 U1642 ( .A(\mem<27><15> ), .B(n1261), .Y(n2035) );
  OAI21X1 U1643 ( .A(n1260), .B(n1943), .C(n2035), .Y(n2592) );
  NAND3X1 U1644 ( .A(n1949), .B(n1947), .C(n1946), .Y(n2036) );
  NAND2X1 U1645 ( .A(\mem<26><0> ), .B(n1266), .Y(n2037) );
  OAI21X1 U1646 ( .A(n1264), .B(n1912), .C(n2037), .Y(n2591) );
  NAND2X1 U1647 ( .A(\mem<26><1> ), .B(n1266), .Y(n2038) );
  OAI21X1 U1648 ( .A(n1264), .B(n1915), .C(n2038), .Y(n2590) );
  NAND2X1 U1649 ( .A(\mem<26><2> ), .B(n1266), .Y(n2039) );
  OAI21X1 U1650 ( .A(n1264), .B(n1917), .C(n2039), .Y(n2589) );
  NAND2X1 U1651 ( .A(\mem<26><3> ), .B(n1266), .Y(n2040) );
  OAI21X1 U1652 ( .A(n1264), .B(n1919), .C(n2040), .Y(n2588) );
  NAND2X1 U1653 ( .A(\mem<26><4> ), .B(n1266), .Y(n2041) );
  OAI21X1 U1654 ( .A(n1264), .B(n1921), .C(n2041), .Y(n2587) );
  NAND2X1 U1655 ( .A(\mem<26><5> ), .B(n1266), .Y(n2042) );
  OAI21X1 U1656 ( .A(n1264), .B(n1923), .C(n2042), .Y(n2586) );
  NAND2X1 U1657 ( .A(\mem<26><6> ), .B(n1266), .Y(n2043) );
  OAI21X1 U1658 ( .A(n1264), .B(n1925), .C(n2043), .Y(n2585) );
  NAND2X1 U1659 ( .A(\mem<26><7> ), .B(n1266), .Y(n2044) );
  OAI21X1 U1660 ( .A(n1264), .B(n1927), .C(n2044), .Y(n2584) );
  NAND2X1 U1661 ( .A(\mem<26><8> ), .B(n1265), .Y(n2045) );
  OAI21X1 U1662 ( .A(n1264), .B(n1928), .C(n2045), .Y(n2583) );
  NAND2X1 U1663 ( .A(\mem<26><9> ), .B(n1265), .Y(n2046) );
  OAI21X1 U1664 ( .A(n1264), .B(n1930), .C(n2046), .Y(n2582) );
  NAND2X1 U1665 ( .A(\mem<26><10> ), .B(n1265), .Y(n2047) );
  OAI21X1 U1666 ( .A(n1264), .B(n1932), .C(n2047), .Y(n2581) );
  NAND2X1 U1667 ( .A(\mem<26><11> ), .B(n1265), .Y(n2048) );
  OAI21X1 U1668 ( .A(n1264), .B(n1934), .C(n2048), .Y(n2580) );
  NAND2X1 U1669 ( .A(\mem<26><12> ), .B(n1265), .Y(n2049) );
  OAI21X1 U1670 ( .A(n1264), .B(n1936), .C(n2049), .Y(n2579) );
  NAND2X1 U1671 ( .A(\mem<26><13> ), .B(n1265), .Y(n2050) );
  OAI21X1 U1672 ( .A(n1264), .B(n1938), .C(n2050), .Y(n2578) );
  NAND2X1 U1673 ( .A(\mem<26><14> ), .B(n1265), .Y(n2051) );
  OAI21X1 U1674 ( .A(n1264), .B(n1940), .C(n2051), .Y(n2577) );
  NAND2X1 U1675 ( .A(\mem<26><15> ), .B(n1265), .Y(n2052) );
  OAI21X1 U1676 ( .A(n1264), .B(n1942), .C(n2052), .Y(n2576) );
  NAND3X1 U1677 ( .A(n1945), .B(n1949), .C(n1948), .Y(n2053) );
  NAND2X1 U1678 ( .A(\mem<25><0> ), .B(n1270), .Y(n2054) );
  OAI21X1 U1679 ( .A(n1268), .B(n1912), .C(n2054), .Y(n2575) );
  NAND2X1 U1680 ( .A(\mem<25><1> ), .B(n1270), .Y(n2055) );
  OAI21X1 U1681 ( .A(n1268), .B(n1914), .C(n2055), .Y(n2574) );
  NAND2X1 U1682 ( .A(\mem<25><2> ), .B(n1270), .Y(n2056) );
  OAI21X1 U1683 ( .A(n1268), .B(n1916), .C(n2056), .Y(n2573) );
  NAND2X1 U1684 ( .A(\mem<25><3> ), .B(n1270), .Y(n2057) );
  OAI21X1 U1685 ( .A(n1268), .B(n1918), .C(n2057), .Y(n2572) );
  NAND2X1 U1686 ( .A(\mem<25><4> ), .B(n1270), .Y(n2058) );
  OAI21X1 U1687 ( .A(n1268), .B(n1920), .C(n2058), .Y(n2571) );
  NAND2X1 U1688 ( .A(\mem<25><5> ), .B(n1270), .Y(n2059) );
  OAI21X1 U1689 ( .A(n1268), .B(n1922), .C(n2059), .Y(n2570) );
  NAND2X1 U1690 ( .A(\mem<25><6> ), .B(n1270), .Y(n2060) );
  OAI21X1 U1691 ( .A(n1268), .B(n1924), .C(n2060), .Y(n2569) );
  NAND2X1 U1692 ( .A(\mem<25><7> ), .B(n1270), .Y(n2061) );
  OAI21X1 U1693 ( .A(n1268), .B(n1926), .C(n2061), .Y(n2568) );
  NAND2X1 U1694 ( .A(\mem<25><8> ), .B(n1269), .Y(n2062) );
  OAI21X1 U1695 ( .A(n1268), .B(n1929), .C(n2062), .Y(n2567) );
  NAND2X1 U1696 ( .A(\mem<25><9> ), .B(n1269), .Y(n2063) );
  OAI21X1 U1697 ( .A(n1268), .B(n1931), .C(n2063), .Y(n2566) );
  NAND2X1 U1698 ( .A(\mem<25><10> ), .B(n1269), .Y(n2064) );
  OAI21X1 U1699 ( .A(n1268), .B(n1933), .C(n2064), .Y(n2565) );
  NAND2X1 U1700 ( .A(\mem<25><11> ), .B(n1269), .Y(n2065) );
  OAI21X1 U1701 ( .A(n1268), .B(n1935), .C(n2065), .Y(n2564) );
  NAND2X1 U1702 ( .A(\mem<25><12> ), .B(n1269), .Y(n2066) );
  OAI21X1 U1703 ( .A(n1268), .B(n1937), .C(n2066), .Y(n2563) );
  NAND2X1 U1704 ( .A(\mem<25><13> ), .B(n1269), .Y(n2067) );
  OAI21X1 U1705 ( .A(n1268), .B(n1939), .C(n2067), .Y(n2562) );
  NAND2X1 U1706 ( .A(\mem<25><14> ), .B(n1269), .Y(n2068) );
  OAI21X1 U1707 ( .A(n1268), .B(n1941), .C(n2068), .Y(n2561) );
  NAND2X1 U1708 ( .A(\mem<25><15> ), .B(n1269), .Y(n2069) );
  OAI21X1 U1709 ( .A(n1268), .B(n1943), .C(n2069), .Y(n2560) );
  NOR3X1 U1710 ( .A(n1945), .B(n1947), .C(n1827), .Y(n2159) );
  NAND2X1 U1711 ( .A(\mem<24><0> ), .B(n1272), .Y(n2070) );
  OAI21X1 U1712 ( .A(n1863), .B(n1912), .C(n2070), .Y(n2559) );
  NAND2X1 U1713 ( .A(\mem<24><1> ), .B(n1272), .Y(n2071) );
  OAI21X1 U1714 ( .A(n1863), .B(n1914), .C(n2071), .Y(n2558) );
  NAND2X1 U1715 ( .A(\mem<24><2> ), .B(n1272), .Y(n2072) );
  OAI21X1 U1716 ( .A(n1863), .B(n1916), .C(n2072), .Y(n2557) );
  NAND2X1 U1717 ( .A(\mem<24><3> ), .B(n1272), .Y(n2073) );
  OAI21X1 U1718 ( .A(n1863), .B(n1918), .C(n2073), .Y(n2556) );
  NAND2X1 U1719 ( .A(\mem<24><4> ), .B(n1272), .Y(n2074) );
  OAI21X1 U1720 ( .A(n1863), .B(n1920), .C(n2074), .Y(n2555) );
  NAND2X1 U1721 ( .A(\mem<24><5> ), .B(n1272), .Y(n2075) );
  OAI21X1 U1722 ( .A(n1863), .B(n1922), .C(n2075), .Y(n2554) );
  NAND2X1 U1723 ( .A(\mem<24><6> ), .B(n1272), .Y(n2076) );
  OAI21X1 U1724 ( .A(n1863), .B(n1924), .C(n2076), .Y(n2553) );
  NAND2X1 U1725 ( .A(\mem<24><7> ), .B(n1272), .Y(n2077) );
  OAI21X1 U1726 ( .A(n1863), .B(n1926), .C(n2077), .Y(n2552) );
  NAND2X1 U1727 ( .A(\mem<24><8> ), .B(n1271), .Y(n2078) );
  OAI21X1 U1728 ( .A(n1863), .B(n1928), .C(n2078), .Y(n2551) );
  NAND2X1 U1729 ( .A(\mem<24><9> ), .B(n1271), .Y(n2079) );
  OAI21X1 U1730 ( .A(n1863), .B(n1930), .C(n2079), .Y(n2550) );
  NAND2X1 U1731 ( .A(\mem<24><10> ), .B(n1271), .Y(n2080) );
  OAI21X1 U1732 ( .A(n1863), .B(n1932), .C(n2080), .Y(n2549) );
  NAND2X1 U1733 ( .A(\mem<24><11> ), .B(n1271), .Y(n2081) );
  OAI21X1 U1734 ( .A(n1863), .B(n1934), .C(n2081), .Y(n2548) );
  NAND2X1 U1735 ( .A(\mem<24><12> ), .B(n1271), .Y(n2082) );
  OAI21X1 U1736 ( .A(n1863), .B(n1936), .C(n2082), .Y(n2547) );
  NAND2X1 U1737 ( .A(\mem<24><13> ), .B(n1271), .Y(n2083) );
  OAI21X1 U1738 ( .A(n1863), .B(n1938), .C(n2083), .Y(n2546) );
  NAND2X1 U1739 ( .A(\mem<24><14> ), .B(n1271), .Y(n2084) );
  OAI21X1 U1740 ( .A(n1863), .B(n1940), .C(n2084), .Y(n2545) );
  NAND2X1 U1741 ( .A(\mem<24><15> ), .B(n1271), .Y(n2085) );
  OAI21X1 U1742 ( .A(n1863), .B(n1942), .C(n2085), .Y(n2544) );
  NAND2X1 U1743 ( .A(\mem<23><0> ), .B(n1276), .Y(n2086) );
  OAI21X1 U1744 ( .A(n1274), .B(n1912), .C(n2086), .Y(n2543) );
  NAND2X1 U1745 ( .A(\mem<23><1> ), .B(n1276), .Y(n2087) );
  OAI21X1 U1746 ( .A(n1274), .B(n1915), .C(n2087), .Y(n2542) );
  NAND2X1 U1747 ( .A(\mem<23><2> ), .B(n1276), .Y(n2088) );
  OAI21X1 U1748 ( .A(n1274), .B(n1917), .C(n2088), .Y(n2541) );
  NAND2X1 U1749 ( .A(\mem<23><3> ), .B(n1276), .Y(n2089) );
  OAI21X1 U1750 ( .A(n1274), .B(n1919), .C(n2089), .Y(n2540) );
  NAND2X1 U1751 ( .A(\mem<23><4> ), .B(n1276), .Y(n2090) );
  OAI21X1 U1752 ( .A(n1274), .B(n1921), .C(n2090), .Y(n2539) );
  NAND2X1 U1753 ( .A(\mem<23><5> ), .B(n1276), .Y(n2091) );
  OAI21X1 U1754 ( .A(n1274), .B(n1923), .C(n2091), .Y(n2538) );
  NAND2X1 U1755 ( .A(\mem<23><6> ), .B(n1276), .Y(n2092) );
  OAI21X1 U1756 ( .A(n1274), .B(n1925), .C(n2092), .Y(n2537) );
  NAND2X1 U1757 ( .A(\mem<23><7> ), .B(n1276), .Y(n2093) );
  OAI21X1 U1758 ( .A(n1274), .B(n1927), .C(n2093), .Y(n2536) );
  NAND2X1 U1759 ( .A(\mem<23><8> ), .B(n1275), .Y(n2094) );
  OAI21X1 U1760 ( .A(n1274), .B(n1929), .C(n2094), .Y(n2535) );
  NAND2X1 U1761 ( .A(\mem<23><9> ), .B(n1275), .Y(n2095) );
  OAI21X1 U1762 ( .A(n1274), .B(n1931), .C(n2095), .Y(n2534) );
  NAND2X1 U1763 ( .A(\mem<23><10> ), .B(n1275), .Y(n2096) );
  OAI21X1 U1764 ( .A(n1274), .B(n1933), .C(n2096), .Y(n2533) );
  NAND2X1 U1765 ( .A(\mem<23><11> ), .B(n1275), .Y(n2097) );
  OAI21X1 U1766 ( .A(n1274), .B(n1935), .C(n2097), .Y(n2532) );
  NAND2X1 U1767 ( .A(\mem<23><12> ), .B(n1275), .Y(n2098) );
  OAI21X1 U1768 ( .A(n1274), .B(n1937), .C(n2098), .Y(n2531) );
  NAND2X1 U1769 ( .A(\mem<23><13> ), .B(n1275), .Y(n2099) );
  OAI21X1 U1770 ( .A(n1274), .B(n1939), .C(n2099), .Y(n2530) );
  NAND2X1 U1771 ( .A(\mem<23><14> ), .B(n1275), .Y(n2100) );
  OAI21X1 U1772 ( .A(n1274), .B(n1941), .C(n2100), .Y(n2529) );
  NAND2X1 U1773 ( .A(\mem<23><15> ), .B(n1275), .Y(n2101) );
  OAI21X1 U1774 ( .A(n1274), .B(n1943), .C(n2101), .Y(n2528) );
  NAND2X1 U1775 ( .A(\mem<22><0> ), .B(n1280), .Y(n2102) );
  OAI21X1 U1776 ( .A(n1278), .B(n1912), .C(n2102), .Y(n2527) );
  NAND2X1 U1777 ( .A(\mem<22><1> ), .B(n1280), .Y(n2103) );
  OAI21X1 U1778 ( .A(n1278), .B(n1915), .C(n2103), .Y(n2526) );
  NAND2X1 U1779 ( .A(\mem<22><2> ), .B(n1280), .Y(n2104) );
  OAI21X1 U1780 ( .A(n1278), .B(n1917), .C(n2104), .Y(n2525) );
  NAND2X1 U1781 ( .A(\mem<22><3> ), .B(n1280), .Y(n2105) );
  OAI21X1 U1782 ( .A(n1278), .B(n1919), .C(n2105), .Y(n2524) );
  NAND2X1 U1783 ( .A(\mem<22><4> ), .B(n1280), .Y(n2106) );
  OAI21X1 U1784 ( .A(n1278), .B(n1921), .C(n2106), .Y(n2523) );
  NAND2X1 U1785 ( .A(\mem<22><5> ), .B(n1280), .Y(n2107) );
  OAI21X1 U1786 ( .A(n1278), .B(n1923), .C(n2107), .Y(n2522) );
  NAND2X1 U1787 ( .A(\mem<22><6> ), .B(n1280), .Y(n2108) );
  OAI21X1 U1788 ( .A(n1278), .B(n1925), .C(n2108), .Y(n2521) );
  NAND2X1 U1789 ( .A(\mem<22><7> ), .B(n1280), .Y(n2109) );
  OAI21X1 U1790 ( .A(n1278), .B(n1927), .C(n2109), .Y(n2520) );
  NAND2X1 U1791 ( .A(\mem<22><8> ), .B(n1279), .Y(n2110) );
  OAI21X1 U1792 ( .A(n1278), .B(n1929), .C(n2110), .Y(n2519) );
  NAND2X1 U1793 ( .A(\mem<22><9> ), .B(n1279), .Y(n2111) );
  OAI21X1 U1794 ( .A(n1278), .B(n1931), .C(n2111), .Y(n2518) );
  NAND2X1 U1795 ( .A(\mem<22><10> ), .B(n1279), .Y(n2112) );
  OAI21X1 U1796 ( .A(n1278), .B(n1933), .C(n2112), .Y(n2517) );
  NAND2X1 U1797 ( .A(\mem<22><11> ), .B(n1279), .Y(n2113) );
  OAI21X1 U1798 ( .A(n1278), .B(n1935), .C(n2113), .Y(n2516) );
  NAND2X1 U1799 ( .A(\mem<22><12> ), .B(n1279), .Y(n2114) );
  OAI21X1 U1800 ( .A(n1278), .B(n1937), .C(n2114), .Y(n2515) );
  NAND2X1 U1801 ( .A(\mem<22><13> ), .B(n1279), .Y(n2115) );
  OAI21X1 U1802 ( .A(n1278), .B(n1939), .C(n2115), .Y(n2514) );
  NAND2X1 U1803 ( .A(\mem<22><14> ), .B(n1279), .Y(n2116) );
  OAI21X1 U1804 ( .A(n1278), .B(n1941), .C(n2116), .Y(n2513) );
  NAND2X1 U1805 ( .A(\mem<22><15> ), .B(n1279), .Y(n2117) );
  OAI21X1 U1806 ( .A(n1278), .B(n1943), .C(n2117), .Y(n2512) );
  NAND2X1 U1807 ( .A(\mem<21><0> ), .B(n1284), .Y(n2118) );
  OAI21X1 U1808 ( .A(n1282), .B(n1912), .C(n2118), .Y(n2511) );
  NAND2X1 U1809 ( .A(\mem<21><1> ), .B(n1284), .Y(n2119) );
  OAI21X1 U1810 ( .A(n1282), .B(n1915), .C(n2119), .Y(n2510) );
  NAND2X1 U1811 ( .A(\mem<21><2> ), .B(n1284), .Y(n2120) );
  OAI21X1 U1812 ( .A(n1282), .B(n1917), .C(n2120), .Y(n2509) );
  NAND2X1 U1813 ( .A(\mem<21><3> ), .B(n1284), .Y(n2121) );
  OAI21X1 U1814 ( .A(n1282), .B(n1919), .C(n2121), .Y(n2508) );
  NAND2X1 U1815 ( .A(\mem<21><4> ), .B(n1284), .Y(n2122) );
  OAI21X1 U1816 ( .A(n1282), .B(n1921), .C(n2122), .Y(n2507) );
  NAND2X1 U1817 ( .A(\mem<21><5> ), .B(n1284), .Y(n2123) );
  OAI21X1 U1818 ( .A(n1282), .B(n1923), .C(n2123), .Y(n2506) );
  NAND2X1 U1819 ( .A(\mem<21><6> ), .B(n1284), .Y(n2124) );
  OAI21X1 U1820 ( .A(n1282), .B(n1925), .C(n2124), .Y(n2505) );
  NAND2X1 U1821 ( .A(\mem<21><7> ), .B(n1284), .Y(n2125) );
  OAI21X1 U1822 ( .A(n1282), .B(n1927), .C(n2125), .Y(n2504) );
  NAND2X1 U1823 ( .A(\mem<21><8> ), .B(n1283), .Y(n2126) );
  OAI21X1 U1824 ( .A(n1282), .B(n1929), .C(n2126), .Y(n2503) );
  NAND2X1 U1825 ( .A(\mem<21><9> ), .B(n1283), .Y(n2127) );
  OAI21X1 U1826 ( .A(n1282), .B(n1931), .C(n2127), .Y(n2502) );
  NAND2X1 U1827 ( .A(\mem<21><10> ), .B(n1283), .Y(n2128) );
  OAI21X1 U1828 ( .A(n1282), .B(n1933), .C(n2128), .Y(n2501) );
  NAND2X1 U1829 ( .A(\mem<21><11> ), .B(n1283), .Y(n2129) );
  OAI21X1 U1830 ( .A(n1282), .B(n1935), .C(n2129), .Y(n2500) );
  NAND2X1 U1831 ( .A(\mem<21><12> ), .B(n1283), .Y(n2130) );
  OAI21X1 U1832 ( .A(n1282), .B(n1937), .C(n2130), .Y(n2499) );
  NAND2X1 U1833 ( .A(\mem<21><13> ), .B(n1283), .Y(n2131) );
  OAI21X1 U1834 ( .A(n1282), .B(n1939), .C(n2131), .Y(n2498) );
  NAND2X1 U1835 ( .A(\mem<21><14> ), .B(n1283), .Y(n2132) );
  OAI21X1 U1836 ( .A(n1282), .B(n1941), .C(n2132), .Y(n2497) );
  NAND2X1 U1837 ( .A(\mem<21><15> ), .B(n1283), .Y(n2133) );
  OAI21X1 U1838 ( .A(n1282), .B(n1943), .C(n2133), .Y(n2496) );
  NAND2X1 U1839 ( .A(\mem<20><0> ), .B(n1288), .Y(n2134) );
  OAI21X1 U1840 ( .A(n1286), .B(n1912), .C(n2134), .Y(n2495) );
  NAND2X1 U1841 ( .A(\mem<20><1> ), .B(n1288), .Y(n2135) );
  OAI21X1 U1842 ( .A(n1286), .B(n1915), .C(n2135), .Y(n2494) );
  NAND2X1 U1843 ( .A(\mem<20><2> ), .B(n1288), .Y(n2136) );
  OAI21X1 U1844 ( .A(n1286), .B(n1917), .C(n2136), .Y(n2493) );
  NAND2X1 U1845 ( .A(\mem<20><3> ), .B(n1288), .Y(n2137) );
  OAI21X1 U1846 ( .A(n1286), .B(n1919), .C(n2137), .Y(n2492) );
  NAND2X1 U1847 ( .A(\mem<20><4> ), .B(n1288), .Y(n2138) );
  OAI21X1 U1848 ( .A(n1286), .B(n1921), .C(n2138), .Y(n2491) );
  NAND2X1 U1849 ( .A(\mem<20><5> ), .B(n1288), .Y(n2139) );
  OAI21X1 U1850 ( .A(n1286), .B(n1923), .C(n2139), .Y(n2490) );
  NAND2X1 U1851 ( .A(\mem<20><6> ), .B(n1288), .Y(n2140) );
  OAI21X1 U1852 ( .A(n1286), .B(n1925), .C(n2140), .Y(n2489) );
  NAND2X1 U1853 ( .A(\mem<20><7> ), .B(n1288), .Y(n2141) );
  OAI21X1 U1854 ( .A(n1286), .B(n1927), .C(n2141), .Y(n2488) );
  NAND2X1 U1855 ( .A(\mem<20><8> ), .B(n1287), .Y(n2142) );
  OAI21X1 U1856 ( .A(n1286), .B(n1929), .C(n2142), .Y(n2487) );
  NAND2X1 U1857 ( .A(\mem<20><9> ), .B(n1287), .Y(n2143) );
  OAI21X1 U1858 ( .A(n1286), .B(n1931), .C(n2143), .Y(n2486) );
  NAND2X1 U1859 ( .A(\mem<20><10> ), .B(n1287), .Y(n2144) );
  OAI21X1 U1860 ( .A(n1286), .B(n1933), .C(n2144), .Y(n2485) );
  NAND2X1 U1861 ( .A(\mem<20><11> ), .B(n1287), .Y(n2145) );
  OAI21X1 U1862 ( .A(n1286), .B(n1935), .C(n2145), .Y(n2484) );
  NAND2X1 U1863 ( .A(\mem<20><12> ), .B(n1287), .Y(n2146) );
  OAI21X1 U1864 ( .A(n1286), .B(n1937), .C(n2146), .Y(n2483) );
  NAND2X1 U1865 ( .A(\mem<20><13> ), .B(n1287), .Y(n2147) );
  OAI21X1 U1866 ( .A(n1286), .B(n1939), .C(n2147), .Y(n2482) );
  NAND2X1 U1867 ( .A(\mem<20><14> ), .B(n1287), .Y(n2148) );
  OAI21X1 U1868 ( .A(n1286), .B(n1941), .C(n2148), .Y(n2481) );
  NAND2X1 U1869 ( .A(\mem<20><15> ), .B(n1287), .Y(n2149) );
  OAI21X1 U1870 ( .A(n1286), .B(n1943), .C(n2149), .Y(n2480) );
  OAI21X1 U1871 ( .A(n1290), .B(n1913), .C(n74), .Y(n2479) );
  OAI21X1 U1872 ( .A(n1290), .B(n1915), .C(n76), .Y(n2478) );
  OAI21X1 U1873 ( .A(n1290), .B(n1917), .C(n78), .Y(n2477) );
  OAI21X1 U1874 ( .A(n1290), .B(n1919), .C(n80), .Y(n2476) );
  OAI21X1 U1875 ( .A(n1290), .B(n1921), .C(n82), .Y(n2475) );
  OAI21X1 U1876 ( .A(n1290), .B(n1923), .C(n84), .Y(n2474) );
  OAI21X1 U1877 ( .A(n1290), .B(n1925), .C(n86), .Y(n2473) );
  OAI21X1 U1878 ( .A(n1290), .B(n1927), .C(n88), .Y(n2472) );
  OAI21X1 U1879 ( .A(n1290), .B(n1929), .C(n90), .Y(n2471) );
  OAI21X1 U1880 ( .A(n1290), .B(n1931), .C(n92), .Y(n2470) );
  OAI21X1 U1881 ( .A(n1290), .B(n1933), .C(n94), .Y(n2469) );
  OAI21X1 U1882 ( .A(n1290), .B(n1935), .C(n96), .Y(n2468) );
  OAI21X1 U1883 ( .A(n1290), .B(n1937), .C(n98), .Y(n2467) );
  OAI21X1 U1884 ( .A(n1290), .B(n1939), .C(n100), .Y(n2466) );
  OAI21X1 U1885 ( .A(n1290), .B(n1941), .C(n102), .Y(n2465) );
  OAI21X1 U1886 ( .A(n1290), .B(n1943), .C(n104), .Y(n2464) );
  OAI21X1 U1887 ( .A(n1292), .B(n1913), .C(n106), .Y(n2463) );
  OAI21X1 U1888 ( .A(n1292), .B(n1915), .C(n108), .Y(n2462) );
  OAI21X1 U1889 ( .A(n1292), .B(n1917), .C(n110), .Y(n2461) );
  OAI21X1 U1890 ( .A(n1292), .B(n1919), .C(n112), .Y(n2460) );
  OAI21X1 U1891 ( .A(n1292), .B(n1921), .C(n114), .Y(n2459) );
  OAI21X1 U1892 ( .A(n1292), .B(n1923), .C(n116), .Y(n2458) );
  OAI21X1 U1893 ( .A(n1292), .B(n1925), .C(n118), .Y(n2457) );
  OAI21X1 U1894 ( .A(n1292), .B(n1927), .C(n120), .Y(n2456) );
  OAI21X1 U1895 ( .A(n1292), .B(n1929), .C(n122), .Y(n2455) );
  OAI21X1 U1896 ( .A(n1292), .B(n1931), .C(n124), .Y(n2454) );
  OAI21X1 U1897 ( .A(n1292), .B(n1933), .C(n126), .Y(n2453) );
  OAI21X1 U1898 ( .A(n1292), .B(n1935), .C(n128), .Y(n2452) );
  OAI21X1 U1899 ( .A(n1292), .B(n1937), .C(n130), .Y(n2451) );
  OAI21X1 U1900 ( .A(n1292), .B(n1939), .C(n132), .Y(n2450) );
  OAI21X1 U1901 ( .A(n1292), .B(n1941), .C(n134), .Y(n2449) );
  OAI21X1 U1902 ( .A(n1292), .B(n1943), .C(n136), .Y(n2448) );
  OAI21X1 U1903 ( .A(n1294), .B(n1913), .C(n138), .Y(n2447) );
  OAI21X1 U1904 ( .A(n1294), .B(n1915), .C(n140), .Y(n2446) );
  OAI21X1 U1905 ( .A(n1294), .B(n1917), .C(n142), .Y(n2445) );
  OAI21X1 U1906 ( .A(n1294), .B(n1919), .C(n144), .Y(n2444) );
  OAI21X1 U1907 ( .A(n1294), .B(n1921), .C(n146), .Y(n2443) );
  OAI21X1 U1908 ( .A(n1294), .B(n1923), .C(n148), .Y(n2442) );
  OAI21X1 U1909 ( .A(n1294), .B(n1925), .C(n150), .Y(n2441) );
  OAI21X1 U1910 ( .A(n1294), .B(n1927), .C(n152), .Y(n2440) );
  OAI21X1 U1911 ( .A(n1294), .B(n1929), .C(n154), .Y(n2439) );
  OAI21X1 U1912 ( .A(n1294), .B(n1931), .C(n156), .Y(n2438) );
  OAI21X1 U1913 ( .A(n1294), .B(n1933), .C(n158), .Y(n2437) );
  OAI21X1 U1914 ( .A(n1294), .B(n1935), .C(n160), .Y(n2436) );
  OAI21X1 U1915 ( .A(n1294), .B(n1937), .C(n162), .Y(n2435) );
  OAI21X1 U1916 ( .A(n1294), .B(n1939), .C(n164), .Y(n2434) );
  OAI21X1 U1917 ( .A(n1294), .B(n1941), .C(n166), .Y(n2433) );
  OAI21X1 U1918 ( .A(n1294), .B(n1943), .C(n168), .Y(n2432) );
  OAI21X1 U1919 ( .A(n1870), .B(n1913), .C(n170), .Y(n2431) );
  OAI21X1 U1920 ( .A(n1870), .B(n1915), .C(n172), .Y(n2430) );
  OAI21X1 U1921 ( .A(n1870), .B(n1917), .C(n174), .Y(n2429) );
  OAI21X1 U1922 ( .A(n1870), .B(n1919), .C(n176), .Y(n2428) );
  OAI21X1 U1923 ( .A(n1870), .B(n1921), .C(n178), .Y(n2427) );
  OAI21X1 U1924 ( .A(n1870), .B(n1923), .C(n180), .Y(n2426) );
  OAI21X1 U1925 ( .A(n1870), .B(n1925), .C(n182), .Y(n2425) );
  OAI21X1 U1926 ( .A(n1870), .B(n1927), .C(n184), .Y(n2424) );
  OAI21X1 U1927 ( .A(n1870), .B(n1929), .C(n186), .Y(n2423) );
  OAI21X1 U1928 ( .A(n1870), .B(n1931), .C(n188), .Y(n2422) );
  OAI21X1 U1929 ( .A(n1870), .B(n1933), .C(n190), .Y(n2421) );
  OAI21X1 U1930 ( .A(n1870), .B(n1935), .C(n192), .Y(n2420) );
  OAI21X1 U1931 ( .A(n1870), .B(n1937), .C(n194), .Y(n2419) );
  OAI21X1 U1932 ( .A(n1870), .B(n1939), .C(n196), .Y(n2418) );
  OAI21X1 U1933 ( .A(n1870), .B(n1941), .C(n198), .Y(n2417) );
  OAI21X1 U1934 ( .A(n1870), .B(n1943), .C(n200), .Y(n2416) );
  NAND3X1 U1935 ( .A(n1950), .B(n2672), .C(n1952), .Y(n2150) );
  OAI21X1 U1936 ( .A(n1296), .B(n1913), .C(n202), .Y(n2415) );
  OAI21X1 U1937 ( .A(n1296), .B(n1915), .C(n204), .Y(n2414) );
  OAI21X1 U1938 ( .A(n1296), .B(n1917), .C(n206), .Y(n2413) );
  OAI21X1 U1939 ( .A(n1296), .B(n1919), .C(n208), .Y(n2412) );
  OAI21X1 U1940 ( .A(n1296), .B(n1921), .C(n210), .Y(n2411) );
  OAI21X1 U1941 ( .A(n1296), .B(n1923), .C(n212), .Y(n2410) );
  OAI21X1 U1942 ( .A(n1296), .B(n1925), .C(n215), .Y(n2409) );
  OAI21X1 U1943 ( .A(n1296), .B(n1927), .C(n217), .Y(n2408) );
  OAI21X1 U1944 ( .A(n1296), .B(n1929), .C(n219), .Y(n2407) );
  OAI21X1 U1945 ( .A(n1296), .B(n1931), .C(n221), .Y(n2406) );
  OAI21X1 U1946 ( .A(n1296), .B(n1933), .C(n223), .Y(n2405) );
  OAI21X1 U1947 ( .A(n1296), .B(n1935), .C(n225), .Y(n2404) );
  OAI21X1 U1948 ( .A(n1296), .B(n1937), .C(n227), .Y(n2403) );
  OAI21X1 U1949 ( .A(n1296), .B(n1939), .C(n229), .Y(n2402) );
  OAI21X1 U1950 ( .A(n1296), .B(n1941), .C(n231), .Y(n2401) );
  OAI21X1 U1951 ( .A(n1296), .B(n1943), .C(n233), .Y(n2400) );
  OAI21X1 U1952 ( .A(n1298), .B(n1913), .C(n235), .Y(n2399) );
  OAI21X1 U1953 ( .A(n1298), .B(n1915), .C(n237), .Y(n2398) );
  OAI21X1 U1954 ( .A(n1298), .B(n1917), .C(n239), .Y(n2397) );
  OAI21X1 U1955 ( .A(n1298), .B(n1919), .C(n241), .Y(n2396) );
  OAI21X1 U1956 ( .A(n1298), .B(n1921), .C(n243), .Y(n2395) );
  OAI21X1 U1957 ( .A(n1298), .B(n1923), .C(n245), .Y(n2394) );
  OAI21X1 U1958 ( .A(n1298), .B(n1925), .C(n247), .Y(n2393) );
  OAI21X1 U1959 ( .A(n1298), .B(n1927), .C(n249), .Y(n2392) );
  OAI21X1 U1960 ( .A(n1298), .B(n1929), .C(n251), .Y(n2391) );
  OAI21X1 U1961 ( .A(n1298), .B(n1931), .C(n253), .Y(n2390) );
  OAI21X1 U1962 ( .A(n1298), .B(n1933), .C(n255), .Y(n2389) );
  OAI21X1 U1963 ( .A(n1298), .B(n1935), .C(n257), .Y(n2388) );
  OAI21X1 U1964 ( .A(n1298), .B(n1937), .C(n259), .Y(n2387) );
  OAI21X1 U1965 ( .A(n1298), .B(n1939), .C(n261), .Y(n2386) );
  OAI21X1 U1966 ( .A(n1298), .B(n1941), .C(n263), .Y(n2385) );
  OAI21X1 U1967 ( .A(n1298), .B(n1943), .C(n265), .Y(n2384) );
  OAI21X1 U1968 ( .A(n1300), .B(n1913), .C(n267), .Y(n2383) );
  OAI21X1 U1969 ( .A(n1300), .B(n1915), .C(n269), .Y(n2382) );
  OAI21X1 U1970 ( .A(n1300), .B(n1917), .C(n271), .Y(n2381) );
  OAI21X1 U1971 ( .A(n1300), .B(n1919), .C(n273), .Y(n2380) );
  OAI21X1 U1972 ( .A(n1300), .B(n1921), .C(n275), .Y(n2379) );
  OAI21X1 U1973 ( .A(n1300), .B(n1923), .C(n277), .Y(n2378) );
  OAI21X1 U1974 ( .A(n1300), .B(n1925), .C(n279), .Y(n2377) );
  OAI21X1 U1975 ( .A(n1300), .B(n1927), .C(n281), .Y(n2376) );
  OAI21X1 U1976 ( .A(n1300), .B(n1929), .C(n283), .Y(n2375) );
  OAI21X1 U1977 ( .A(n1300), .B(n1931), .C(n285), .Y(n2374) );
  OAI21X1 U1978 ( .A(n1300), .B(n1933), .C(n287), .Y(n2373) );
  OAI21X1 U1979 ( .A(n1300), .B(n1935), .C(n289), .Y(n2372) );
  OAI21X1 U1980 ( .A(n1300), .B(n1937), .C(n291), .Y(n2371) );
  OAI21X1 U1981 ( .A(n1300), .B(n1939), .C(n293), .Y(n2370) );
  OAI21X1 U1982 ( .A(n1300), .B(n1941), .C(n295), .Y(n2369) );
  OAI21X1 U1983 ( .A(n1300), .B(n1943), .C(n297), .Y(n2368) );
  OAI21X1 U1984 ( .A(n1302), .B(n1913), .C(n299), .Y(n2367) );
  OAI21X1 U1985 ( .A(n1302), .B(n1915), .C(n301), .Y(n2366) );
  OAI21X1 U1986 ( .A(n1302), .B(n1917), .C(n303), .Y(n2365) );
  OAI21X1 U1987 ( .A(n1302), .B(n1919), .C(n305), .Y(n2364) );
  OAI21X1 U1988 ( .A(n1302), .B(n1921), .C(n307), .Y(n2363) );
  OAI21X1 U1989 ( .A(n1302), .B(n1923), .C(n309), .Y(n2362) );
  OAI21X1 U1990 ( .A(n1302), .B(n1925), .C(n311), .Y(n2361) );
  OAI21X1 U1991 ( .A(n1302), .B(n1927), .C(n313), .Y(n2360) );
  OAI21X1 U1992 ( .A(n1302), .B(n1929), .C(n315), .Y(n2359) );
  OAI21X1 U1993 ( .A(n1302), .B(n1931), .C(n317), .Y(n2358) );
  OAI21X1 U1994 ( .A(n1302), .B(n1933), .C(n319), .Y(n2357) );
  OAI21X1 U1995 ( .A(n1302), .B(n1935), .C(n321), .Y(n2356) );
  OAI21X1 U1996 ( .A(n1302), .B(n1937), .C(n323), .Y(n2355) );
  OAI21X1 U1997 ( .A(n1302), .B(n1939), .C(n325), .Y(n2354) );
  OAI21X1 U1998 ( .A(n1302), .B(n1941), .C(n327), .Y(n2353) );
  OAI21X1 U1999 ( .A(n1302), .B(n1943), .C(n329), .Y(n2352) );
  OAI21X1 U2000 ( .A(n1304), .B(n1913), .C(n331), .Y(n2351) );
  OAI21X1 U2001 ( .A(n1304), .B(n1914), .C(n333), .Y(n2350) );
  OAI21X1 U2002 ( .A(n1304), .B(n1916), .C(n335), .Y(n2349) );
  OAI21X1 U2003 ( .A(n1304), .B(n1918), .C(n337), .Y(n2348) );
  OAI21X1 U2004 ( .A(n1304), .B(n1920), .C(n339), .Y(n2347) );
  OAI21X1 U2005 ( .A(n1304), .B(n1922), .C(n341), .Y(n2346) );
  OAI21X1 U2006 ( .A(n1304), .B(n1924), .C(n343), .Y(n2345) );
  OAI21X1 U2007 ( .A(n1304), .B(n1926), .C(n345), .Y(n2344) );
  OAI21X1 U2008 ( .A(n1304), .B(n1928), .C(n347), .Y(n2343) );
  OAI21X1 U2009 ( .A(n1304), .B(n1930), .C(n349), .Y(n2342) );
  OAI21X1 U2010 ( .A(n1304), .B(n1932), .C(n351), .Y(n2341) );
  OAI21X1 U2011 ( .A(n1304), .B(n1934), .C(n353), .Y(n2340) );
  OAI21X1 U2012 ( .A(n1304), .B(n1936), .C(n355), .Y(n2339) );
  OAI21X1 U2013 ( .A(n1304), .B(n1938), .C(n357), .Y(n2338) );
  OAI21X1 U2014 ( .A(n1304), .B(n1940), .C(n359), .Y(n2337) );
  OAI21X1 U2015 ( .A(n1304), .B(n1942), .C(n361), .Y(n2336) );
  OAI21X1 U2016 ( .A(n1306), .B(n1913), .C(n363), .Y(n2335) );
  OAI21X1 U2017 ( .A(n1306), .B(n1914), .C(n365), .Y(n2334) );
  OAI21X1 U2018 ( .A(n1306), .B(n1916), .C(n367), .Y(n2333) );
  OAI21X1 U2019 ( .A(n1306), .B(n1918), .C(n369), .Y(n2332) );
  OAI21X1 U2020 ( .A(n1306), .B(n1920), .C(n371), .Y(n2331) );
  OAI21X1 U2021 ( .A(n1306), .B(n1922), .C(n373), .Y(n2330) );
  OAI21X1 U2022 ( .A(n1306), .B(n1924), .C(n375), .Y(n2329) );
  OAI21X1 U2023 ( .A(n1306), .B(n1926), .C(n377), .Y(n2328) );
  OAI21X1 U2024 ( .A(n1306), .B(n1928), .C(n379), .Y(n2327) );
  OAI21X1 U2025 ( .A(n1306), .B(n1930), .C(n381), .Y(n2326) );
  OAI21X1 U2026 ( .A(n1306), .B(n1932), .C(n383), .Y(n2325) );
  OAI21X1 U2027 ( .A(n1306), .B(n1934), .C(n385), .Y(n2324) );
  OAI21X1 U2028 ( .A(n1306), .B(n1936), .C(n387), .Y(n2323) );
  OAI21X1 U2029 ( .A(n1306), .B(n1938), .C(n389), .Y(n2322) );
  OAI21X1 U2030 ( .A(n1306), .B(n1940), .C(n391), .Y(n2321) );
  OAI21X1 U2031 ( .A(n1306), .B(n1942), .C(n393), .Y(n2320) );
  OAI21X1 U2032 ( .A(n1308), .B(n1913), .C(n395), .Y(n2319) );
  OAI21X1 U2033 ( .A(n1308), .B(n1914), .C(n397), .Y(n2318) );
  OAI21X1 U2034 ( .A(n1308), .B(n1916), .C(n399), .Y(n2317) );
  OAI21X1 U2035 ( .A(n1308), .B(n1918), .C(n401), .Y(n2316) );
  OAI21X1 U2036 ( .A(n1308), .B(n1920), .C(n403), .Y(n2315) );
  OAI21X1 U2037 ( .A(n1308), .B(n1922), .C(n405), .Y(n2314) );
  OAI21X1 U2038 ( .A(n1308), .B(n1924), .C(n407), .Y(n2313) );
  OAI21X1 U2039 ( .A(n1308), .B(n1926), .C(n409), .Y(n2312) );
  OAI21X1 U2040 ( .A(n1308), .B(n1928), .C(n411), .Y(n2311) );
  OAI21X1 U2041 ( .A(n1308), .B(n1930), .C(n413), .Y(n2310) );
  OAI21X1 U2042 ( .A(n1308), .B(n1932), .C(n415), .Y(n2309) );
  OAI21X1 U2043 ( .A(n1308), .B(n1934), .C(n417), .Y(n2308) );
  OAI21X1 U2044 ( .A(n1308), .B(n1936), .C(n419), .Y(n2307) );
  OAI21X1 U2045 ( .A(n1308), .B(n1938), .C(n421), .Y(n2306) );
  OAI21X1 U2046 ( .A(n1308), .B(n1940), .C(n423), .Y(n2305) );
  OAI21X1 U2047 ( .A(n1308), .B(n1942), .C(n425), .Y(n2304) );
  OAI21X1 U2048 ( .A(n1887), .B(n1913), .C(n427), .Y(n2303) );
  OAI21X1 U2049 ( .A(n1887), .B(n1914), .C(n429), .Y(n2302) );
  OAI21X1 U2050 ( .A(n1887), .B(n1916), .C(n431), .Y(n2301) );
  OAI21X1 U2051 ( .A(n1887), .B(n1918), .C(n433), .Y(n2300) );
  OAI21X1 U2052 ( .A(n1887), .B(n1920), .C(n435), .Y(n2299) );
  OAI21X1 U2053 ( .A(n1887), .B(n1922), .C(n437), .Y(n2298) );
  OAI21X1 U2054 ( .A(n1887), .B(n1924), .C(n439), .Y(n2297) );
  OAI21X1 U2055 ( .A(n1887), .B(n1926), .C(n441), .Y(n2296) );
  OAI21X1 U2056 ( .A(n1887), .B(n1928), .C(n443), .Y(n2295) );
  OAI21X1 U2057 ( .A(n1887), .B(n1930), .C(n445), .Y(n2294) );
  OAI21X1 U2058 ( .A(n1887), .B(n1932), .C(n447), .Y(n2293) );
  OAI21X1 U2059 ( .A(n1887), .B(n1934), .C(n449), .Y(n2292) );
  OAI21X1 U2060 ( .A(n1887), .B(n1936), .C(n451), .Y(n2291) );
  OAI21X1 U2061 ( .A(n1887), .B(n1938), .C(n453), .Y(n2290) );
  OAI21X1 U2062 ( .A(n1887), .B(n1940), .C(n455), .Y(n2289) );
  OAI21X1 U2063 ( .A(n1887), .B(n1942), .C(n457), .Y(n2288) );
  NAND3X1 U2064 ( .A(n1951), .B(n2672), .C(n1952), .Y(n2152) );
  OAI21X1 U2065 ( .A(n1310), .B(n1912), .C(n459), .Y(n2287) );
  OAI21X1 U2066 ( .A(n1310), .B(n1914), .C(n461), .Y(n2286) );
  OAI21X1 U2067 ( .A(n1310), .B(n1916), .C(n463), .Y(n2285) );
  OAI21X1 U2068 ( .A(n1310), .B(n1918), .C(n465), .Y(n2284) );
  OAI21X1 U2069 ( .A(n1310), .B(n1920), .C(n467), .Y(n2283) );
  OAI21X1 U2070 ( .A(n1310), .B(n1922), .C(n469), .Y(n2282) );
  OAI21X1 U2071 ( .A(n1310), .B(n1924), .C(n471), .Y(n2281) );
  OAI21X1 U2072 ( .A(n1310), .B(n1926), .C(n473), .Y(n2280) );
  OAI21X1 U2073 ( .A(n1310), .B(n1928), .C(n475), .Y(n2279) );
  OAI21X1 U2074 ( .A(n1310), .B(n1930), .C(n477), .Y(n2278) );
  OAI21X1 U2075 ( .A(n1310), .B(n1932), .C(n479), .Y(n2277) );
  OAI21X1 U2076 ( .A(n1310), .B(n1934), .C(n481), .Y(n2276) );
  OAI21X1 U2077 ( .A(n1310), .B(n1936), .C(n483), .Y(n2275) );
  OAI21X1 U2078 ( .A(n1310), .B(n1938), .C(n485), .Y(n2274) );
  OAI21X1 U2079 ( .A(n1310), .B(n1940), .C(n487), .Y(n2273) );
  OAI21X1 U2080 ( .A(n1310), .B(n1942), .C(n489), .Y(n2272) );
  OAI21X1 U2081 ( .A(n1312), .B(n1913), .C(n491), .Y(n2271) );
  OAI21X1 U2082 ( .A(n1312), .B(n1914), .C(n493), .Y(n2270) );
  OAI21X1 U2083 ( .A(n1312), .B(n1916), .C(n495), .Y(n2269) );
  OAI21X1 U2084 ( .A(n1312), .B(n1918), .C(n497), .Y(n2268) );
  OAI21X1 U2085 ( .A(n1312), .B(n1920), .C(n499), .Y(n2267) );
  OAI21X1 U2086 ( .A(n1312), .B(n1922), .C(n501), .Y(n2266) );
  OAI21X1 U2087 ( .A(n1312), .B(n1924), .C(n503), .Y(n2265) );
  OAI21X1 U2088 ( .A(n1312), .B(n1926), .C(n505), .Y(n2264) );
  OAI21X1 U2089 ( .A(n1312), .B(n1928), .C(n507), .Y(n2263) );
  OAI21X1 U2090 ( .A(n1312), .B(n1930), .C(n509), .Y(n2262) );
  OAI21X1 U2091 ( .A(n1312), .B(n1932), .C(n511), .Y(n2261) );
  OAI21X1 U2092 ( .A(n1312), .B(n1934), .C(n513), .Y(n2260) );
  OAI21X1 U2093 ( .A(n1312), .B(n1936), .C(n515), .Y(n2259) );
  OAI21X1 U2094 ( .A(n1312), .B(n1938), .C(n517), .Y(n2258) );
  OAI21X1 U2095 ( .A(n1312), .B(n1940), .C(n519), .Y(n2257) );
  OAI21X1 U2096 ( .A(n1312), .B(n1942), .C(n521), .Y(n2256) );
  OAI21X1 U2097 ( .A(n1314), .B(n1912), .C(n523), .Y(n2255) );
  OAI21X1 U2098 ( .A(n1314), .B(n1914), .C(n525), .Y(n2254) );
  OAI21X1 U2099 ( .A(n1314), .B(n1916), .C(n527), .Y(n2253) );
  OAI21X1 U2100 ( .A(n1314), .B(n1918), .C(n529), .Y(n2252) );
  OAI21X1 U2101 ( .A(n1314), .B(n1920), .C(n531), .Y(n2251) );
  OAI21X1 U2102 ( .A(n1314), .B(n1922), .C(n533), .Y(n2250) );
  OAI21X1 U2103 ( .A(n1314), .B(n1924), .C(n535), .Y(n2249) );
  OAI21X1 U2104 ( .A(n1314), .B(n1926), .C(n537), .Y(n2248) );
  OAI21X1 U2105 ( .A(n1314), .B(n1928), .C(n539), .Y(n2247) );
  OAI21X1 U2106 ( .A(n1314), .B(n1930), .C(n541), .Y(n2246) );
  OAI21X1 U2107 ( .A(n1314), .B(n1932), .C(n543), .Y(n2245) );
  OAI21X1 U2108 ( .A(n1314), .B(n1934), .C(n545), .Y(n2244) );
  OAI21X1 U2109 ( .A(n1314), .B(n1936), .C(n547), .Y(n2243) );
  OAI21X1 U2110 ( .A(n1314), .B(n1938), .C(n549), .Y(n2242) );
  OAI21X1 U2111 ( .A(n1314), .B(n1940), .C(n551), .Y(n2241) );
  OAI21X1 U2112 ( .A(n1314), .B(n1942), .C(n553), .Y(n2240) );
  OAI21X1 U2113 ( .A(n1316), .B(n1913), .C(n555), .Y(n2239) );
  OAI21X1 U2114 ( .A(n1316), .B(n1914), .C(n557), .Y(n2238) );
  OAI21X1 U2115 ( .A(n1316), .B(n1916), .C(n559), .Y(n2237) );
  OAI21X1 U2116 ( .A(n1316), .B(n1918), .C(n561), .Y(n2236) );
  OAI21X1 U2117 ( .A(n1316), .B(n1920), .C(n563), .Y(n2235) );
  OAI21X1 U2118 ( .A(n1316), .B(n1922), .C(n565), .Y(n2234) );
  OAI21X1 U2119 ( .A(n1316), .B(n1924), .C(n567), .Y(n2233) );
  OAI21X1 U2120 ( .A(n1316), .B(n1926), .C(n569), .Y(n2232) );
  OAI21X1 U2121 ( .A(n1316), .B(n1928), .C(n571), .Y(n2231) );
  OAI21X1 U2122 ( .A(n1316), .B(n1930), .C(n573), .Y(n2230) );
  OAI21X1 U2123 ( .A(n1316), .B(n1932), .C(n575), .Y(n2229) );
  OAI21X1 U2124 ( .A(n1316), .B(n1934), .C(n577), .Y(n2228) );
  OAI21X1 U2125 ( .A(n1316), .B(n1936), .C(n579), .Y(n2227) );
  OAI21X1 U2126 ( .A(n1316), .B(n1938), .C(n581), .Y(n2226) );
  OAI21X1 U2127 ( .A(n1316), .B(n1940), .C(n583), .Y(n2225) );
  OAI21X1 U2128 ( .A(n1316), .B(n1942), .C(n585), .Y(n2224) );
  OAI21X1 U2129 ( .A(n1318), .B(n1912), .C(n587), .Y(n2223) );
  OAI21X1 U2130 ( .A(n1318), .B(n1914), .C(n589), .Y(n2222) );
  OAI21X1 U2131 ( .A(n1318), .B(n1916), .C(n591), .Y(n2221) );
  OAI21X1 U2132 ( .A(n1318), .B(n1918), .C(n593), .Y(n2220) );
  OAI21X1 U2133 ( .A(n1318), .B(n1920), .C(n595), .Y(n2219) );
  OAI21X1 U2134 ( .A(n1318), .B(n1922), .C(n597), .Y(n2218) );
  OAI21X1 U2135 ( .A(n1318), .B(n1924), .C(n599), .Y(n2217) );
  OAI21X1 U2136 ( .A(n1318), .B(n1926), .C(n601), .Y(n2216) );
  OAI21X1 U2137 ( .A(n1318), .B(n1928), .C(n603), .Y(n2215) );
  OAI21X1 U2138 ( .A(n1318), .B(n1930), .C(n605), .Y(n2214) );
  OAI21X1 U2139 ( .A(n1318), .B(n1932), .C(n607), .Y(n2213) );
  OAI21X1 U2140 ( .A(n1318), .B(n1934), .C(n609), .Y(n2212) );
  OAI21X1 U2141 ( .A(n1318), .B(n1936), .C(n611), .Y(n2211) );
  OAI21X1 U2142 ( .A(n1318), .B(n1938), .C(n613), .Y(n2210) );
  OAI21X1 U2143 ( .A(n1318), .B(n1940), .C(n615), .Y(n2209) );
  OAI21X1 U2144 ( .A(n1318), .B(n1942), .C(n617), .Y(n2208) );
  OAI21X1 U2145 ( .A(n1320), .B(n1913), .C(n619), .Y(n2207) );
  OAI21X1 U2146 ( .A(n1320), .B(n1914), .C(n621), .Y(n2206) );
  OAI21X1 U2147 ( .A(n1320), .B(n1916), .C(n623), .Y(n2205) );
  OAI21X1 U2148 ( .A(n1320), .B(n1918), .C(n625), .Y(n2204) );
  OAI21X1 U2149 ( .A(n1320), .B(n1920), .C(n627), .Y(n2203) );
  OAI21X1 U2150 ( .A(n1320), .B(n1922), .C(n629), .Y(n2202) );
  OAI21X1 U2151 ( .A(n1320), .B(n1924), .C(n631), .Y(n2201) );
  OAI21X1 U2152 ( .A(n1320), .B(n1926), .C(n633), .Y(n2200) );
  OAI21X1 U2153 ( .A(n1320), .B(n1928), .C(n635), .Y(n2199) );
  OAI21X1 U2154 ( .A(n1320), .B(n1930), .C(n637), .Y(n2198) );
  OAI21X1 U2155 ( .A(n1320), .B(n1932), .C(n639), .Y(n2197) );
  OAI21X1 U2156 ( .A(n1320), .B(n1934), .C(n641), .Y(n2196) );
  OAI21X1 U2157 ( .A(n1320), .B(n1936), .C(n643), .Y(n2195) );
  OAI21X1 U2158 ( .A(n1320), .B(n1938), .C(n645), .Y(n2194) );
  OAI21X1 U2159 ( .A(n1320), .B(n1940), .C(n647), .Y(n2193) );
  OAI21X1 U2160 ( .A(n1320), .B(n1942), .C(n649), .Y(n2192) );
  OAI21X1 U2161 ( .A(n1322), .B(n1912), .C(n1163), .Y(n2191) );
  OAI21X1 U2162 ( .A(n1322), .B(n1914), .C(n1165), .Y(n2190) );
  OAI21X1 U2163 ( .A(n1322), .B(n1916), .C(n1167), .Y(n2189) );
  OAI21X1 U2164 ( .A(n1322), .B(n1918), .C(n1169), .Y(n2188) );
  OAI21X1 U2165 ( .A(n1322), .B(n1920), .C(n1171), .Y(n2187) );
  OAI21X1 U2166 ( .A(n1322), .B(n1922), .C(n1173), .Y(n2186) );
  OAI21X1 U2167 ( .A(n1322), .B(n1924), .C(n1175), .Y(n2185) );
  OAI21X1 U2168 ( .A(n1322), .B(n1926), .C(n1177), .Y(n2184) );
  OAI21X1 U2169 ( .A(n1322), .B(n1928), .C(n1179), .Y(n2183) );
  OAI21X1 U2170 ( .A(n1322), .B(n1930), .C(n1181), .Y(n2182) );
  OAI21X1 U2171 ( .A(n1322), .B(n1932), .C(n1183), .Y(n2181) );
  OAI21X1 U2172 ( .A(n1322), .B(n1934), .C(n1185), .Y(n2180) );
  OAI21X1 U2173 ( .A(n1322), .B(n1936), .C(n1187), .Y(n2179) );
  OAI21X1 U2174 ( .A(n1322), .B(n1938), .C(n1189), .Y(n2178) );
  OAI21X1 U2175 ( .A(n1322), .B(n1940), .C(n1191), .Y(n2177) );
  OAI21X1 U2176 ( .A(n1322), .B(n1942), .C(n1193), .Y(n2176) );
  OAI21X1 U2177 ( .A(n1904), .B(n1913), .C(n1195), .Y(n2175) );
  OAI21X1 U2178 ( .A(n1904), .B(n1914), .C(n1197), .Y(n2174) );
  OAI21X1 U2179 ( .A(n1904), .B(n1916), .C(n1199), .Y(n2173) );
  OAI21X1 U2180 ( .A(n1904), .B(n1918), .C(n1201), .Y(n2172) );
  OAI21X1 U2181 ( .A(n1904), .B(n1920), .C(n1203), .Y(n2171) );
  OAI21X1 U2182 ( .A(n1904), .B(n1922), .C(n1205), .Y(n2170) );
  OAI21X1 U2183 ( .A(n1904), .B(n1924), .C(n1207), .Y(n2169) );
  OAI21X1 U2184 ( .A(n1904), .B(n1926), .C(n1209), .Y(n2168) );
  OAI21X1 U2185 ( .A(n1904), .B(n1928), .C(n1211), .Y(n2167) );
  OAI21X1 U2186 ( .A(n1904), .B(n1930), .C(n1213), .Y(n2166) );
  OAI21X1 U2187 ( .A(n1904), .B(n1932), .C(n1215), .Y(n2165) );
  OAI21X1 U2188 ( .A(n1904), .B(n1934), .C(n1217), .Y(n2164) );
  OAI21X1 U2189 ( .A(n1904), .B(n1936), .C(n1219), .Y(n2163) );
  OAI21X1 U2190 ( .A(n1904), .B(n1938), .C(n1221), .Y(n2162) );
  OAI21X1 U2191 ( .A(n1904), .B(n1940), .C(n1223), .Y(n2161) );
  OAI21X1 U2192 ( .A(n1904), .B(n1942), .C(n1225), .Y(n2160) );
endmodule


module memc_Size16_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n1852), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n1853), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n1854), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n1855), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n1856), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n1857), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n1858), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n1859), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n1860), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1861), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1862), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1863), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1864), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1865), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1866), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1867), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n1868), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n1869), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n1870), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n1871), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n1872), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n1873), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n1874), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n1875), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1876), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1877), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1878), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1879), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1880), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1881), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1882), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1883), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n1884), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n1885), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n1886), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n1887), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n1888), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n1889), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n1890), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n1891), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1892), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1893), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1894), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1895), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1896), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1897), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1898), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1899), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n1900), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n1901), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n1902), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n1903), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n1904), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n1905), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n1906), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n1907), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1908), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1909), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1910), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1911), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1912), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1913), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1914), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1915), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n1916), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n1917), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n1918), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n1919), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n1920), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n1921), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n1922), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n1923), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1924), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1925), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1926), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1927), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1928), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1929), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1930), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1931), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n1932), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n1933), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n1934), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n1935), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n1936), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n1937), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n1938), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n1939), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1940), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1941), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1942), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1943), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1944), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1945), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1946), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1947), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n1948), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n1949), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n1950), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n1951), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n1952), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n1953), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n1954), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n1955), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1956), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1957), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1958), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1959), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1960), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1961), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1962), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1963), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n1964), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n1965), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n1966), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n1967), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n1968), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n1969), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n1970), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n1971), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1972), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1973), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1974), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1975), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1976), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1977), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1978), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1979), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n1980), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n1981), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n1982), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n1983), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n1984), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n1985), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n1986), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n1987), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1988), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1989), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1990), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1991), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1992), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1993), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1994), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1995), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n1996), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n1997), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n1998), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n1999), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2000), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2001), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2002), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2003), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2004), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2005), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2006), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2007), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2008), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2009), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2010), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2011), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2012), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2013), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2014), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2015), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2016), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2017), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2018), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2019), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2020), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2021), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2022), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2023), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2024), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2025), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2026), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2027), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2028), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2029), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2030), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2031), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2032), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2033), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2034), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2035), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2036), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2037), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2038), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2039), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2040), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2041), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2042), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2043), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2044), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2045), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2046), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2047), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2048), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2049), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2050), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2051), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2052), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2053), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2054), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2055), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2056), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2057), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2058), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2059), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2060), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2061), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2062), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2063), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2064), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2065), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2066), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2067), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2068), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2069), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2070), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2071), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2072), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2073), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2074), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2075), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2076), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2077), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2078), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2079), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2080), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2081), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2082), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2083), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2084), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2085), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2086), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2087), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2088), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2089), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2090), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2091), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2092), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2093), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2094), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2095), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2096), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2097), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2098), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2099), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2100), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2101), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2102), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2103), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2104), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2105), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2106), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2107), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2108), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2109), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2110), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2111), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2112), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2113), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2114), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2115), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2116), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2117), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2118), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2119), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2120), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2121), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2122), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2123), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2124), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2125), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2126), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2127), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2128), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2129), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2130), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2131), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2132), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2133), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2134), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2135), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2136), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2137), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2138), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2139), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2140), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2141), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2142), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2143), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2144), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2145), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2146), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2147), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2148), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2149), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2150), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2151), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2152), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2153), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2154), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2155), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2156), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2157), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2158), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2159), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2160), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2161), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2162), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2163), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2164), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2165), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2166), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2167), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2168), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2169), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2170), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2171), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2172), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2173), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2174), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2175), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2176), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2177), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2178), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2179), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2180), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2181), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2182), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2183), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2184), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2185), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2186), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2187), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2188), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2189), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2190), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2191), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2192), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2193), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2194), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2195), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2196), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2197), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2198), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2199), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2200), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2201), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2202), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2203), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2204), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2205), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2206), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2207), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2208), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2209), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2210), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2211), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2212), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2213), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2214), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2215), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2216), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2217), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2218), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2219), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2220), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2221), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2222), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2223), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2224), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2225), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2226), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2227), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2228), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2229), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2230), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2231), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2232), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2233), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2234), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2235), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2236), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2237), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2238), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2239), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2240), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2241), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2242), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2243), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2244), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2245), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2246), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2247), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2248), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2249), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2250), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2251), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2252), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2253), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2254), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2255), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2256), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2257), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2258), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2259), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2260), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2261), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2262), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2263), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2264), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2265), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2266), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2267), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2268), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2269), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2270), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2271), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2272), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2273), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2274), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2275), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2276), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2277), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2278), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2279), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2280), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2281), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2282), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2283), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2284), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2285), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2286), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2287), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2288), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2289), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2290), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2291), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2292), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2293), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2294), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2295), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2296), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2297), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2298), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2299), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2300), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2301), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2302), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2303), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2304), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2305), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2306), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2307), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2308), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2309), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2310), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2311), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2312), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2313), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2314), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2315), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2316), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2317), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2318), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2319), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2320), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2321), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2322), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2323), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2324), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2325), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2326), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2327), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2328), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2329), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2330), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2331), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2332), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2333), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2334), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2335), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2336), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2337), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2338), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2339), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2340), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2341), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2342), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2343), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2344), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2345), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2346), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2347), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2348), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2349), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2350), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2351), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2352), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2353), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2354), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2355), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2356), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2357), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2358), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2359), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2360), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2361), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2362), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2363), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2364) );
  INVX2 U2 ( .A(n1192), .Y(n1205) );
  INVX2 U3 ( .A(n1318), .Y(n1207) );
  INVX1 U4 ( .A(n1210), .Y(n1192) );
  INVX2 U5 ( .A(n1318), .Y(n1206) );
  INVX2 U6 ( .A(n1192), .Y(n1198) );
  INVX2 U7 ( .A(n1192), .Y(n1209) );
  INVX2 U8 ( .A(n1192), .Y(n1194) );
  INVX2 U9 ( .A(n1192), .Y(n1200) );
  INVX2 U10 ( .A(n1192), .Y(n1199) );
  INVX2 U11 ( .A(n87), .Y(n1282) );
  INVX1 U12 ( .A(n642), .Y(N32) );
  INVX1 U13 ( .A(n643), .Y(N31) );
  INVX1 U14 ( .A(n644), .Y(N30) );
  INVX1 U15 ( .A(n645), .Y(N29) );
  INVX1 U16 ( .A(n646), .Y(N28) );
  INVX1 U17 ( .A(n647), .Y(N27) );
  INVX1 U18 ( .A(n648), .Y(N26) );
  INVX1 U19 ( .A(n649), .Y(N25) );
  INVX1 U20 ( .A(n650), .Y(N24) );
  INVX1 U21 ( .A(n1163), .Y(N23) );
  INVX1 U22 ( .A(n1164), .Y(N22) );
  INVX1 U23 ( .A(n1165), .Y(N21) );
  INVX1 U24 ( .A(n1166), .Y(N20) );
  INVX1 U25 ( .A(n1167), .Y(N19) );
  INVX1 U26 ( .A(n1168), .Y(N18) );
  INVX1 U27 ( .A(n1169), .Y(N17) );
  INVX1 U28 ( .A(n1210), .Y(n1193) );
  INVX1 U29 ( .A(n1191), .Y(n1180) );
  INVX1 U30 ( .A(n1191), .Y(n1181) );
  INVX1 U31 ( .A(n1191), .Y(n1182) );
  INVX1 U32 ( .A(n1179), .Y(n1183) );
  INVX2 U33 ( .A(n1192), .Y(n1201) );
  INVX1 U34 ( .A(n1179), .Y(n1184) );
  INVX2 U35 ( .A(n1318), .Y(n1202) );
  INVX2 U36 ( .A(n1192), .Y(n1203) );
  INVX2 U37 ( .A(n1179), .Y(n1185) );
  INVX2 U38 ( .A(n1192), .Y(n1204) );
  INVX1 U39 ( .A(n1178), .Y(n1186) );
  INVX1 U40 ( .A(n1178), .Y(n1187) );
  INVX2 U41 ( .A(n1178), .Y(n1188) );
  INVX2 U42 ( .A(n1178), .Y(n1189) );
  INVX2 U43 ( .A(n1179), .Y(n1190) );
  BUFX2 U44 ( .A(n9), .Y(n1211) );
  BUFX2 U45 ( .A(n9), .Y(n1212) );
  BUFX2 U46 ( .A(n26), .Y(n1213) );
  BUFX2 U47 ( .A(n26), .Y(n1214) );
  BUFX2 U48 ( .A(n28), .Y(n1215) );
  BUFX2 U49 ( .A(n28), .Y(n1216) );
  BUFX2 U50 ( .A(n30), .Y(n1217) );
  BUFX2 U51 ( .A(n30), .Y(n1218) );
  BUFX2 U52 ( .A(n32), .Y(n1219) );
  BUFX2 U53 ( .A(n32), .Y(n1220) );
  BUFX2 U54 ( .A(n34), .Y(n1221) );
  BUFX2 U55 ( .A(n34), .Y(n1222) );
  BUFX2 U56 ( .A(n36), .Y(n1223) );
  BUFX2 U57 ( .A(n36), .Y(n1224) );
  BUFX2 U58 ( .A(n38), .Y(n1226) );
  BUFX2 U59 ( .A(n38), .Y(n1227) );
  BUFX2 U60 ( .A(n40), .Y(n1228) );
  BUFX2 U61 ( .A(n40), .Y(n1229) );
  BUFX2 U62 ( .A(n42), .Y(n1230) );
  BUFX2 U63 ( .A(n42), .Y(n1231) );
  BUFX2 U64 ( .A(n44), .Y(n1232) );
  BUFX2 U65 ( .A(n44), .Y(n1233) );
  BUFX2 U66 ( .A(n46), .Y(n1234) );
  BUFX2 U67 ( .A(n46), .Y(n1235) );
  BUFX2 U68 ( .A(n48), .Y(n1236) );
  BUFX2 U69 ( .A(n48), .Y(n1237) );
  BUFX2 U70 ( .A(n50), .Y(n1238) );
  BUFX2 U71 ( .A(n50), .Y(n1239) );
  BUFX2 U72 ( .A(n52), .Y(n1240) );
  BUFX2 U73 ( .A(n52), .Y(n1241) );
  BUFX2 U74 ( .A(n54), .Y(n1243) );
  BUFX2 U75 ( .A(n54), .Y(n1244) );
  BUFX2 U76 ( .A(n56), .Y(n1245) );
  BUFX2 U77 ( .A(n56), .Y(n1246) );
  BUFX2 U78 ( .A(n58), .Y(n1247) );
  BUFX2 U79 ( .A(n58), .Y(n1248) );
  BUFX2 U80 ( .A(n60), .Y(n1249) );
  BUFX2 U81 ( .A(n60), .Y(n1250) );
  BUFX2 U82 ( .A(n62), .Y(n1251) );
  BUFX2 U83 ( .A(n62), .Y(n1252) );
  BUFX2 U84 ( .A(n64), .Y(n1253) );
  BUFX2 U85 ( .A(n64), .Y(n1254) );
  BUFX2 U86 ( .A(n66), .Y(n1255) );
  BUFX2 U87 ( .A(n66), .Y(n1256) );
  BUFX2 U88 ( .A(n68), .Y(n1257) );
  BUFX2 U89 ( .A(n68), .Y(n1258) );
  BUFX2 U90 ( .A(n70), .Y(n1260) );
  BUFX2 U91 ( .A(n70), .Y(n1261) );
  BUFX2 U92 ( .A(n72), .Y(n1262) );
  BUFX2 U93 ( .A(n72), .Y(n1263) );
  BUFX2 U94 ( .A(n74), .Y(n1264) );
  BUFX2 U95 ( .A(n74), .Y(n1265) );
  BUFX2 U96 ( .A(n76), .Y(n1266) );
  BUFX2 U97 ( .A(n76), .Y(n1267) );
  BUFX2 U98 ( .A(n78), .Y(n1268) );
  BUFX2 U99 ( .A(n78), .Y(n1269) );
  BUFX2 U100 ( .A(n80), .Y(n1270) );
  BUFX2 U101 ( .A(n80), .Y(n1271) );
  BUFX2 U102 ( .A(n82), .Y(n1272) );
  BUFX2 U103 ( .A(n82), .Y(n1273) );
  BUFX2 U104 ( .A(n84), .Y(n1274) );
  BUFX2 U105 ( .A(n84), .Y(n1275) );
  BUFX2 U106 ( .A(n86), .Y(n1277) );
  BUFX2 U107 ( .A(n86), .Y(n1278) );
  INVX1 U108 ( .A(n1318), .Y(n1210) );
  INVX1 U109 ( .A(n1319), .Y(n1191) );
  INVX1 U110 ( .A(N14), .Y(n1324) );
  INVX2 U111 ( .A(n1322), .Y(n1177) );
  INVX1 U112 ( .A(n1321), .Y(n1173) );
  INVX1 U113 ( .A(n1173), .Y(n1175) );
  INVX1 U114 ( .A(n1322), .Y(n1176) );
  INVX1 U115 ( .A(n1173), .Y(n1174) );
  INVX1 U116 ( .A(n1324), .Y(n1170) );
  INVX1 U117 ( .A(n1323), .Y(n1171) );
  INVX1 U118 ( .A(n1323), .Y(n1172) );
  INVX1 U119 ( .A(rst), .Y(n1316) );
  INVX1 U120 ( .A(n1319), .Y(n1179) );
  INVX1 U121 ( .A(n1319), .Y(n1178) );
  INVX1 U122 ( .A(n101), .Y(n1225) );
  INVX1 U123 ( .A(n102), .Y(n1242) );
  INVX1 U124 ( .A(n103), .Y(n1259) );
  INVX1 U125 ( .A(n104), .Y(n1276) );
  INVX4 U126 ( .A(n1282), .Y(n1280) );
  INVX4 U127 ( .A(n1282), .Y(n1281) );
  INVX1 U128 ( .A(n5), .Y(n4) );
  INVX2 U129 ( .A(n5), .Y(n1) );
  INVX1 U130 ( .A(write), .Y(n2) );
  INVX1 U131 ( .A(n2), .Y(n3) );
  INVX2 U132 ( .A(n5), .Y(n6) );
  OR2X2 U133 ( .A(write), .B(rst), .Y(n5) );
  AND2X2 U134 ( .A(\data_in<0> ), .B(n1280), .Y(n7) );
  AND2X2 U135 ( .A(n1279), .B(n105), .Y(n8) );
  INVX1 U136 ( .A(n8), .Y(n9) );
  AND2X2 U137 ( .A(\data_in<1> ), .B(n1281), .Y(n10) );
  AND2X2 U138 ( .A(\data_in<2> ), .B(n1280), .Y(n11) );
  AND2X2 U139 ( .A(\data_in<3> ), .B(n1280), .Y(n12) );
  AND2X2 U140 ( .A(\data_in<4> ), .B(n1281), .Y(n13) );
  AND2X2 U141 ( .A(\data_in<5> ), .B(n1280), .Y(n14) );
  AND2X2 U142 ( .A(\data_in<6> ), .B(n1281), .Y(n15) );
  AND2X2 U143 ( .A(\data_in<7> ), .B(n1280), .Y(n16) );
  AND2X2 U144 ( .A(\data_in<8> ), .B(n1281), .Y(n17) );
  AND2X2 U145 ( .A(\data_in<9> ), .B(n1280), .Y(n18) );
  AND2X2 U146 ( .A(\data_in<10> ), .B(n1281), .Y(n19) );
  AND2X2 U147 ( .A(\data_in<11> ), .B(n1281), .Y(n20) );
  AND2X2 U148 ( .A(\data_in<12> ), .B(n1281), .Y(n21) );
  AND2X2 U149 ( .A(\data_in<13> ), .B(n1281), .Y(n22) );
  AND2X2 U150 ( .A(\data_in<14> ), .B(n1281), .Y(n23) );
  AND2X2 U151 ( .A(\data_in<15> ), .B(n1281), .Y(n24) );
  AND2X2 U152 ( .A(n1279), .B(n107), .Y(n25) );
  INVX1 U153 ( .A(n25), .Y(n26) );
  AND2X2 U154 ( .A(n1279), .B(n109), .Y(n27) );
  INVX1 U155 ( .A(n27), .Y(n28) );
  AND2X2 U156 ( .A(n1279), .B(n111), .Y(n29) );
  INVX1 U157 ( .A(n29), .Y(n30) );
  AND2X2 U158 ( .A(n1279), .B(n113), .Y(n31) );
  INVX1 U159 ( .A(n31), .Y(n32) );
  AND2X2 U160 ( .A(n1279), .B(n115), .Y(n33) );
  INVX1 U161 ( .A(n33), .Y(n34) );
  AND2X2 U162 ( .A(n1279), .B(n117), .Y(n35) );
  INVX1 U163 ( .A(n35), .Y(n36) );
  AND2X2 U164 ( .A(n1279), .B(n101), .Y(n37) );
  INVX1 U165 ( .A(n37), .Y(n38) );
  AND2X2 U166 ( .A(n1279), .B(n119), .Y(n39) );
  INVX1 U167 ( .A(n39), .Y(n40) );
  AND2X2 U168 ( .A(n1279), .B(n121), .Y(n41) );
  INVX1 U169 ( .A(n41), .Y(n42) );
  AND2X2 U170 ( .A(n1279), .B(n123), .Y(n43) );
  INVX1 U171 ( .A(n43), .Y(n44) );
  AND2X2 U172 ( .A(n1279), .B(n125), .Y(n45) );
  INVX1 U173 ( .A(n45), .Y(n46) );
  AND2X2 U174 ( .A(n1280), .B(n127), .Y(n47) );
  INVX1 U175 ( .A(n47), .Y(n48) );
  AND2X2 U176 ( .A(n1280), .B(n129), .Y(n49) );
  INVX1 U177 ( .A(n49), .Y(n50) );
  AND2X2 U178 ( .A(n1280), .B(n131), .Y(n51) );
  INVX1 U179 ( .A(n51), .Y(n52) );
  AND2X2 U180 ( .A(n1280), .B(n102), .Y(n53) );
  INVX1 U181 ( .A(n53), .Y(n54) );
  AND2X2 U182 ( .A(n1280), .B(n133), .Y(n55) );
  INVX1 U183 ( .A(n55), .Y(n56) );
  AND2X2 U184 ( .A(n1280), .B(n135), .Y(n57) );
  INVX1 U185 ( .A(n57), .Y(n58) );
  AND2X2 U186 ( .A(n1280), .B(n137), .Y(n59) );
  INVX1 U187 ( .A(n59), .Y(n60) );
  AND2X2 U188 ( .A(n1280), .B(n139), .Y(n61) );
  INVX1 U189 ( .A(n61), .Y(n62) );
  AND2X2 U190 ( .A(n1280), .B(n141), .Y(n63) );
  INVX1 U191 ( .A(n63), .Y(n64) );
  AND2X2 U192 ( .A(n1280), .B(n143), .Y(n65) );
  INVX1 U193 ( .A(n65), .Y(n66) );
  AND2X2 U194 ( .A(n1280), .B(n145), .Y(n67) );
  INVX1 U195 ( .A(n67), .Y(n68) );
  AND2X2 U196 ( .A(n1281), .B(n103), .Y(n69) );
  INVX1 U197 ( .A(n69), .Y(n70) );
  AND2X2 U198 ( .A(n1281), .B(n147), .Y(n71) );
  INVX1 U199 ( .A(n71), .Y(n72) );
  AND2X2 U200 ( .A(n1281), .B(n149), .Y(n73) );
  INVX1 U201 ( .A(n73), .Y(n74) );
  AND2X2 U202 ( .A(n1281), .B(n151), .Y(n75) );
  INVX1 U203 ( .A(n75), .Y(n76) );
  AND2X2 U204 ( .A(n1281), .B(n153), .Y(n77) );
  INVX1 U205 ( .A(n77), .Y(n78) );
  AND2X2 U206 ( .A(n1281), .B(n155), .Y(n79) );
  INVX1 U207 ( .A(n79), .Y(n80) );
  AND2X2 U208 ( .A(n1281), .B(n157), .Y(n81) );
  INVX1 U209 ( .A(n81), .Y(n82) );
  AND2X2 U210 ( .A(n1281), .B(n159), .Y(n83) );
  INVX1 U211 ( .A(n83), .Y(n84) );
  AND2X2 U212 ( .A(n1280), .B(n104), .Y(n85) );
  INVX1 U213 ( .A(n85), .Y(n86) );
  AND2X2 U214 ( .A(n3), .B(n1316), .Y(n87) );
  INVX1 U215 ( .A(n1320), .Y(n1319) );
  INVX1 U216 ( .A(n1318), .Y(n1317) );
  INVX1 U217 ( .A(N13), .Y(n1323) );
  AND2X1 U218 ( .A(n1321), .B(n1319), .Y(n88) );
  INVX1 U219 ( .A(n1322), .Y(n1321) );
  AND2X1 U220 ( .A(n2364), .B(N14), .Y(n89) );
  INVX2 U221 ( .A(n1283), .Y(n1279) );
  BUFX2 U222 ( .A(n1357), .Y(n90) );
  INVX1 U223 ( .A(n90), .Y(n1749) );
  BUFX2 U224 ( .A(n1374), .Y(n91) );
  INVX1 U225 ( .A(n91), .Y(n1766) );
  BUFX2 U226 ( .A(n1391), .Y(n92) );
  INVX1 U227 ( .A(n92), .Y(n1783) );
  BUFX2 U228 ( .A(n1408), .Y(n93) );
  INVX1 U229 ( .A(n93), .Y(n1800) );
  BUFX2 U230 ( .A(n1425), .Y(n94) );
  INVX1 U231 ( .A(n94), .Y(n1817) );
  BUFX2 U232 ( .A(n1586), .Y(n95) );
  INVX1 U233 ( .A(n95), .Y(n1699) );
  BUFX2 U234 ( .A(n1716), .Y(n96) );
  INVX1 U235 ( .A(n96), .Y(n1834) );
  AND2X1 U236 ( .A(n1317), .B(n88), .Y(n97) );
  AND2X1 U237 ( .A(n1172), .B(n89), .Y(n98) );
  INVX1 U238 ( .A(n87), .Y(n1283) );
  AND2X1 U239 ( .A(n1318), .B(n88), .Y(n99) );
  AND2X1 U240 ( .A(n1323), .B(n89), .Y(n100) );
  AND2X1 U241 ( .A(n98), .B(n1835), .Y(n101) );
  AND2X1 U242 ( .A(n1835), .B(n100), .Y(n102) );
  AND2X1 U243 ( .A(n1835), .B(n1699), .Y(n103) );
  AND2X1 U244 ( .A(n1835), .B(n1834), .Y(n104) );
  AND2X1 U245 ( .A(n97), .B(n98), .Y(n105) );
  INVX1 U246 ( .A(n105), .Y(n106) );
  AND2X1 U247 ( .A(n98), .B(n99), .Y(n107) );
  INVX1 U248 ( .A(n107), .Y(n108) );
  AND2X1 U249 ( .A(n98), .B(n1749), .Y(n109) );
  INVX1 U250 ( .A(n109), .Y(n110) );
  AND2X1 U251 ( .A(n98), .B(n1766), .Y(n111) );
  INVX1 U252 ( .A(n111), .Y(n112) );
  AND2X1 U253 ( .A(n98), .B(n1783), .Y(n113) );
  INVX1 U254 ( .A(n113), .Y(n114) );
  AND2X1 U255 ( .A(n98), .B(n1800), .Y(n115) );
  INVX1 U256 ( .A(n115), .Y(n116) );
  AND2X1 U257 ( .A(n98), .B(n1817), .Y(n117) );
  INVX1 U258 ( .A(n117), .Y(n118) );
  AND2X1 U259 ( .A(n97), .B(n100), .Y(n119) );
  INVX1 U260 ( .A(n119), .Y(n120) );
  AND2X1 U261 ( .A(n99), .B(n100), .Y(n121) );
  INVX1 U262 ( .A(n121), .Y(n122) );
  AND2X1 U263 ( .A(n1749), .B(n100), .Y(n123) );
  INVX1 U264 ( .A(n123), .Y(n124) );
  AND2X1 U265 ( .A(n1766), .B(n100), .Y(n125) );
  INVX1 U266 ( .A(n125), .Y(n126) );
  AND2X1 U267 ( .A(n1783), .B(n100), .Y(n127) );
  INVX1 U268 ( .A(n127), .Y(n128) );
  AND2X1 U269 ( .A(n1800), .B(n100), .Y(n129) );
  INVX1 U270 ( .A(n129), .Y(n130) );
  AND2X1 U271 ( .A(n1817), .B(n100), .Y(n131) );
  INVX1 U272 ( .A(n131), .Y(n132) );
  AND2X1 U273 ( .A(n97), .B(n1699), .Y(n133) );
  INVX1 U274 ( .A(n133), .Y(n134) );
  AND2X1 U275 ( .A(n99), .B(n1699), .Y(n135) );
  INVX1 U276 ( .A(n135), .Y(n136) );
  AND2X1 U277 ( .A(n1749), .B(n1699), .Y(n137) );
  INVX1 U278 ( .A(n137), .Y(n138) );
  AND2X1 U279 ( .A(n1766), .B(n1699), .Y(n139) );
  INVX1 U280 ( .A(n139), .Y(n140) );
  AND2X1 U281 ( .A(n1783), .B(n1699), .Y(n141) );
  INVX1 U282 ( .A(n141), .Y(n142) );
  AND2X1 U283 ( .A(n1800), .B(n1699), .Y(n143) );
  INVX1 U284 ( .A(n143), .Y(n144) );
  AND2X1 U285 ( .A(n1817), .B(n1699), .Y(n145) );
  INVX1 U286 ( .A(n145), .Y(n146) );
  AND2X1 U287 ( .A(n97), .B(n1834), .Y(n147) );
  INVX1 U288 ( .A(n147), .Y(n148) );
  AND2X1 U289 ( .A(n99), .B(n1834), .Y(n149) );
  INVX1 U290 ( .A(n149), .Y(n150) );
  AND2X1 U291 ( .A(n1749), .B(n1834), .Y(n151) );
  INVX1 U292 ( .A(n151), .Y(n152) );
  AND2X1 U293 ( .A(n1766), .B(n1834), .Y(n153) );
  INVX1 U294 ( .A(n153), .Y(n154) );
  AND2X1 U295 ( .A(n1783), .B(n1834), .Y(n155) );
  INVX1 U296 ( .A(n155), .Y(n156) );
  AND2X1 U297 ( .A(n1800), .B(n1834), .Y(n157) );
  INVX1 U298 ( .A(n157), .Y(n158) );
  AND2X1 U299 ( .A(n1817), .B(n1834), .Y(n159) );
  INVX1 U300 ( .A(n159), .Y(n160) );
  MUX2X1 U301 ( .B(n162), .A(n163), .S(n1180), .Y(n161) );
  MUX2X1 U302 ( .B(n165), .A(n166), .S(n1180), .Y(n164) );
  MUX2X1 U303 ( .B(n168), .A(n169), .S(n1180), .Y(n167) );
  MUX2X1 U304 ( .B(n171), .A(n172), .S(n1180), .Y(n170) );
  MUX2X1 U305 ( .B(n174), .A(n175), .S(n1172), .Y(n173) );
  MUX2X1 U306 ( .B(n177), .A(n178), .S(n1180), .Y(n176) );
  MUX2X1 U307 ( .B(n180), .A(n181), .S(n1180), .Y(n179) );
  MUX2X1 U308 ( .B(n183), .A(n184), .S(n1180), .Y(n182) );
  MUX2X1 U309 ( .B(n186), .A(n187), .S(n1180), .Y(n185) );
  MUX2X1 U310 ( .B(n189), .A(n190), .S(n1172), .Y(n188) );
  MUX2X1 U311 ( .B(n192), .A(n193), .S(n1181), .Y(n191) );
  MUX2X1 U312 ( .B(n195), .A(n196), .S(n1181), .Y(n194) );
  MUX2X1 U313 ( .B(n198), .A(n199), .S(n1181), .Y(n197) );
  MUX2X1 U314 ( .B(n201), .A(n202), .S(n1181), .Y(n200) );
  MUX2X1 U315 ( .B(n204), .A(n205), .S(n1172), .Y(n203) );
  MUX2X1 U316 ( .B(n207), .A(n208), .S(n1181), .Y(n206) );
  MUX2X1 U317 ( .B(n210), .A(n211), .S(n1181), .Y(n209) );
  MUX2X1 U318 ( .B(n213), .A(n215), .S(n1181), .Y(n212) );
  MUX2X1 U319 ( .B(n217), .A(n218), .S(n1181), .Y(n216) );
  MUX2X1 U320 ( .B(n220), .A(n221), .S(n1172), .Y(n219) );
  MUX2X1 U321 ( .B(n223), .A(n224), .S(n1181), .Y(n222) );
  MUX2X1 U322 ( .B(n226), .A(n227), .S(n1181), .Y(n225) );
  MUX2X1 U323 ( .B(n229), .A(n230), .S(n1181), .Y(n228) );
  MUX2X1 U324 ( .B(n232), .A(n233), .S(n1181), .Y(n231) );
  MUX2X1 U325 ( .B(n235), .A(n236), .S(n1172), .Y(n234) );
  MUX2X1 U326 ( .B(n238), .A(n239), .S(n1182), .Y(n237) );
  MUX2X1 U327 ( .B(n241), .A(n242), .S(n1182), .Y(n240) );
  MUX2X1 U328 ( .B(n244), .A(n245), .S(n1182), .Y(n243) );
  MUX2X1 U329 ( .B(n247), .A(n248), .S(n1182), .Y(n246) );
  MUX2X1 U330 ( .B(n250), .A(n251), .S(n1172), .Y(n249) );
  MUX2X1 U331 ( .B(n253), .A(n254), .S(n1182), .Y(n252) );
  MUX2X1 U332 ( .B(n256), .A(n257), .S(n1182), .Y(n255) );
  MUX2X1 U333 ( .B(n259), .A(n260), .S(n1182), .Y(n258) );
  MUX2X1 U334 ( .B(n262), .A(n263), .S(n1182), .Y(n261) );
  MUX2X1 U335 ( .B(n265), .A(n266), .S(n1172), .Y(n264) );
  MUX2X1 U336 ( .B(n268), .A(n269), .S(n1182), .Y(n267) );
  MUX2X1 U337 ( .B(n271), .A(n272), .S(n1182), .Y(n270) );
  MUX2X1 U338 ( .B(n274), .A(n275), .S(n1182), .Y(n273) );
  MUX2X1 U339 ( .B(n277), .A(n278), .S(n1182), .Y(n276) );
  MUX2X1 U340 ( .B(n280), .A(n281), .S(n1172), .Y(n279) );
  MUX2X1 U341 ( .B(n283), .A(n284), .S(n1183), .Y(n282) );
  MUX2X1 U342 ( .B(n286), .A(n287), .S(n1183), .Y(n285) );
  MUX2X1 U343 ( .B(n289), .A(n290), .S(n1183), .Y(n288) );
  MUX2X1 U344 ( .B(n292), .A(n293), .S(n1183), .Y(n291) );
  MUX2X1 U345 ( .B(n295), .A(n296), .S(n1172), .Y(n294) );
  MUX2X1 U346 ( .B(n298), .A(n299), .S(n1183), .Y(n297) );
  MUX2X1 U347 ( .B(n301), .A(n302), .S(n1183), .Y(n300) );
  MUX2X1 U348 ( .B(n304), .A(n305), .S(n1183), .Y(n303) );
  MUX2X1 U349 ( .B(n307), .A(n308), .S(n1183), .Y(n306) );
  MUX2X1 U350 ( .B(n310), .A(n311), .S(n1172), .Y(n309) );
  MUX2X1 U351 ( .B(n313), .A(n314), .S(n1183), .Y(n312) );
  MUX2X1 U352 ( .B(n316), .A(n317), .S(n1183), .Y(n315) );
  MUX2X1 U353 ( .B(n319), .A(n320), .S(n1183), .Y(n318) );
  MUX2X1 U354 ( .B(n322), .A(n323), .S(n1183), .Y(n321) );
  MUX2X1 U355 ( .B(n325), .A(n326), .S(n1172), .Y(n324) );
  MUX2X1 U356 ( .B(n328), .A(n329), .S(n1184), .Y(n327) );
  MUX2X1 U357 ( .B(n331), .A(n332), .S(n1184), .Y(n330) );
  MUX2X1 U358 ( .B(n334), .A(n335), .S(n1184), .Y(n333) );
  MUX2X1 U359 ( .B(n337), .A(n338), .S(n1184), .Y(n336) );
  MUX2X1 U360 ( .B(n340), .A(n341), .S(n1172), .Y(n339) );
  MUX2X1 U361 ( .B(n343), .A(n344), .S(n1184), .Y(n342) );
  MUX2X1 U362 ( .B(n346), .A(n347), .S(n1184), .Y(n345) );
  MUX2X1 U363 ( .B(n349), .A(n350), .S(n1184), .Y(n348) );
  MUX2X1 U364 ( .B(n352), .A(n353), .S(n1184), .Y(n351) );
  MUX2X1 U365 ( .B(n355), .A(n356), .S(n1171), .Y(n354) );
  MUX2X1 U366 ( .B(n358), .A(n359), .S(n1184), .Y(n357) );
  MUX2X1 U367 ( .B(n361), .A(n362), .S(n1184), .Y(n360) );
  MUX2X1 U368 ( .B(n364), .A(n365), .S(n1184), .Y(n363) );
  MUX2X1 U369 ( .B(n367), .A(n368), .S(n1184), .Y(n366) );
  MUX2X1 U370 ( .B(n370), .A(n371), .S(n1171), .Y(n369) );
  MUX2X1 U371 ( .B(n373), .A(n374), .S(n1185), .Y(n372) );
  MUX2X1 U372 ( .B(n376), .A(n377), .S(n1185), .Y(n375) );
  MUX2X1 U373 ( .B(n379), .A(n380), .S(n1185), .Y(n378) );
  MUX2X1 U374 ( .B(n382), .A(n383), .S(n1185), .Y(n381) );
  MUX2X1 U375 ( .B(n385), .A(n386), .S(n1171), .Y(n384) );
  MUX2X1 U376 ( .B(n388), .A(n389), .S(n1185), .Y(n387) );
  MUX2X1 U377 ( .B(n391), .A(n392), .S(n1185), .Y(n390) );
  MUX2X1 U378 ( .B(n394), .A(n395), .S(n1185), .Y(n393) );
  MUX2X1 U379 ( .B(n397), .A(n398), .S(n1185), .Y(n396) );
  MUX2X1 U380 ( .B(n400), .A(n401), .S(n1171), .Y(n399) );
  MUX2X1 U381 ( .B(n403), .A(n404), .S(n1185), .Y(n402) );
  MUX2X1 U382 ( .B(n406), .A(n407), .S(n1185), .Y(n405) );
  MUX2X1 U383 ( .B(n409), .A(n410), .S(n1185), .Y(n408) );
  MUX2X1 U384 ( .B(n412), .A(n413), .S(n1185), .Y(n411) );
  MUX2X1 U385 ( .B(n415), .A(n416), .S(n1171), .Y(n414) );
  MUX2X1 U386 ( .B(n418), .A(n419), .S(n1186), .Y(n417) );
  MUX2X1 U387 ( .B(n421), .A(n422), .S(n1186), .Y(n420) );
  MUX2X1 U388 ( .B(n424), .A(n425), .S(n1186), .Y(n423) );
  MUX2X1 U389 ( .B(n427), .A(n428), .S(n1186), .Y(n426) );
  MUX2X1 U390 ( .B(n430), .A(n431), .S(n1171), .Y(n429) );
  MUX2X1 U391 ( .B(n433), .A(n434), .S(n1186), .Y(n432) );
  MUX2X1 U392 ( .B(n436), .A(n437), .S(n1186), .Y(n435) );
  MUX2X1 U393 ( .B(n439), .A(n440), .S(n1186), .Y(n438) );
  MUX2X1 U394 ( .B(n442), .A(n443), .S(n1186), .Y(n441) );
  MUX2X1 U395 ( .B(n445), .A(n446), .S(n1171), .Y(n444) );
  MUX2X1 U396 ( .B(n448), .A(n449), .S(n1186), .Y(n447) );
  MUX2X1 U397 ( .B(n451), .A(n452), .S(n1186), .Y(n450) );
  MUX2X1 U398 ( .B(n454), .A(n455), .S(n1186), .Y(n453) );
  MUX2X1 U399 ( .B(n457), .A(n458), .S(n1186), .Y(n456) );
  MUX2X1 U400 ( .B(n460), .A(n461), .S(n1171), .Y(n459) );
  MUX2X1 U401 ( .B(n463), .A(n464), .S(n1187), .Y(n462) );
  MUX2X1 U402 ( .B(n466), .A(n467), .S(n1187), .Y(n465) );
  MUX2X1 U403 ( .B(n469), .A(n470), .S(n1187), .Y(n468) );
  MUX2X1 U404 ( .B(n472), .A(n473), .S(n1187), .Y(n471) );
  MUX2X1 U405 ( .B(n475), .A(n476), .S(n1171), .Y(n474) );
  MUX2X1 U406 ( .B(n478), .A(n479), .S(n1187), .Y(n477) );
  MUX2X1 U407 ( .B(n481), .A(n482), .S(n1187), .Y(n480) );
  MUX2X1 U408 ( .B(n484), .A(n485), .S(n1187), .Y(n483) );
  MUX2X1 U409 ( .B(n487), .A(n488), .S(n1187), .Y(n486) );
  MUX2X1 U410 ( .B(n490), .A(n491), .S(n1171), .Y(n489) );
  MUX2X1 U411 ( .B(n493), .A(n494), .S(n1187), .Y(n492) );
  MUX2X1 U412 ( .B(n496), .A(n497), .S(n1187), .Y(n495) );
  MUX2X1 U413 ( .B(n499), .A(n500), .S(n1187), .Y(n498) );
  MUX2X1 U414 ( .B(n502), .A(n503), .S(n1187), .Y(n501) );
  MUX2X1 U415 ( .B(n505), .A(n506), .S(n1171), .Y(n504) );
  MUX2X1 U416 ( .B(n508), .A(n509), .S(n1188), .Y(n507) );
  MUX2X1 U417 ( .B(n511), .A(n512), .S(n1188), .Y(n510) );
  MUX2X1 U418 ( .B(n514), .A(n515), .S(n1188), .Y(n513) );
  MUX2X1 U419 ( .B(n517), .A(n518), .S(n1188), .Y(n516) );
  MUX2X1 U420 ( .B(n520), .A(n521), .S(n1171), .Y(n519) );
  MUX2X1 U421 ( .B(n523), .A(n524), .S(n1188), .Y(n522) );
  MUX2X1 U422 ( .B(n526), .A(n527), .S(n1188), .Y(n525) );
  MUX2X1 U423 ( .B(n529), .A(n530), .S(n1188), .Y(n528) );
  MUX2X1 U424 ( .B(n532), .A(n533), .S(n1188), .Y(n531) );
  MUX2X1 U425 ( .B(n535), .A(n536), .S(n1171), .Y(n534) );
  MUX2X1 U426 ( .B(n538), .A(n539), .S(n1188), .Y(n537) );
  MUX2X1 U427 ( .B(n541), .A(n542), .S(n1188), .Y(n540) );
  MUX2X1 U428 ( .B(n544), .A(n545), .S(n1188), .Y(n543) );
  MUX2X1 U429 ( .B(n547), .A(n548), .S(n1188), .Y(n546) );
  MUX2X1 U430 ( .B(n550), .A(n551), .S(n1171), .Y(n549) );
  MUX2X1 U431 ( .B(n553), .A(n554), .S(n1189), .Y(n552) );
  MUX2X1 U432 ( .B(n556), .A(n557), .S(n1189), .Y(n555) );
  MUX2X1 U433 ( .B(n559), .A(n560), .S(n1189), .Y(n558) );
  MUX2X1 U434 ( .B(n562), .A(n563), .S(n1189), .Y(n561) );
  MUX2X1 U435 ( .B(n565), .A(n566), .S(n1171), .Y(n564) );
  MUX2X1 U436 ( .B(n568), .A(n569), .S(n1189), .Y(n567) );
  MUX2X1 U437 ( .B(n571), .A(n572), .S(n1189), .Y(n570) );
  MUX2X1 U438 ( .B(n574), .A(n575), .S(n1189), .Y(n573) );
  MUX2X1 U439 ( .B(n577), .A(n578), .S(n1189), .Y(n576) );
  MUX2X1 U440 ( .B(n580), .A(n581), .S(n1171), .Y(n579) );
  MUX2X1 U441 ( .B(n583), .A(n584), .S(n1189), .Y(n582) );
  MUX2X1 U442 ( .B(n586), .A(n587), .S(n1189), .Y(n585) );
  MUX2X1 U443 ( .B(n589), .A(n590), .S(n1189), .Y(n588) );
  MUX2X1 U444 ( .B(n592), .A(n593), .S(n1189), .Y(n591) );
  MUX2X1 U445 ( .B(n595), .A(n596), .S(n1172), .Y(n594) );
  MUX2X1 U446 ( .B(n598), .A(n599), .S(n1190), .Y(n597) );
  MUX2X1 U447 ( .B(n601), .A(n602), .S(n1190), .Y(n600) );
  MUX2X1 U448 ( .B(n604), .A(n605), .S(n1190), .Y(n603) );
  MUX2X1 U449 ( .B(n607), .A(n608), .S(n1190), .Y(n606) );
  MUX2X1 U450 ( .B(n610), .A(n611), .S(n1171), .Y(n609) );
  MUX2X1 U451 ( .B(n613), .A(n614), .S(n1190), .Y(n612) );
  MUX2X1 U452 ( .B(n616), .A(n617), .S(n1190), .Y(n615) );
  MUX2X1 U453 ( .B(n619), .A(n620), .S(n1190), .Y(n618) );
  MUX2X1 U454 ( .B(n622), .A(n623), .S(n1190), .Y(n621) );
  MUX2X1 U455 ( .B(n625), .A(n626), .S(n1171), .Y(n624) );
  MUX2X1 U456 ( .B(n628), .A(n629), .S(n1190), .Y(n627) );
  MUX2X1 U457 ( .B(n631), .A(n632), .S(n1190), .Y(n630) );
  MUX2X1 U458 ( .B(n634), .A(n635), .S(n1190), .Y(n633) );
  MUX2X1 U459 ( .B(n637), .A(n638), .S(n1190), .Y(n636) );
  MUX2X1 U460 ( .B(n640), .A(n641), .S(n1171), .Y(n639) );
  MUX2X1 U461 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1199), .Y(n163) );
  MUX2X1 U462 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1200), .Y(n162) );
  MUX2X1 U463 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1200), .Y(n166) );
  MUX2X1 U464 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1199), .Y(n165) );
  MUX2X1 U465 ( .B(n164), .A(n161), .S(n1177), .Y(n175) );
  MUX2X1 U466 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1194), .Y(n169) );
  MUX2X1 U467 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1194), .Y(n168) );
  MUX2X1 U468 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1194), .Y(n172) );
  MUX2X1 U469 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1194), .Y(n171) );
  MUX2X1 U470 ( .B(n170), .A(n167), .S(n1177), .Y(n174) );
  MUX2X1 U471 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1194), .Y(n178) );
  MUX2X1 U472 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1194), .Y(n177) );
  MUX2X1 U473 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1194), .Y(n181) );
  MUX2X1 U474 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1194), .Y(n180) );
  MUX2X1 U475 ( .B(n179), .A(n176), .S(n1177), .Y(n190) );
  MUX2X1 U476 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1194), .Y(n184) );
  MUX2X1 U477 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1194), .Y(n183) );
  MUX2X1 U478 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1194), .Y(n187) );
  MUX2X1 U479 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1194), .Y(n186) );
  MUX2X1 U480 ( .B(n185), .A(n182), .S(n1177), .Y(n189) );
  MUX2X1 U481 ( .B(n188), .A(n173), .S(n1170), .Y(n642) );
  MUX2X1 U482 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1209), .Y(n193) );
  MUX2X1 U483 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1208), .Y(n192) );
  MUX2X1 U484 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1209), .Y(n196) );
  MUX2X1 U485 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1209), .Y(n195) );
  MUX2X1 U486 ( .B(n194), .A(n191), .S(n1177), .Y(n205) );
  MUX2X1 U487 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1194), .Y(n199) );
  MUX2X1 U488 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1198), .Y(n198) );
  MUX2X1 U489 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1198), .Y(n202) );
  MUX2X1 U490 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1198), .Y(n201) );
  MUX2X1 U491 ( .B(n200), .A(n197), .S(n1177), .Y(n204) );
  MUX2X1 U492 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1209), .Y(n208) );
  MUX2X1 U493 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1194), .Y(n207) );
  MUX2X1 U494 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1198), .Y(n211) );
  MUX2X1 U495 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1209), .Y(n210) );
  MUX2X1 U496 ( .B(n209), .A(n206), .S(n1177), .Y(n221) );
  MUX2X1 U497 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1195), .Y(n215) );
  MUX2X1 U498 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1195), .Y(n213) );
  MUX2X1 U499 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1195), .Y(n218) );
  MUX2X1 U500 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1195), .Y(n217) );
  MUX2X1 U501 ( .B(n216), .A(n212), .S(n1177), .Y(n220) );
  MUX2X1 U502 ( .B(n219), .A(n203), .S(n1170), .Y(n643) );
  MUX2X1 U503 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1195), .Y(n224) );
  MUX2X1 U504 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1195), .Y(n223) );
  MUX2X1 U505 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1195), .Y(n227) );
  MUX2X1 U506 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1195), .Y(n226) );
  MUX2X1 U507 ( .B(n225), .A(n222), .S(n1177), .Y(n236) );
  MUX2X1 U508 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1195), .Y(n230) );
  MUX2X1 U509 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1195), .Y(n229) );
  MUX2X1 U510 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1195), .Y(n233) );
  MUX2X1 U511 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1195), .Y(n232) );
  MUX2X1 U512 ( .B(n231), .A(n228), .S(n1177), .Y(n235) );
  MUX2X1 U513 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1196), .Y(n239) );
  MUX2X1 U514 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1196), .Y(n238) );
  MUX2X1 U515 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1196), .Y(n242) );
  MUX2X1 U516 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1196), .Y(n241) );
  MUX2X1 U517 ( .B(n240), .A(n237), .S(n1177), .Y(n251) );
  MUX2X1 U518 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1196), .Y(n245) );
  MUX2X1 U519 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1196), .Y(n244) );
  MUX2X1 U520 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1196), .Y(n248) );
  MUX2X1 U521 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1196), .Y(n247) );
  MUX2X1 U522 ( .B(n246), .A(n243), .S(n1177), .Y(n250) );
  MUX2X1 U523 ( .B(n249), .A(n234), .S(n1170), .Y(n644) );
  MUX2X1 U524 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1196), .Y(n254) );
  MUX2X1 U525 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1196), .Y(n253) );
  MUX2X1 U526 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1196), .Y(n257) );
  MUX2X1 U527 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1196), .Y(n256) );
  MUX2X1 U528 ( .B(n255), .A(n252), .S(n1176), .Y(n266) );
  MUX2X1 U529 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1197), .Y(n260) );
  MUX2X1 U530 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1197), .Y(n259) );
  MUX2X1 U531 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1197), .Y(n263) );
  MUX2X1 U532 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1197), .Y(n262) );
  MUX2X1 U533 ( .B(n261), .A(n258), .S(n1176), .Y(n265) );
  MUX2X1 U534 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1197), .Y(n269) );
  MUX2X1 U535 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1197), .Y(n268) );
  MUX2X1 U536 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1197), .Y(n272) );
  MUX2X1 U537 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1197), .Y(n271) );
  MUX2X1 U538 ( .B(n270), .A(n267), .S(n1176), .Y(n281) );
  MUX2X1 U539 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1197), .Y(n275) );
  MUX2X1 U540 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1197), .Y(n274) );
  MUX2X1 U541 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1197), .Y(n278) );
  MUX2X1 U542 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1197), .Y(n277) );
  MUX2X1 U543 ( .B(n276), .A(n273), .S(n1176), .Y(n280) );
  MUX2X1 U544 ( .B(n279), .A(n264), .S(n1170), .Y(n645) );
  MUX2X1 U545 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1198), .Y(n284) );
  MUX2X1 U546 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1198), .Y(n283) );
  MUX2X1 U547 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1198), .Y(n287) );
  MUX2X1 U548 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1198), .Y(n286) );
  MUX2X1 U549 ( .B(n285), .A(n282), .S(n1176), .Y(n296) );
  MUX2X1 U550 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1198), .Y(n290) );
  MUX2X1 U551 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1198), .Y(n289) );
  MUX2X1 U552 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1198), .Y(n293) );
  MUX2X1 U553 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1198), .Y(n292) );
  MUX2X1 U554 ( .B(n291), .A(n288), .S(n1176), .Y(n295) );
  MUX2X1 U555 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1198), .Y(n299) );
  MUX2X1 U556 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1198), .Y(n298) );
  MUX2X1 U557 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1198), .Y(n302) );
  MUX2X1 U558 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1198), .Y(n301) );
  MUX2X1 U559 ( .B(n300), .A(n297), .S(n1176), .Y(n311) );
  MUX2X1 U560 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1199), .Y(n305) );
  MUX2X1 U561 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1199), .Y(n304) );
  MUX2X1 U562 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1199), .Y(n308) );
  MUX2X1 U563 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1199), .Y(n307) );
  MUX2X1 U564 ( .B(n306), .A(n303), .S(n1176), .Y(n310) );
  MUX2X1 U565 ( .B(n309), .A(n294), .S(n1170), .Y(n646) );
  MUX2X1 U566 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1199), .Y(n314) );
  MUX2X1 U567 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1199), .Y(n313) );
  MUX2X1 U568 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1199), .Y(n317) );
  MUX2X1 U569 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1199), .Y(n316) );
  MUX2X1 U570 ( .B(n315), .A(n312), .S(n1176), .Y(n326) );
  MUX2X1 U571 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1199), .Y(n320) );
  MUX2X1 U572 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1199), .Y(n319) );
  MUX2X1 U573 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1199), .Y(n323) );
  MUX2X1 U574 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1199), .Y(n322) );
  MUX2X1 U575 ( .B(n321), .A(n318), .S(n1176), .Y(n325) );
  MUX2X1 U576 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1200), .Y(n329) );
  MUX2X1 U577 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1200), .Y(n328) );
  MUX2X1 U578 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1200), .Y(n332) );
  MUX2X1 U579 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1200), .Y(n331) );
  MUX2X1 U580 ( .B(n330), .A(n327), .S(n1176), .Y(n341) );
  MUX2X1 U581 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1200), .Y(n335) );
  MUX2X1 U582 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1200), .Y(n334) );
  MUX2X1 U583 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1200), .Y(n338) );
  MUX2X1 U584 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1200), .Y(n337) );
  MUX2X1 U585 ( .B(n336), .A(n333), .S(n1176), .Y(n340) );
  MUX2X1 U586 ( .B(n339), .A(n324), .S(n1170), .Y(n647) );
  MUX2X1 U587 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1200), .Y(n344) );
  MUX2X1 U588 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1200), .Y(n343) );
  MUX2X1 U589 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1200), .Y(n347) );
  MUX2X1 U590 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1200), .Y(n346) );
  MUX2X1 U591 ( .B(n345), .A(n342), .S(n1177), .Y(n356) );
  MUX2X1 U592 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1201), .Y(n350) );
  MUX2X1 U593 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1201), .Y(n349) );
  MUX2X1 U594 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1201), .Y(n353) );
  MUX2X1 U595 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1201), .Y(n352) );
  MUX2X1 U596 ( .B(n351), .A(n348), .S(n1177), .Y(n355) );
  MUX2X1 U597 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1201), .Y(n359) );
  MUX2X1 U598 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1201), .Y(n358) );
  MUX2X1 U599 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1201), .Y(n362) );
  MUX2X1 U600 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1201), .Y(n361) );
  MUX2X1 U601 ( .B(n360), .A(n357), .S(n1177), .Y(n371) );
  MUX2X1 U602 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1201), .Y(n365) );
  MUX2X1 U603 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1201), .Y(n364) );
  MUX2X1 U604 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1201), .Y(n368) );
  MUX2X1 U605 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1201), .Y(n367) );
  MUX2X1 U606 ( .B(n366), .A(n363), .S(n1177), .Y(n370) );
  MUX2X1 U607 ( .B(n369), .A(n354), .S(n1170), .Y(n648) );
  MUX2X1 U608 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1202), .Y(n374) );
  MUX2X1 U609 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1202), .Y(n373) );
  MUX2X1 U610 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1202), .Y(n377) );
  MUX2X1 U611 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1202), .Y(n376) );
  MUX2X1 U612 ( .B(n375), .A(n372), .S(n1177), .Y(n386) );
  MUX2X1 U613 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1202), .Y(n380) );
  MUX2X1 U614 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1202), .Y(n379) );
  MUX2X1 U615 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1202), .Y(n383) );
  MUX2X1 U616 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1202), .Y(n382) );
  MUX2X1 U617 ( .B(n381), .A(n378), .S(n1177), .Y(n385) );
  MUX2X1 U618 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1202), .Y(n389) );
  MUX2X1 U619 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1202), .Y(n388) );
  MUX2X1 U620 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1202), .Y(n392) );
  MUX2X1 U621 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1202), .Y(n391) );
  MUX2X1 U622 ( .B(n390), .A(n387), .S(n1177), .Y(n401) );
  MUX2X1 U623 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1203), .Y(n395) );
  MUX2X1 U624 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1203), .Y(n394) );
  MUX2X1 U625 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1203), .Y(n398) );
  MUX2X1 U626 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1203), .Y(n397) );
  MUX2X1 U627 ( .B(n396), .A(n393), .S(n1177), .Y(n400) );
  MUX2X1 U628 ( .B(n399), .A(n384), .S(n1170), .Y(n649) );
  MUX2X1 U629 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1203), .Y(n404) );
  MUX2X1 U630 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1203), .Y(n403) );
  MUX2X1 U631 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1203), .Y(n407) );
  MUX2X1 U632 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1203), .Y(n406) );
  MUX2X1 U633 ( .B(n405), .A(n402), .S(n1177), .Y(n416) );
  MUX2X1 U634 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1203), .Y(n410) );
  MUX2X1 U635 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1203), .Y(n409) );
  MUX2X1 U636 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1203), .Y(n413) );
  MUX2X1 U637 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1203), .Y(n412) );
  MUX2X1 U638 ( .B(n411), .A(n408), .S(n1177), .Y(n415) );
  MUX2X1 U639 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1204), .Y(n419) );
  MUX2X1 U640 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1204), .Y(n418) );
  MUX2X1 U641 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1204), .Y(n422) );
  MUX2X1 U642 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1204), .Y(n421) );
  MUX2X1 U643 ( .B(n420), .A(n417), .S(n1177), .Y(n431) );
  MUX2X1 U644 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1204), .Y(n425) );
  MUX2X1 U645 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1204), .Y(n424) );
  MUX2X1 U646 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1204), .Y(n428) );
  MUX2X1 U647 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1204), .Y(n427) );
  MUX2X1 U648 ( .B(n426), .A(n423), .S(n1177), .Y(n430) );
  MUX2X1 U649 ( .B(n429), .A(n414), .S(n1170), .Y(n650) );
  MUX2X1 U650 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1204), .Y(n434) );
  MUX2X1 U651 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1204), .Y(n433) );
  MUX2X1 U652 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1204), .Y(n437) );
  MUX2X1 U653 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1204), .Y(n436) );
  MUX2X1 U654 ( .B(n435), .A(n432), .S(n1175), .Y(n446) );
  MUX2X1 U655 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1205), .Y(n440) );
  MUX2X1 U656 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1205), .Y(n439) );
  MUX2X1 U657 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1205), .Y(n443) );
  MUX2X1 U658 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1205), .Y(n442) );
  MUX2X1 U659 ( .B(n441), .A(n438), .S(n1175), .Y(n445) );
  MUX2X1 U660 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1205), .Y(n449) );
  MUX2X1 U661 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1205), .Y(n448) );
  MUX2X1 U662 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1205), .Y(n452) );
  MUX2X1 U663 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1205), .Y(n451) );
  MUX2X1 U664 ( .B(n450), .A(n447), .S(n1175), .Y(n461) );
  MUX2X1 U665 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1205), .Y(n455) );
  MUX2X1 U666 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1205), .Y(n454) );
  MUX2X1 U667 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1205), .Y(n458) );
  MUX2X1 U668 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1205), .Y(n457) );
  MUX2X1 U669 ( .B(n456), .A(n453), .S(n1175), .Y(n460) );
  MUX2X1 U670 ( .B(n459), .A(n444), .S(n1170), .Y(n1163) );
  MUX2X1 U671 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1205), .Y(n464) );
  MUX2X1 U672 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1207), .Y(n463) );
  MUX2X1 U673 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1317), .Y(n467) );
  MUX2X1 U674 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1317), .Y(n466) );
  MUX2X1 U675 ( .B(n465), .A(n462), .S(n1175), .Y(n476) );
  MUX2X1 U676 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1317), .Y(n470) );
  MUX2X1 U677 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1205), .Y(n469) );
  MUX2X1 U678 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1317), .Y(n473) );
  MUX2X1 U679 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1205), .Y(n472) );
  MUX2X1 U680 ( .B(n471), .A(n468), .S(n1175), .Y(n475) );
  MUX2X1 U681 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1317), .Y(n479) );
  MUX2X1 U682 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1205), .Y(n478) );
  MUX2X1 U683 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1317), .Y(n482) );
  MUX2X1 U684 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1317), .Y(n481) );
  MUX2X1 U685 ( .B(n480), .A(n477), .S(n1175), .Y(n491) );
  MUX2X1 U686 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1201), .Y(n485) );
  MUX2X1 U687 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1201), .Y(n484) );
  MUX2X1 U688 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1203), .Y(n488) );
  MUX2X1 U689 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1201), .Y(n487) );
  MUX2X1 U690 ( .B(n486), .A(n483), .S(n1175), .Y(n490) );
  MUX2X1 U691 ( .B(n489), .A(n474), .S(n1170), .Y(n1164) );
  MUX2X1 U692 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1202), .Y(n494) );
  MUX2X1 U693 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1206), .Y(n493) );
  MUX2X1 U694 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1202), .Y(n497) );
  MUX2X1 U695 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1202), .Y(n496) );
  MUX2X1 U696 ( .B(n495), .A(n492), .S(n1175), .Y(n506) );
  MUX2X1 U697 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1201), .Y(n500) );
  MUX2X1 U698 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1317), .Y(n499) );
  MUX2X1 U699 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1203), .Y(n503) );
  MUX2X1 U700 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1203), .Y(n502) );
  MUX2X1 U701 ( .B(n501), .A(n498), .S(n1175), .Y(n505) );
  MUX2X1 U702 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1206), .Y(n509) );
  MUX2X1 U703 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1206), .Y(n508) );
  MUX2X1 U704 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1206), .Y(n512) );
  MUX2X1 U705 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1206), .Y(n511) );
  MUX2X1 U706 ( .B(n510), .A(n507), .S(n1175), .Y(n521) );
  MUX2X1 U707 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1206), .Y(n515) );
  MUX2X1 U708 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1206), .Y(n514) );
  MUX2X1 U709 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1206), .Y(n518) );
  MUX2X1 U710 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1206), .Y(n517) );
  MUX2X1 U711 ( .B(n516), .A(n513), .S(n1175), .Y(n520) );
  MUX2X1 U712 ( .B(n519), .A(n504), .S(n1170), .Y(n1165) );
  MUX2X1 U713 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1206), .Y(n524) );
  MUX2X1 U714 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1206), .Y(n523) );
  MUX2X1 U715 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1206), .Y(n527) );
  MUX2X1 U716 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1206), .Y(n526) );
  MUX2X1 U717 ( .B(n525), .A(n522), .S(n1174), .Y(n536) );
  MUX2X1 U718 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1207), .Y(n530) );
  MUX2X1 U719 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1207), .Y(n529) );
  MUX2X1 U720 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1207), .Y(n533) );
  MUX2X1 U721 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1207), .Y(n532) );
  MUX2X1 U722 ( .B(n531), .A(n528), .S(n1174), .Y(n535) );
  MUX2X1 U723 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1207), .Y(n539) );
  MUX2X1 U724 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1207), .Y(n538) );
  MUX2X1 U725 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1207), .Y(n542) );
  MUX2X1 U726 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1207), .Y(n541) );
  MUX2X1 U727 ( .B(n540), .A(n537), .S(n1174), .Y(n551) );
  MUX2X1 U728 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1207), .Y(n545) );
  MUX2X1 U729 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1207), .Y(n544) );
  MUX2X1 U730 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1207), .Y(n548) );
  MUX2X1 U731 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1207), .Y(n547) );
  MUX2X1 U732 ( .B(n546), .A(n543), .S(n1174), .Y(n550) );
  MUX2X1 U733 ( .B(n549), .A(n534), .S(n1170), .Y(n1166) );
  MUX2X1 U734 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1208), .Y(n554) );
  MUX2X1 U735 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1208), .Y(n553) );
  MUX2X1 U736 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1208), .Y(n557) );
  MUX2X1 U737 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1208), .Y(n556) );
  MUX2X1 U738 ( .B(n555), .A(n552), .S(n1174), .Y(n566) );
  MUX2X1 U739 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1208), .Y(n560) );
  MUX2X1 U740 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1208), .Y(n559) );
  MUX2X1 U741 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1208), .Y(n563) );
  MUX2X1 U742 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1208), .Y(n562) );
  MUX2X1 U743 ( .B(n561), .A(n558), .S(n1174), .Y(n565) );
  MUX2X1 U744 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1208), .Y(n569) );
  MUX2X1 U745 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1208), .Y(n568) );
  MUX2X1 U746 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1208), .Y(n572) );
  MUX2X1 U747 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1208), .Y(n571) );
  MUX2X1 U748 ( .B(n570), .A(n567), .S(n1174), .Y(n581) );
  MUX2X1 U749 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1207), .Y(n575) );
  MUX2X1 U750 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1207), .Y(n574) );
  MUX2X1 U751 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1207), .Y(n578) );
  MUX2X1 U752 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1207), .Y(n577) );
  MUX2X1 U753 ( .B(n576), .A(n573), .S(n1174), .Y(n580) );
  MUX2X1 U754 ( .B(n579), .A(n564), .S(N14), .Y(n1167) );
  MUX2X1 U755 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1207), .Y(n584) );
  MUX2X1 U756 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1207), .Y(n583) );
  MUX2X1 U757 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1207), .Y(n587) );
  MUX2X1 U758 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1207), .Y(n586) );
  MUX2X1 U759 ( .B(n585), .A(n582), .S(n1174), .Y(n596) );
  MUX2X1 U760 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1207), .Y(n590) );
  MUX2X1 U761 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1207), .Y(n589) );
  MUX2X1 U762 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1207), .Y(n593) );
  MUX2X1 U763 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1207), .Y(n592) );
  MUX2X1 U764 ( .B(n591), .A(n588), .S(n1174), .Y(n595) );
  MUX2X1 U765 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1208), .Y(n599) );
  MUX2X1 U766 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1208), .Y(n598) );
  MUX2X1 U767 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1208), .Y(n602) );
  MUX2X1 U768 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1208), .Y(n601) );
  MUX2X1 U769 ( .B(n600), .A(n597), .S(n1174), .Y(n611) );
  MUX2X1 U770 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1208), .Y(n605) );
  MUX2X1 U771 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1208), .Y(n604) );
  MUX2X1 U772 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1208), .Y(n608) );
  MUX2X1 U773 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1208), .Y(n607) );
  MUX2X1 U774 ( .B(n606), .A(n603), .S(n1174), .Y(n610) );
  MUX2X1 U775 ( .B(n609), .A(n594), .S(N14), .Y(n1168) );
  MUX2X1 U776 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1206), .Y(n614) );
  MUX2X1 U777 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1206), .Y(n613) );
  MUX2X1 U778 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1208), .Y(n617) );
  MUX2X1 U779 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1208), .Y(n616) );
  MUX2X1 U780 ( .B(n615), .A(n612), .S(n1174), .Y(n626) );
  MUX2X1 U781 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1209), .Y(n620) );
  MUX2X1 U782 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1209), .Y(n619) );
  MUX2X1 U783 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1209), .Y(n623) );
  MUX2X1 U784 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1209), .Y(n622) );
  MUX2X1 U785 ( .B(n621), .A(n618), .S(n1176), .Y(n625) );
  MUX2X1 U786 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1209), .Y(n629) );
  MUX2X1 U787 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1209), .Y(n628) );
  MUX2X1 U788 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1209), .Y(n632) );
  MUX2X1 U789 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1209), .Y(n631) );
  MUX2X1 U790 ( .B(n630), .A(n627), .S(n1175), .Y(n641) );
  MUX2X1 U791 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1209), .Y(n635) );
  MUX2X1 U792 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1209), .Y(n634) );
  MUX2X1 U793 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1209), .Y(n638) );
  MUX2X1 U794 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1209), .Y(n637) );
  MUX2X1 U795 ( .B(n636), .A(n633), .S(n1176), .Y(n640) );
  MUX2X1 U796 ( .B(n639), .A(n624), .S(n1170), .Y(n1169) );
  INVX8 U797 ( .A(n1193), .Y(n1195) );
  INVX8 U798 ( .A(n1193), .Y(n1196) );
  INVX8 U799 ( .A(n1193), .Y(n1197) );
  INVX8 U800 ( .A(n1193), .Y(n1208) );
  INVX1 U801 ( .A(N12), .Y(n1322) );
  AND2X2 U802 ( .A(n1), .B(N29), .Y(\data_out<3> ) );
  INVX1 U803 ( .A(N11), .Y(n1320) );
  INVX1 U804 ( .A(N10), .Y(n1318) );
  INVX8 U805 ( .A(n7), .Y(n1284) );
  INVX8 U806 ( .A(n7), .Y(n1285) );
  INVX8 U807 ( .A(n10), .Y(n1286) );
  INVX8 U808 ( .A(n10), .Y(n1287) );
  INVX8 U809 ( .A(n11), .Y(n1288) );
  INVX8 U810 ( .A(n11), .Y(n1289) );
  INVX8 U811 ( .A(n12), .Y(n1290) );
  INVX8 U812 ( .A(n12), .Y(n1291) );
  INVX8 U813 ( .A(n13), .Y(n1292) );
  INVX8 U814 ( .A(n13), .Y(n1293) );
  INVX8 U815 ( .A(n14), .Y(n1294) );
  INVX8 U816 ( .A(n14), .Y(n1295) );
  INVX8 U817 ( .A(n15), .Y(n1296) );
  INVX8 U818 ( .A(n15), .Y(n1297) );
  INVX8 U819 ( .A(n16), .Y(n1298) );
  INVX8 U820 ( .A(n16), .Y(n1299) );
  INVX8 U821 ( .A(n17), .Y(n1300) );
  INVX8 U822 ( .A(n17), .Y(n1301) );
  INVX8 U823 ( .A(n18), .Y(n1302) );
  INVX8 U824 ( .A(n18), .Y(n1303) );
  INVX8 U825 ( .A(n19), .Y(n1304) );
  INVX8 U826 ( .A(n19), .Y(n1305) );
  INVX8 U827 ( .A(n20), .Y(n1306) );
  INVX8 U828 ( .A(n20), .Y(n1307) );
  INVX8 U829 ( .A(n21), .Y(n1308) );
  INVX8 U830 ( .A(n21), .Y(n1309) );
  INVX8 U831 ( .A(n22), .Y(n1310) );
  INVX8 U832 ( .A(n22), .Y(n1311) );
  INVX8 U833 ( .A(n23), .Y(n1312) );
  INVX8 U834 ( .A(n23), .Y(n1313) );
  INVX8 U835 ( .A(n24), .Y(n1314) );
  INVX8 U836 ( .A(n24), .Y(n1315) );
  AND2X2 U837 ( .A(n4), .B(N32), .Y(\data_out<0> ) );
  AND2X2 U838 ( .A(n1), .B(N31), .Y(\data_out<1> ) );
  AND2X2 U839 ( .A(n6), .B(N30), .Y(\data_out<2> ) );
  AND2X2 U840 ( .A(n1), .B(N28), .Y(\data_out<4> ) );
  AND2X2 U841 ( .A(n6), .B(N27), .Y(\data_out<5> ) );
  AND2X2 U842 ( .A(n6), .B(N26), .Y(\data_out<6> ) );
  AND2X2 U843 ( .A(n6), .B(N25), .Y(\data_out<7> ) );
  AND2X2 U844 ( .A(n1), .B(N24), .Y(\data_out<8> ) );
  AND2X2 U845 ( .A(n6), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U846 ( .A(n1), .B(N22), .Y(\data_out<10> ) );
  AND2X2 U847 ( .A(n1), .B(N21), .Y(\data_out<11> ) );
  AND2X2 U848 ( .A(n1), .B(N20), .Y(\data_out<12> ) );
  AND2X2 U849 ( .A(n6), .B(N19), .Y(\data_out<13> ) );
  AND2X2 U850 ( .A(n4), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U851 ( .A(n4), .B(N17), .Y(\data_out<15> ) );
  NAND2X1 U852 ( .A(\mem<31><0> ), .B(n1211), .Y(n1325) );
  OAI21X1 U853 ( .A(n106), .B(n1284), .C(n1325), .Y(n2363) );
  NAND2X1 U854 ( .A(\mem<31><1> ), .B(n1211), .Y(n1326) );
  OAI21X1 U855 ( .A(n1287), .B(n106), .C(n1326), .Y(n2362) );
  NAND2X1 U856 ( .A(\mem<31><2> ), .B(n1211), .Y(n1327) );
  OAI21X1 U857 ( .A(n1289), .B(n106), .C(n1327), .Y(n2361) );
  NAND2X1 U858 ( .A(\mem<31><3> ), .B(n1211), .Y(n1328) );
  OAI21X1 U859 ( .A(n1291), .B(n106), .C(n1328), .Y(n2360) );
  NAND2X1 U860 ( .A(\mem<31><4> ), .B(n1211), .Y(n1329) );
  OAI21X1 U861 ( .A(n1293), .B(n106), .C(n1329), .Y(n2359) );
  NAND2X1 U862 ( .A(\mem<31><5> ), .B(n1211), .Y(n1330) );
  OAI21X1 U863 ( .A(n1295), .B(n106), .C(n1330), .Y(n2358) );
  NAND2X1 U864 ( .A(\mem<31><6> ), .B(n1211), .Y(n1331) );
  OAI21X1 U865 ( .A(n1297), .B(n106), .C(n1331), .Y(n2357) );
  NAND2X1 U866 ( .A(\mem<31><7> ), .B(n1211), .Y(n1332) );
  OAI21X1 U867 ( .A(n1299), .B(n106), .C(n1332), .Y(n2356) );
  NAND2X1 U868 ( .A(\mem<31><8> ), .B(n1212), .Y(n1333) );
  OAI21X1 U869 ( .A(n1301), .B(n106), .C(n1333), .Y(n2355) );
  NAND2X1 U870 ( .A(\mem<31><9> ), .B(n1212), .Y(n1334) );
  OAI21X1 U871 ( .A(n1303), .B(n106), .C(n1334), .Y(n2354) );
  NAND2X1 U872 ( .A(\mem<31><10> ), .B(n1212), .Y(n1335) );
  OAI21X1 U873 ( .A(n1305), .B(n106), .C(n1335), .Y(n2353) );
  NAND2X1 U874 ( .A(\mem<31><11> ), .B(n1212), .Y(n1336) );
  OAI21X1 U875 ( .A(n1307), .B(n106), .C(n1336), .Y(n2352) );
  NAND2X1 U876 ( .A(\mem<31><12> ), .B(n1212), .Y(n1337) );
  OAI21X1 U877 ( .A(n1309), .B(n106), .C(n1337), .Y(n2351) );
  NAND2X1 U878 ( .A(\mem<31><13> ), .B(n1212), .Y(n1338) );
  OAI21X1 U879 ( .A(n1311), .B(n106), .C(n1338), .Y(n2350) );
  NAND2X1 U880 ( .A(\mem<31><14> ), .B(n1212), .Y(n1339) );
  OAI21X1 U881 ( .A(n1313), .B(n106), .C(n1339), .Y(n2349) );
  NAND2X1 U882 ( .A(\mem<31><15> ), .B(n1212), .Y(n1340) );
  OAI21X1 U883 ( .A(n1315), .B(n106), .C(n1340), .Y(n2348) );
  NAND2X1 U884 ( .A(\mem<30><0> ), .B(n1213), .Y(n1341) );
  OAI21X1 U885 ( .A(n108), .B(n1284), .C(n1341), .Y(n2347) );
  NAND2X1 U886 ( .A(\mem<30><1> ), .B(n1213), .Y(n1342) );
  OAI21X1 U887 ( .A(n108), .B(n1287), .C(n1342), .Y(n2346) );
  NAND2X1 U888 ( .A(\mem<30><2> ), .B(n1213), .Y(n1343) );
  OAI21X1 U889 ( .A(n108), .B(n1289), .C(n1343), .Y(n2345) );
  NAND2X1 U890 ( .A(\mem<30><3> ), .B(n1213), .Y(n1344) );
  OAI21X1 U891 ( .A(n108), .B(n1291), .C(n1344), .Y(n2344) );
  NAND2X1 U892 ( .A(\mem<30><4> ), .B(n1213), .Y(n1345) );
  OAI21X1 U893 ( .A(n108), .B(n1293), .C(n1345), .Y(n2343) );
  NAND2X1 U894 ( .A(\mem<30><5> ), .B(n1213), .Y(n1346) );
  OAI21X1 U895 ( .A(n108), .B(n1295), .C(n1346), .Y(n2342) );
  NAND2X1 U896 ( .A(\mem<30><6> ), .B(n1213), .Y(n1347) );
  OAI21X1 U897 ( .A(n108), .B(n1297), .C(n1347), .Y(n2341) );
  NAND2X1 U898 ( .A(\mem<30><7> ), .B(n1213), .Y(n1348) );
  OAI21X1 U899 ( .A(n108), .B(n1299), .C(n1348), .Y(n2340) );
  NAND2X1 U900 ( .A(\mem<30><8> ), .B(n1214), .Y(n1349) );
  OAI21X1 U901 ( .A(n108), .B(n1300), .C(n1349), .Y(n2339) );
  NAND2X1 U902 ( .A(\mem<30><9> ), .B(n1214), .Y(n1350) );
  OAI21X1 U903 ( .A(n108), .B(n1302), .C(n1350), .Y(n2338) );
  NAND2X1 U904 ( .A(\mem<30><10> ), .B(n1214), .Y(n1351) );
  OAI21X1 U905 ( .A(n108), .B(n1304), .C(n1351), .Y(n2337) );
  NAND2X1 U906 ( .A(\mem<30><11> ), .B(n1214), .Y(n1352) );
  OAI21X1 U907 ( .A(n108), .B(n1306), .C(n1352), .Y(n2336) );
  NAND2X1 U908 ( .A(\mem<30><12> ), .B(n1214), .Y(n1353) );
  OAI21X1 U909 ( .A(n108), .B(n1308), .C(n1353), .Y(n2335) );
  NAND2X1 U910 ( .A(\mem<30><13> ), .B(n1214), .Y(n1354) );
  OAI21X1 U911 ( .A(n108), .B(n1310), .C(n1354), .Y(n2334) );
  NAND2X1 U912 ( .A(\mem<30><14> ), .B(n1214), .Y(n1355) );
  OAI21X1 U913 ( .A(n108), .B(n1312), .C(n1355), .Y(n2333) );
  NAND2X1 U914 ( .A(\mem<30><15> ), .B(n1214), .Y(n1356) );
  OAI21X1 U915 ( .A(n108), .B(n1314), .C(n1356), .Y(n2332) );
  NAND3X1 U916 ( .A(n1317), .B(n1321), .C(n1320), .Y(n1357) );
  NAND2X1 U917 ( .A(\mem<29><0> ), .B(n1215), .Y(n1358) );
  OAI21X1 U918 ( .A(n110), .B(n1284), .C(n1358), .Y(n2331) );
  NAND2X1 U919 ( .A(\mem<29><1> ), .B(n1215), .Y(n1359) );
  OAI21X1 U920 ( .A(n110), .B(n1286), .C(n1359), .Y(n2330) );
  NAND2X1 U921 ( .A(\mem<29><2> ), .B(n1215), .Y(n1360) );
  OAI21X1 U922 ( .A(n110), .B(n1288), .C(n1360), .Y(n2329) );
  NAND2X1 U923 ( .A(\mem<29><3> ), .B(n1215), .Y(n1361) );
  OAI21X1 U924 ( .A(n110), .B(n1290), .C(n1361), .Y(n2328) );
  NAND2X1 U925 ( .A(\mem<29><4> ), .B(n1215), .Y(n1362) );
  OAI21X1 U926 ( .A(n110), .B(n1292), .C(n1362), .Y(n2327) );
  NAND2X1 U927 ( .A(\mem<29><5> ), .B(n1215), .Y(n1363) );
  OAI21X1 U928 ( .A(n110), .B(n1294), .C(n1363), .Y(n2326) );
  NAND2X1 U929 ( .A(\mem<29><6> ), .B(n1215), .Y(n1364) );
  OAI21X1 U930 ( .A(n110), .B(n1296), .C(n1364), .Y(n2325) );
  NAND2X1 U931 ( .A(\mem<29><7> ), .B(n1215), .Y(n1365) );
  OAI21X1 U932 ( .A(n110), .B(n1298), .C(n1365), .Y(n2324) );
  NAND2X1 U933 ( .A(\mem<29><8> ), .B(n1216), .Y(n1366) );
  OAI21X1 U934 ( .A(n110), .B(n1301), .C(n1366), .Y(n2323) );
  NAND2X1 U935 ( .A(\mem<29><9> ), .B(n1216), .Y(n1367) );
  OAI21X1 U936 ( .A(n110), .B(n1303), .C(n1367), .Y(n2322) );
  NAND2X1 U937 ( .A(\mem<29><10> ), .B(n1216), .Y(n1368) );
  OAI21X1 U938 ( .A(n110), .B(n1305), .C(n1368), .Y(n2321) );
  NAND2X1 U939 ( .A(\mem<29><11> ), .B(n1216), .Y(n1369) );
  OAI21X1 U940 ( .A(n110), .B(n1307), .C(n1369), .Y(n2320) );
  NAND2X1 U941 ( .A(\mem<29><12> ), .B(n1216), .Y(n1370) );
  OAI21X1 U942 ( .A(n110), .B(n1309), .C(n1370), .Y(n2319) );
  NAND2X1 U943 ( .A(\mem<29><13> ), .B(n1216), .Y(n1371) );
  OAI21X1 U944 ( .A(n110), .B(n1311), .C(n1371), .Y(n2318) );
  NAND2X1 U945 ( .A(\mem<29><14> ), .B(n1216), .Y(n1372) );
  OAI21X1 U946 ( .A(n110), .B(n1313), .C(n1372), .Y(n2317) );
  NAND2X1 U947 ( .A(\mem<29><15> ), .B(n1216), .Y(n1373) );
  OAI21X1 U948 ( .A(n110), .B(n1315), .C(n1373), .Y(n2316) );
  NAND3X1 U949 ( .A(n1321), .B(n1320), .C(n1318), .Y(n1374) );
  NAND2X1 U950 ( .A(\mem<28><0> ), .B(n1217), .Y(n1375) );
  OAI21X1 U951 ( .A(n112), .B(n1284), .C(n1375), .Y(n2315) );
  NAND2X1 U952 ( .A(\mem<28><1> ), .B(n1217), .Y(n1376) );
  OAI21X1 U953 ( .A(n112), .B(n1287), .C(n1376), .Y(n2314) );
  NAND2X1 U954 ( .A(\mem<28><2> ), .B(n1217), .Y(n1377) );
  OAI21X1 U955 ( .A(n112), .B(n1289), .C(n1377), .Y(n2313) );
  NAND2X1 U956 ( .A(\mem<28><3> ), .B(n1217), .Y(n1378) );
  OAI21X1 U957 ( .A(n112), .B(n1291), .C(n1378), .Y(n2312) );
  NAND2X1 U958 ( .A(\mem<28><4> ), .B(n1217), .Y(n1379) );
  OAI21X1 U959 ( .A(n112), .B(n1293), .C(n1379), .Y(n2311) );
  NAND2X1 U960 ( .A(\mem<28><5> ), .B(n1217), .Y(n1380) );
  OAI21X1 U961 ( .A(n112), .B(n1295), .C(n1380), .Y(n2310) );
  NAND2X1 U962 ( .A(\mem<28><6> ), .B(n1217), .Y(n1381) );
  OAI21X1 U963 ( .A(n112), .B(n1297), .C(n1381), .Y(n2309) );
  NAND2X1 U964 ( .A(\mem<28><7> ), .B(n1217), .Y(n1382) );
  OAI21X1 U965 ( .A(n112), .B(n1299), .C(n1382), .Y(n2308) );
  NAND2X1 U966 ( .A(\mem<28><8> ), .B(n1218), .Y(n1383) );
  OAI21X1 U967 ( .A(n112), .B(n1300), .C(n1383), .Y(n2307) );
  NAND2X1 U968 ( .A(\mem<28><9> ), .B(n1218), .Y(n1384) );
  OAI21X1 U969 ( .A(n112), .B(n1302), .C(n1384), .Y(n2306) );
  NAND2X1 U970 ( .A(\mem<28><10> ), .B(n1218), .Y(n1385) );
  OAI21X1 U971 ( .A(n112), .B(n1304), .C(n1385), .Y(n2305) );
  NAND2X1 U972 ( .A(\mem<28><11> ), .B(n1218), .Y(n1386) );
  OAI21X1 U973 ( .A(n112), .B(n1306), .C(n1386), .Y(n2304) );
  NAND2X1 U974 ( .A(\mem<28><12> ), .B(n1218), .Y(n1387) );
  OAI21X1 U975 ( .A(n112), .B(n1308), .C(n1387), .Y(n2303) );
  NAND2X1 U976 ( .A(\mem<28><13> ), .B(n1218), .Y(n1388) );
  OAI21X1 U977 ( .A(n112), .B(n1310), .C(n1388), .Y(n2302) );
  NAND2X1 U978 ( .A(\mem<28><14> ), .B(n1218), .Y(n1389) );
  OAI21X1 U979 ( .A(n112), .B(n1312), .C(n1389), .Y(n2301) );
  NAND2X1 U980 ( .A(\mem<28><15> ), .B(n1218), .Y(n1390) );
  OAI21X1 U981 ( .A(n112), .B(n1314), .C(n1390), .Y(n2300) );
  NAND3X1 U982 ( .A(n1317), .B(n1319), .C(n1322), .Y(n1391) );
  NAND2X1 U983 ( .A(\mem<27><0> ), .B(n1219), .Y(n1392) );
  OAI21X1 U984 ( .A(n114), .B(n1284), .C(n1392), .Y(n2299) );
  NAND2X1 U985 ( .A(\mem<27><1> ), .B(n1219), .Y(n1393) );
  OAI21X1 U986 ( .A(n114), .B(n1286), .C(n1393), .Y(n2298) );
  NAND2X1 U987 ( .A(\mem<27><2> ), .B(n1219), .Y(n1394) );
  OAI21X1 U988 ( .A(n114), .B(n1288), .C(n1394), .Y(n2297) );
  NAND2X1 U989 ( .A(\mem<27><3> ), .B(n1219), .Y(n1395) );
  OAI21X1 U990 ( .A(n114), .B(n1290), .C(n1395), .Y(n2296) );
  NAND2X1 U991 ( .A(\mem<27><4> ), .B(n1219), .Y(n1396) );
  OAI21X1 U992 ( .A(n114), .B(n1292), .C(n1396), .Y(n2295) );
  NAND2X1 U993 ( .A(\mem<27><5> ), .B(n1219), .Y(n1397) );
  OAI21X1 U994 ( .A(n114), .B(n1294), .C(n1397), .Y(n2294) );
  NAND2X1 U995 ( .A(\mem<27><6> ), .B(n1219), .Y(n1398) );
  OAI21X1 U996 ( .A(n114), .B(n1296), .C(n1398), .Y(n2293) );
  NAND2X1 U997 ( .A(\mem<27><7> ), .B(n1219), .Y(n1399) );
  OAI21X1 U998 ( .A(n114), .B(n1298), .C(n1399), .Y(n2292) );
  NAND2X1 U999 ( .A(\mem<27><8> ), .B(n1220), .Y(n1400) );
  OAI21X1 U1000 ( .A(n114), .B(n1301), .C(n1400), .Y(n2291) );
  NAND2X1 U1001 ( .A(\mem<27><9> ), .B(n1220), .Y(n1401) );
  OAI21X1 U1002 ( .A(n114), .B(n1303), .C(n1401), .Y(n2290) );
  NAND2X1 U1003 ( .A(\mem<27><10> ), .B(n1220), .Y(n1402) );
  OAI21X1 U1004 ( .A(n114), .B(n1305), .C(n1402), .Y(n2289) );
  NAND2X1 U1005 ( .A(\mem<27><11> ), .B(n1220), .Y(n1403) );
  OAI21X1 U1006 ( .A(n114), .B(n1307), .C(n1403), .Y(n2288) );
  NAND2X1 U1007 ( .A(\mem<27><12> ), .B(n1220), .Y(n1404) );
  OAI21X1 U1008 ( .A(n114), .B(n1309), .C(n1404), .Y(n2287) );
  NAND2X1 U1009 ( .A(\mem<27><13> ), .B(n1220), .Y(n1405) );
  OAI21X1 U1010 ( .A(n114), .B(n1311), .C(n1405), .Y(n2286) );
  NAND2X1 U1011 ( .A(\mem<27><14> ), .B(n1220), .Y(n1406) );
  OAI21X1 U1012 ( .A(n114), .B(n1313), .C(n1406), .Y(n2285) );
  NAND2X1 U1013 ( .A(\mem<27><15> ), .B(n1220), .Y(n1407) );
  OAI21X1 U1014 ( .A(n114), .B(n1315), .C(n1407), .Y(n2284) );
  NAND3X1 U1015 ( .A(n1322), .B(n1319), .C(n1318), .Y(n1408) );
  NAND2X1 U1016 ( .A(\mem<26><0> ), .B(n1221), .Y(n1409) );
  OAI21X1 U1017 ( .A(n116), .B(n1284), .C(n1409), .Y(n2283) );
  NAND2X1 U1018 ( .A(\mem<26><1> ), .B(n1221), .Y(n1410) );
  OAI21X1 U1019 ( .A(n116), .B(n1287), .C(n1410), .Y(n2282) );
  NAND2X1 U1020 ( .A(\mem<26><2> ), .B(n1221), .Y(n1411) );
  OAI21X1 U1021 ( .A(n116), .B(n1289), .C(n1411), .Y(n2281) );
  NAND2X1 U1022 ( .A(\mem<26><3> ), .B(n1221), .Y(n1412) );
  OAI21X1 U1023 ( .A(n116), .B(n1291), .C(n1412), .Y(n2280) );
  NAND2X1 U1024 ( .A(\mem<26><4> ), .B(n1221), .Y(n1413) );
  OAI21X1 U1025 ( .A(n116), .B(n1293), .C(n1413), .Y(n2279) );
  NAND2X1 U1026 ( .A(\mem<26><5> ), .B(n1221), .Y(n1414) );
  OAI21X1 U1027 ( .A(n116), .B(n1295), .C(n1414), .Y(n2278) );
  NAND2X1 U1028 ( .A(\mem<26><6> ), .B(n1221), .Y(n1415) );
  OAI21X1 U1029 ( .A(n116), .B(n1297), .C(n1415), .Y(n2277) );
  NAND2X1 U1030 ( .A(\mem<26><7> ), .B(n1221), .Y(n1416) );
  OAI21X1 U1031 ( .A(n116), .B(n1299), .C(n1416), .Y(n2276) );
  NAND2X1 U1032 ( .A(\mem<26><8> ), .B(n1222), .Y(n1417) );
  OAI21X1 U1033 ( .A(n116), .B(n1300), .C(n1417), .Y(n2275) );
  NAND2X1 U1034 ( .A(\mem<26><9> ), .B(n1222), .Y(n1418) );
  OAI21X1 U1035 ( .A(n116), .B(n1302), .C(n1418), .Y(n2274) );
  NAND2X1 U1036 ( .A(\mem<26><10> ), .B(n1222), .Y(n1419) );
  OAI21X1 U1037 ( .A(n116), .B(n1304), .C(n1419), .Y(n2273) );
  NAND2X1 U1038 ( .A(\mem<26><11> ), .B(n1222), .Y(n1420) );
  OAI21X1 U1039 ( .A(n116), .B(n1306), .C(n1420), .Y(n2272) );
  NAND2X1 U1040 ( .A(\mem<26><12> ), .B(n1222), .Y(n1421) );
  OAI21X1 U1041 ( .A(n116), .B(n1308), .C(n1421), .Y(n2271) );
  NAND2X1 U1042 ( .A(\mem<26><13> ), .B(n1222), .Y(n1422) );
  OAI21X1 U1043 ( .A(n116), .B(n1310), .C(n1422), .Y(n2270) );
  NAND2X1 U1044 ( .A(\mem<26><14> ), .B(n1222), .Y(n1423) );
  OAI21X1 U1045 ( .A(n116), .B(n1312), .C(n1423), .Y(n2269) );
  NAND2X1 U1046 ( .A(\mem<26><15> ), .B(n1222), .Y(n1424) );
  OAI21X1 U1047 ( .A(n116), .B(n1314), .C(n1424), .Y(n2268) );
  NAND3X1 U1048 ( .A(n1317), .B(n1322), .C(n1320), .Y(n1425) );
  NAND2X1 U1049 ( .A(\mem<25><0> ), .B(n1223), .Y(n1426) );
  OAI21X1 U1050 ( .A(n118), .B(n1284), .C(n1426), .Y(n2267) );
  NAND2X1 U1051 ( .A(\mem<25><1> ), .B(n1223), .Y(n1427) );
  OAI21X1 U1052 ( .A(n118), .B(n1286), .C(n1427), .Y(n2266) );
  NAND2X1 U1053 ( .A(\mem<25><2> ), .B(n1223), .Y(n1428) );
  OAI21X1 U1054 ( .A(n118), .B(n1288), .C(n1428), .Y(n2265) );
  NAND2X1 U1055 ( .A(\mem<25><3> ), .B(n1223), .Y(n1429) );
  OAI21X1 U1056 ( .A(n118), .B(n1290), .C(n1429), .Y(n2264) );
  NAND2X1 U1057 ( .A(\mem<25><4> ), .B(n1223), .Y(n1430) );
  OAI21X1 U1058 ( .A(n118), .B(n1292), .C(n1430), .Y(n2263) );
  NAND2X1 U1059 ( .A(\mem<25><5> ), .B(n1223), .Y(n1431) );
  OAI21X1 U1060 ( .A(n118), .B(n1294), .C(n1431), .Y(n2262) );
  NAND2X1 U1061 ( .A(\mem<25><6> ), .B(n1223), .Y(n1432) );
  OAI21X1 U1062 ( .A(n118), .B(n1296), .C(n1432), .Y(n2261) );
  NAND2X1 U1063 ( .A(\mem<25><7> ), .B(n1223), .Y(n1433) );
  OAI21X1 U1064 ( .A(n118), .B(n1298), .C(n1433), .Y(n2260) );
  NAND2X1 U1065 ( .A(\mem<25><8> ), .B(n1224), .Y(n1434) );
  OAI21X1 U1066 ( .A(n118), .B(n1301), .C(n1434), .Y(n2259) );
  NAND2X1 U1067 ( .A(\mem<25><9> ), .B(n1224), .Y(n1435) );
  OAI21X1 U1068 ( .A(n118), .B(n1303), .C(n1435), .Y(n2258) );
  NAND2X1 U1069 ( .A(\mem<25><10> ), .B(n1224), .Y(n1436) );
  OAI21X1 U1070 ( .A(n118), .B(n1305), .C(n1436), .Y(n2257) );
  NAND2X1 U1071 ( .A(\mem<25><11> ), .B(n1224), .Y(n1437) );
  OAI21X1 U1072 ( .A(n118), .B(n1307), .C(n1437), .Y(n2256) );
  NAND2X1 U1073 ( .A(\mem<25><12> ), .B(n1224), .Y(n1438) );
  OAI21X1 U1074 ( .A(n118), .B(n1309), .C(n1438), .Y(n2255) );
  NAND2X1 U1075 ( .A(\mem<25><13> ), .B(n1224), .Y(n1439) );
  OAI21X1 U1076 ( .A(n118), .B(n1311), .C(n1439), .Y(n2254) );
  NAND2X1 U1077 ( .A(\mem<25><14> ), .B(n1224), .Y(n1440) );
  OAI21X1 U1078 ( .A(n118), .B(n1313), .C(n1440), .Y(n2253) );
  NAND2X1 U1079 ( .A(\mem<25><15> ), .B(n1224), .Y(n1441) );
  OAI21X1 U1080 ( .A(n118), .B(n1315), .C(n1441), .Y(n2252) );
  NOR3X1 U1081 ( .A(n1317), .B(n1319), .C(n1321), .Y(n1835) );
  NAND2X1 U1082 ( .A(\mem<24><0> ), .B(n1226), .Y(n1442) );
  OAI21X1 U1083 ( .A(n1225), .B(n1284), .C(n1442), .Y(n2251) );
  NAND2X1 U1084 ( .A(\mem<24><1> ), .B(n1226), .Y(n1443) );
  OAI21X1 U1085 ( .A(n1225), .B(n1286), .C(n1443), .Y(n2250) );
  NAND2X1 U1086 ( .A(\mem<24><2> ), .B(n1226), .Y(n1444) );
  OAI21X1 U1087 ( .A(n1225), .B(n1288), .C(n1444), .Y(n2249) );
  NAND2X1 U1088 ( .A(\mem<24><3> ), .B(n1226), .Y(n1445) );
  OAI21X1 U1089 ( .A(n1225), .B(n1290), .C(n1445), .Y(n2248) );
  NAND2X1 U1090 ( .A(\mem<24><4> ), .B(n1226), .Y(n1446) );
  OAI21X1 U1091 ( .A(n1225), .B(n1292), .C(n1446), .Y(n2247) );
  NAND2X1 U1092 ( .A(\mem<24><5> ), .B(n1226), .Y(n1447) );
  OAI21X1 U1093 ( .A(n1225), .B(n1294), .C(n1447), .Y(n2246) );
  NAND2X1 U1094 ( .A(\mem<24><6> ), .B(n1226), .Y(n1448) );
  OAI21X1 U1095 ( .A(n1225), .B(n1296), .C(n1448), .Y(n2245) );
  NAND2X1 U1096 ( .A(\mem<24><7> ), .B(n1226), .Y(n1449) );
  OAI21X1 U1097 ( .A(n1225), .B(n1298), .C(n1449), .Y(n2244) );
  NAND2X1 U1098 ( .A(\mem<24><8> ), .B(n1227), .Y(n1450) );
  OAI21X1 U1099 ( .A(n1225), .B(n1300), .C(n1450), .Y(n2243) );
  NAND2X1 U1100 ( .A(\mem<24><9> ), .B(n1227), .Y(n1451) );
  OAI21X1 U1101 ( .A(n1225), .B(n1302), .C(n1451), .Y(n2242) );
  NAND2X1 U1102 ( .A(\mem<24><10> ), .B(n1227), .Y(n1452) );
  OAI21X1 U1103 ( .A(n1225), .B(n1304), .C(n1452), .Y(n2241) );
  NAND2X1 U1104 ( .A(\mem<24><11> ), .B(n1227), .Y(n1453) );
  OAI21X1 U1105 ( .A(n1225), .B(n1306), .C(n1453), .Y(n2240) );
  NAND2X1 U1106 ( .A(\mem<24><12> ), .B(n1227), .Y(n1454) );
  OAI21X1 U1107 ( .A(n1225), .B(n1308), .C(n1454), .Y(n2239) );
  NAND2X1 U1108 ( .A(\mem<24><13> ), .B(n1227), .Y(n1455) );
  OAI21X1 U1109 ( .A(n1225), .B(n1310), .C(n1455), .Y(n2238) );
  NAND2X1 U1110 ( .A(\mem<24><14> ), .B(n1227), .Y(n1456) );
  OAI21X1 U1111 ( .A(n1225), .B(n1312), .C(n1456), .Y(n2237) );
  NAND2X1 U1112 ( .A(\mem<24><15> ), .B(n1227), .Y(n1457) );
  OAI21X1 U1113 ( .A(n1225), .B(n1314), .C(n1457), .Y(n2236) );
  NAND2X1 U1114 ( .A(\mem<23><0> ), .B(n1228), .Y(n1458) );
  OAI21X1 U1115 ( .A(n120), .B(n1284), .C(n1458), .Y(n2235) );
  NAND2X1 U1116 ( .A(\mem<23><1> ), .B(n1228), .Y(n1459) );
  OAI21X1 U1117 ( .A(n120), .B(n1287), .C(n1459), .Y(n2234) );
  NAND2X1 U1118 ( .A(\mem<23><2> ), .B(n1228), .Y(n1460) );
  OAI21X1 U1119 ( .A(n120), .B(n1289), .C(n1460), .Y(n2233) );
  NAND2X1 U1120 ( .A(\mem<23><3> ), .B(n1228), .Y(n1461) );
  OAI21X1 U1121 ( .A(n120), .B(n1291), .C(n1461), .Y(n2232) );
  NAND2X1 U1122 ( .A(\mem<23><4> ), .B(n1228), .Y(n1462) );
  OAI21X1 U1123 ( .A(n120), .B(n1293), .C(n1462), .Y(n2231) );
  NAND2X1 U1124 ( .A(\mem<23><5> ), .B(n1228), .Y(n1463) );
  OAI21X1 U1125 ( .A(n120), .B(n1295), .C(n1463), .Y(n2230) );
  NAND2X1 U1126 ( .A(\mem<23><6> ), .B(n1228), .Y(n1464) );
  OAI21X1 U1127 ( .A(n120), .B(n1297), .C(n1464), .Y(n2229) );
  NAND2X1 U1128 ( .A(\mem<23><7> ), .B(n1228), .Y(n1465) );
  OAI21X1 U1129 ( .A(n120), .B(n1299), .C(n1465), .Y(n2228) );
  NAND2X1 U1130 ( .A(\mem<23><8> ), .B(n1229), .Y(n1466) );
  OAI21X1 U1131 ( .A(n120), .B(n1301), .C(n1466), .Y(n2227) );
  NAND2X1 U1132 ( .A(\mem<23><9> ), .B(n1229), .Y(n1467) );
  OAI21X1 U1133 ( .A(n120), .B(n1303), .C(n1467), .Y(n2226) );
  NAND2X1 U1134 ( .A(\mem<23><10> ), .B(n1229), .Y(n1468) );
  OAI21X1 U1135 ( .A(n120), .B(n1305), .C(n1468), .Y(n2225) );
  NAND2X1 U1136 ( .A(\mem<23><11> ), .B(n1229), .Y(n1469) );
  OAI21X1 U1137 ( .A(n120), .B(n1307), .C(n1469), .Y(n2224) );
  NAND2X1 U1138 ( .A(\mem<23><12> ), .B(n1229), .Y(n1470) );
  OAI21X1 U1139 ( .A(n120), .B(n1309), .C(n1470), .Y(n2223) );
  NAND2X1 U1140 ( .A(\mem<23><13> ), .B(n1229), .Y(n1471) );
  OAI21X1 U1141 ( .A(n120), .B(n1311), .C(n1471), .Y(n2222) );
  NAND2X1 U1142 ( .A(\mem<23><14> ), .B(n1229), .Y(n1472) );
  OAI21X1 U1143 ( .A(n120), .B(n1313), .C(n1472), .Y(n2221) );
  NAND2X1 U1144 ( .A(\mem<23><15> ), .B(n1229), .Y(n1473) );
  OAI21X1 U1145 ( .A(n120), .B(n1315), .C(n1473), .Y(n2220) );
  NAND2X1 U1146 ( .A(\mem<22><0> ), .B(n1230), .Y(n1474) );
  OAI21X1 U1147 ( .A(n122), .B(n1284), .C(n1474), .Y(n2219) );
  NAND2X1 U1148 ( .A(\mem<22><1> ), .B(n1230), .Y(n1475) );
  OAI21X1 U1149 ( .A(n122), .B(n1287), .C(n1475), .Y(n2218) );
  NAND2X1 U1150 ( .A(\mem<22><2> ), .B(n1230), .Y(n1476) );
  OAI21X1 U1151 ( .A(n122), .B(n1289), .C(n1476), .Y(n2217) );
  NAND2X1 U1152 ( .A(\mem<22><3> ), .B(n1230), .Y(n1477) );
  OAI21X1 U1153 ( .A(n122), .B(n1291), .C(n1477), .Y(n2216) );
  NAND2X1 U1154 ( .A(\mem<22><4> ), .B(n1230), .Y(n1478) );
  OAI21X1 U1155 ( .A(n122), .B(n1293), .C(n1478), .Y(n2215) );
  NAND2X1 U1156 ( .A(\mem<22><5> ), .B(n1230), .Y(n1479) );
  OAI21X1 U1157 ( .A(n122), .B(n1295), .C(n1479), .Y(n2214) );
  NAND2X1 U1158 ( .A(\mem<22><6> ), .B(n1230), .Y(n1480) );
  OAI21X1 U1159 ( .A(n122), .B(n1297), .C(n1480), .Y(n2213) );
  NAND2X1 U1160 ( .A(\mem<22><7> ), .B(n1230), .Y(n1481) );
  OAI21X1 U1161 ( .A(n122), .B(n1299), .C(n1481), .Y(n2212) );
  NAND2X1 U1162 ( .A(\mem<22><8> ), .B(n1231), .Y(n1482) );
  OAI21X1 U1163 ( .A(n122), .B(n1301), .C(n1482), .Y(n2211) );
  NAND2X1 U1164 ( .A(\mem<22><9> ), .B(n1231), .Y(n1483) );
  OAI21X1 U1165 ( .A(n122), .B(n1303), .C(n1483), .Y(n2210) );
  NAND2X1 U1166 ( .A(\mem<22><10> ), .B(n1231), .Y(n1484) );
  OAI21X1 U1167 ( .A(n122), .B(n1305), .C(n1484), .Y(n2209) );
  NAND2X1 U1168 ( .A(\mem<22><11> ), .B(n1231), .Y(n1485) );
  OAI21X1 U1169 ( .A(n122), .B(n1307), .C(n1485), .Y(n2208) );
  NAND2X1 U1170 ( .A(\mem<22><12> ), .B(n1231), .Y(n1486) );
  OAI21X1 U1171 ( .A(n122), .B(n1309), .C(n1486), .Y(n2207) );
  NAND2X1 U1172 ( .A(\mem<22><13> ), .B(n1231), .Y(n1487) );
  OAI21X1 U1173 ( .A(n122), .B(n1311), .C(n1487), .Y(n2206) );
  NAND2X1 U1174 ( .A(\mem<22><14> ), .B(n1231), .Y(n1488) );
  OAI21X1 U1175 ( .A(n122), .B(n1313), .C(n1488), .Y(n2205) );
  NAND2X1 U1177 ( .A(\mem<22><15> ), .B(n1231), .Y(n1489) );
  OAI21X1 U1178 ( .A(n122), .B(n1315), .C(n1489), .Y(n2204) );
  NAND2X1 U1179 ( .A(\mem<21><0> ), .B(n1232), .Y(n1490) );
  OAI21X1 U1180 ( .A(n124), .B(n1284), .C(n1490), .Y(n2203) );
  NAND2X1 U1181 ( .A(\mem<21><1> ), .B(n1232), .Y(n1491) );
  OAI21X1 U1182 ( .A(n124), .B(n1287), .C(n1491), .Y(n2202) );
  NAND2X1 U1183 ( .A(\mem<21><2> ), .B(n1232), .Y(n1492) );
  OAI21X1 U1184 ( .A(n124), .B(n1289), .C(n1492), .Y(n2201) );
  NAND2X1 U1185 ( .A(\mem<21><3> ), .B(n1232), .Y(n1493) );
  OAI21X1 U1186 ( .A(n124), .B(n1291), .C(n1493), .Y(n2200) );
  NAND2X1 U1187 ( .A(\mem<21><4> ), .B(n1232), .Y(n1494) );
  OAI21X1 U1188 ( .A(n124), .B(n1293), .C(n1494), .Y(n2199) );
  NAND2X1 U1189 ( .A(\mem<21><5> ), .B(n1232), .Y(n1495) );
  OAI21X1 U1190 ( .A(n124), .B(n1295), .C(n1495), .Y(n2198) );
  NAND2X1 U1191 ( .A(\mem<21><6> ), .B(n1232), .Y(n1496) );
  OAI21X1 U1192 ( .A(n124), .B(n1297), .C(n1496), .Y(n2197) );
  NAND2X1 U1193 ( .A(\mem<21><7> ), .B(n1232), .Y(n1497) );
  OAI21X1 U1194 ( .A(n124), .B(n1299), .C(n1497), .Y(n2196) );
  NAND2X1 U1195 ( .A(\mem<21><8> ), .B(n1233), .Y(n1498) );
  OAI21X1 U1196 ( .A(n124), .B(n1301), .C(n1498), .Y(n2195) );
  NAND2X1 U1197 ( .A(\mem<21><9> ), .B(n1233), .Y(n1499) );
  OAI21X1 U1198 ( .A(n124), .B(n1303), .C(n1499), .Y(n2194) );
  NAND2X1 U1199 ( .A(\mem<21><10> ), .B(n1233), .Y(n1500) );
  OAI21X1 U1200 ( .A(n124), .B(n1305), .C(n1500), .Y(n2193) );
  NAND2X1 U1201 ( .A(\mem<21><11> ), .B(n1233), .Y(n1501) );
  OAI21X1 U1202 ( .A(n124), .B(n1307), .C(n1501), .Y(n2192) );
  NAND2X1 U1203 ( .A(\mem<21><12> ), .B(n1233), .Y(n1502) );
  OAI21X1 U1204 ( .A(n124), .B(n1309), .C(n1502), .Y(n2191) );
  NAND2X1 U1205 ( .A(\mem<21><13> ), .B(n1233), .Y(n1503) );
  OAI21X1 U1206 ( .A(n124), .B(n1311), .C(n1503), .Y(n2190) );
  NAND2X1 U1207 ( .A(\mem<21><14> ), .B(n1233), .Y(n1504) );
  OAI21X1 U1208 ( .A(n124), .B(n1313), .C(n1504), .Y(n2189) );
  NAND2X1 U1209 ( .A(\mem<21><15> ), .B(n1233), .Y(n1505) );
  OAI21X1 U1210 ( .A(n124), .B(n1315), .C(n1505), .Y(n2188) );
  NAND2X1 U1211 ( .A(\mem<20><0> ), .B(n1234), .Y(n1506) );
  OAI21X1 U1212 ( .A(n126), .B(n1284), .C(n1506), .Y(n2187) );
  NAND2X1 U1213 ( .A(\mem<20><1> ), .B(n1234), .Y(n1507) );
  OAI21X1 U1214 ( .A(n126), .B(n1287), .C(n1507), .Y(n2186) );
  NAND2X1 U1215 ( .A(\mem<20><2> ), .B(n1234), .Y(n1508) );
  OAI21X1 U1216 ( .A(n126), .B(n1289), .C(n1508), .Y(n2185) );
  NAND2X1 U1217 ( .A(\mem<20><3> ), .B(n1234), .Y(n1509) );
  OAI21X1 U1218 ( .A(n126), .B(n1291), .C(n1509), .Y(n2184) );
  NAND2X1 U1219 ( .A(\mem<20><4> ), .B(n1234), .Y(n1510) );
  OAI21X1 U1220 ( .A(n126), .B(n1293), .C(n1510), .Y(n2183) );
  NAND2X1 U1221 ( .A(\mem<20><5> ), .B(n1234), .Y(n1511) );
  OAI21X1 U1222 ( .A(n126), .B(n1295), .C(n1511), .Y(n2182) );
  NAND2X1 U1223 ( .A(\mem<20><6> ), .B(n1234), .Y(n1512) );
  OAI21X1 U1224 ( .A(n126), .B(n1297), .C(n1512), .Y(n2181) );
  NAND2X1 U1225 ( .A(\mem<20><7> ), .B(n1234), .Y(n1513) );
  OAI21X1 U1226 ( .A(n126), .B(n1299), .C(n1513), .Y(n2180) );
  NAND2X1 U1227 ( .A(\mem<20><8> ), .B(n1235), .Y(n1514) );
  OAI21X1 U1228 ( .A(n126), .B(n1301), .C(n1514), .Y(n2179) );
  NAND2X1 U1229 ( .A(\mem<20><9> ), .B(n1235), .Y(n1515) );
  OAI21X1 U1230 ( .A(n126), .B(n1303), .C(n1515), .Y(n2178) );
  NAND2X1 U1231 ( .A(\mem<20><10> ), .B(n1235), .Y(n1516) );
  OAI21X1 U1232 ( .A(n126), .B(n1305), .C(n1516), .Y(n2177) );
  NAND2X1 U1233 ( .A(\mem<20><11> ), .B(n1235), .Y(n1517) );
  OAI21X1 U1234 ( .A(n126), .B(n1307), .C(n1517), .Y(n2176) );
  NAND2X1 U1235 ( .A(\mem<20><12> ), .B(n1235), .Y(n1518) );
  OAI21X1 U1236 ( .A(n126), .B(n1309), .C(n1518), .Y(n2175) );
  NAND2X1 U1237 ( .A(\mem<20><13> ), .B(n1235), .Y(n1519) );
  OAI21X1 U1238 ( .A(n126), .B(n1311), .C(n1519), .Y(n2174) );
  NAND2X1 U1239 ( .A(\mem<20><14> ), .B(n1235), .Y(n1520) );
  OAI21X1 U1240 ( .A(n126), .B(n1313), .C(n1520), .Y(n2173) );
  NAND2X1 U1241 ( .A(\mem<20><15> ), .B(n1235), .Y(n1521) );
  OAI21X1 U1242 ( .A(n126), .B(n1315), .C(n1521), .Y(n2172) );
  NAND2X1 U1243 ( .A(\mem<19><0> ), .B(n1236), .Y(n1522) );
  OAI21X1 U1244 ( .A(n128), .B(n1285), .C(n1522), .Y(n2171) );
  NAND2X1 U1245 ( .A(\mem<19><1> ), .B(n1236), .Y(n1523) );
  OAI21X1 U1246 ( .A(n128), .B(n1287), .C(n1523), .Y(n2170) );
  NAND2X1 U1247 ( .A(\mem<19><2> ), .B(n1236), .Y(n1524) );
  OAI21X1 U1248 ( .A(n128), .B(n1289), .C(n1524), .Y(n2169) );
  NAND2X1 U1249 ( .A(\mem<19><3> ), .B(n1236), .Y(n1525) );
  OAI21X1 U1250 ( .A(n128), .B(n1291), .C(n1525), .Y(n2168) );
  NAND2X1 U1251 ( .A(\mem<19><4> ), .B(n1236), .Y(n1526) );
  OAI21X1 U1252 ( .A(n128), .B(n1293), .C(n1526), .Y(n2167) );
  NAND2X1 U1253 ( .A(\mem<19><5> ), .B(n1236), .Y(n1527) );
  OAI21X1 U1254 ( .A(n128), .B(n1295), .C(n1527), .Y(n2166) );
  NAND2X1 U1255 ( .A(\mem<19><6> ), .B(n1236), .Y(n1528) );
  OAI21X1 U1256 ( .A(n128), .B(n1297), .C(n1528), .Y(n2165) );
  NAND2X1 U1257 ( .A(\mem<19><7> ), .B(n1236), .Y(n1529) );
  OAI21X1 U1258 ( .A(n128), .B(n1299), .C(n1529), .Y(n2164) );
  NAND2X1 U1259 ( .A(\mem<19><8> ), .B(n1237), .Y(n1530) );
  OAI21X1 U1260 ( .A(n128), .B(n1301), .C(n1530), .Y(n2163) );
  NAND2X1 U1261 ( .A(\mem<19><9> ), .B(n1237), .Y(n1531) );
  OAI21X1 U1262 ( .A(n128), .B(n1303), .C(n1531), .Y(n2162) );
  NAND2X1 U1263 ( .A(\mem<19><10> ), .B(n1237), .Y(n1532) );
  OAI21X1 U1264 ( .A(n128), .B(n1305), .C(n1532), .Y(n2161) );
  NAND2X1 U1265 ( .A(\mem<19><11> ), .B(n1237), .Y(n1533) );
  OAI21X1 U1266 ( .A(n128), .B(n1307), .C(n1533), .Y(n2160) );
  NAND2X1 U1267 ( .A(\mem<19><12> ), .B(n1237), .Y(n1534) );
  OAI21X1 U1268 ( .A(n128), .B(n1309), .C(n1534), .Y(n2159) );
  NAND2X1 U1269 ( .A(\mem<19><13> ), .B(n1237), .Y(n1535) );
  OAI21X1 U1270 ( .A(n128), .B(n1311), .C(n1535), .Y(n2158) );
  NAND2X1 U1271 ( .A(\mem<19><14> ), .B(n1237), .Y(n1536) );
  OAI21X1 U1272 ( .A(n128), .B(n1313), .C(n1536), .Y(n2157) );
  NAND2X1 U1273 ( .A(\mem<19><15> ), .B(n1237), .Y(n1537) );
  OAI21X1 U1274 ( .A(n128), .B(n1315), .C(n1537), .Y(n2156) );
  NAND2X1 U1275 ( .A(\mem<18><0> ), .B(n1238), .Y(n1538) );
  OAI21X1 U1276 ( .A(n130), .B(n1285), .C(n1538), .Y(n2155) );
  NAND2X1 U1277 ( .A(\mem<18><1> ), .B(n1238), .Y(n1539) );
  OAI21X1 U1278 ( .A(n130), .B(n1287), .C(n1539), .Y(n2154) );
  NAND2X1 U1279 ( .A(\mem<18><2> ), .B(n1238), .Y(n1540) );
  OAI21X1 U1280 ( .A(n130), .B(n1289), .C(n1540), .Y(n2153) );
  NAND2X1 U1281 ( .A(\mem<18><3> ), .B(n1238), .Y(n1541) );
  OAI21X1 U1282 ( .A(n130), .B(n1291), .C(n1541), .Y(n2152) );
  NAND2X1 U1283 ( .A(\mem<18><4> ), .B(n1238), .Y(n1542) );
  OAI21X1 U1284 ( .A(n130), .B(n1293), .C(n1542), .Y(n2151) );
  NAND2X1 U1285 ( .A(\mem<18><5> ), .B(n1238), .Y(n1543) );
  OAI21X1 U1286 ( .A(n130), .B(n1295), .C(n1543), .Y(n2150) );
  NAND2X1 U1287 ( .A(\mem<18><6> ), .B(n1238), .Y(n1544) );
  OAI21X1 U1288 ( .A(n130), .B(n1297), .C(n1544), .Y(n2149) );
  NAND2X1 U1289 ( .A(\mem<18><7> ), .B(n1238), .Y(n1545) );
  OAI21X1 U1290 ( .A(n130), .B(n1299), .C(n1545), .Y(n2148) );
  NAND2X1 U1291 ( .A(\mem<18><8> ), .B(n1239), .Y(n1546) );
  OAI21X1 U1292 ( .A(n130), .B(n1301), .C(n1546), .Y(n2147) );
  NAND2X1 U1293 ( .A(\mem<18><9> ), .B(n1239), .Y(n1547) );
  OAI21X1 U1294 ( .A(n130), .B(n1303), .C(n1547), .Y(n2146) );
  NAND2X1 U1295 ( .A(\mem<18><10> ), .B(n1239), .Y(n1548) );
  OAI21X1 U1296 ( .A(n130), .B(n1305), .C(n1548), .Y(n2145) );
  NAND2X1 U1297 ( .A(\mem<18><11> ), .B(n1239), .Y(n1549) );
  OAI21X1 U1298 ( .A(n130), .B(n1307), .C(n1549), .Y(n2144) );
  NAND2X1 U1299 ( .A(\mem<18><12> ), .B(n1239), .Y(n1550) );
  OAI21X1 U1300 ( .A(n130), .B(n1309), .C(n1550), .Y(n2143) );
  NAND2X1 U1301 ( .A(\mem<18><13> ), .B(n1239), .Y(n1551) );
  OAI21X1 U1302 ( .A(n130), .B(n1311), .C(n1551), .Y(n2142) );
  NAND2X1 U1303 ( .A(\mem<18><14> ), .B(n1239), .Y(n1552) );
  OAI21X1 U1304 ( .A(n130), .B(n1313), .C(n1552), .Y(n2141) );
  NAND2X1 U1305 ( .A(\mem<18><15> ), .B(n1239), .Y(n1553) );
  OAI21X1 U1306 ( .A(n130), .B(n1315), .C(n1553), .Y(n2140) );
  NAND2X1 U1307 ( .A(\mem<17><0> ), .B(n1240), .Y(n1554) );
  OAI21X1 U1308 ( .A(n132), .B(n1285), .C(n1554), .Y(n2139) );
  NAND2X1 U1309 ( .A(\mem<17><1> ), .B(n1240), .Y(n1555) );
  OAI21X1 U1310 ( .A(n132), .B(n1287), .C(n1555), .Y(n2138) );
  NAND2X1 U1311 ( .A(\mem<17><2> ), .B(n1240), .Y(n1556) );
  OAI21X1 U1312 ( .A(n132), .B(n1289), .C(n1556), .Y(n2137) );
  NAND2X1 U1313 ( .A(\mem<17><3> ), .B(n1240), .Y(n1557) );
  OAI21X1 U1314 ( .A(n132), .B(n1291), .C(n1557), .Y(n2136) );
  NAND2X1 U1315 ( .A(\mem<17><4> ), .B(n1240), .Y(n1558) );
  OAI21X1 U1316 ( .A(n132), .B(n1293), .C(n1558), .Y(n2135) );
  NAND2X1 U1317 ( .A(\mem<17><5> ), .B(n1240), .Y(n1559) );
  OAI21X1 U1318 ( .A(n132), .B(n1295), .C(n1559), .Y(n2134) );
  NAND2X1 U1319 ( .A(\mem<17><6> ), .B(n1240), .Y(n1560) );
  OAI21X1 U1320 ( .A(n132), .B(n1297), .C(n1560), .Y(n2133) );
  NAND2X1 U1321 ( .A(\mem<17><7> ), .B(n1240), .Y(n1561) );
  OAI21X1 U1322 ( .A(n132), .B(n1299), .C(n1561), .Y(n2132) );
  NAND2X1 U1323 ( .A(\mem<17><8> ), .B(n1241), .Y(n1562) );
  OAI21X1 U1324 ( .A(n132), .B(n1301), .C(n1562), .Y(n2131) );
  NAND2X1 U1325 ( .A(\mem<17><9> ), .B(n1241), .Y(n1563) );
  OAI21X1 U1326 ( .A(n132), .B(n1303), .C(n1563), .Y(n2130) );
  NAND2X1 U1327 ( .A(\mem<17><10> ), .B(n1241), .Y(n1564) );
  OAI21X1 U1328 ( .A(n132), .B(n1305), .C(n1564), .Y(n2129) );
  NAND2X1 U1329 ( .A(\mem<17><11> ), .B(n1241), .Y(n1565) );
  OAI21X1 U1330 ( .A(n132), .B(n1307), .C(n1565), .Y(n2128) );
  NAND2X1 U1331 ( .A(\mem<17><12> ), .B(n1241), .Y(n1566) );
  OAI21X1 U1332 ( .A(n132), .B(n1309), .C(n1566), .Y(n2127) );
  NAND2X1 U1333 ( .A(\mem<17><13> ), .B(n1241), .Y(n1567) );
  OAI21X1 U1334 ( .A(n132), .B(n1311), .C(n1567), .Y(n2126) );
  NAND2X1 U1335 ( .A(\mem<17><14> ), .B(n1241), .Y(n1568) );
  OAI21X1 U1336 ( .A(n132), .B(n1313), .C(n1568), .Y(n2125) );
  NAND2X1 U1337 ( .A(\mem<17><15> ), .B(n1241), .Y(n1569) );
  OAI21X1 U1338 ( .A(n132), .B(n1315), .C(n1569), .Y(n2124) );
  NAND2X1 U1339 ( .A(\mem<16><0> ), .B(n1243), .Y(n1570) );
  OAI21X1 U1340 ( .A(n1242), .B(n1285), .C(n1570), .Y(n2123) );
  NAND2X1 U1341 ( .A(\mem<16><1> ), .B(n1243), .Y(n1571) );
  OAI21X1 U1342 ( .A(n1242), .B(n1287), .C(n1571), .Y(n2122) );
  NAND2X1 U1343 ( .A(\mem<16><2> ), .B(n1243), .Y(n1572) );
  OAI21X1 U1344 ( .A(n1242), .B(n1289), .C(n1572), .Y(n2121) );
  NAND2X1 U1345 ( .A(\mem<16><3> ), .B(n1243), .Y(n1573) );
  OAI21X1 U1346 ( .A(n1242), .B(n1291), .C(n1573), .Y(n2120) );
  NAND2X1 U1347 ( .A(\mem<16><4> ), .B(n1243), .Y(n1574) );
  OAI21X1 U1348 ( .A(n1242), .B(n1293), .C(n1574), .Y(n2119) );
  NAND2X1 U1349 ( .A(\mem<16><5> ), .B(n1243), .Y(n1575) );
  OAI21X1 U1350 ( .A(n1242), .B(n1295), .C(n1575), .Y(n2118) );
  NAND2X1 U1351 ( .A(\mem<16><6> ), .B(n1243), .Y(n1576) );
  OAI21X1 U1352 ( .A(n1242), .B(n1297), .C(n1576), .Y(n2117) );
  NAND2X1 U1353 ( .A(\mem<16><7> ), .B(n1243), .Y(n1577) );
  OAI21X1 U1354 ( .A(n1242), .B(n1299), .C(n1577), .Y(n2116) );
  NAND2X1 U1355 ( .A(\mem<16><8> ), .B(n1244), .Y(n1578) );
  OAI21X1 U1356 ( .A(n1242), .B(n1301), .C(n1578), .Y(n2115) );
  NAND2X1 U1357 ( .A(\mem<16><9> ), .B(n1244), .Y(n1579) );
  OAI21X1 U1358 ( .A(n1242), .B(n1303), .C(n1579), .Y(n2114) );
  NAND2X1 U1359 ( .A(\mem<16><10> ), .B(n1244), .Y(n1580) );
  OAI21X1 U1360 ( .A(n1242), .B(n1305), .C(n1580), .Y(n2113) );
  NAND2X1 U1361 ( .A(\mem<16><11> ), .B(n1244), .Y(n1581) );
  OAI21X1 U1362 ( .A(n1242), .B(n1307), .C(n1581), .Y(n2112) );
  NAND2X1 U1363 ( .A(\mem<16><12> ), .B(n1244), .Y(n1582) );
  OAI21X1 U1364 ( .A(n1242), .B(n1309), .C(n1582), .Y(n2111) );
  NAND2X1 U1365 ( .A(\mem<16><13> ), .B(n1244), .Y(n1583) );
  OAI21X1 U1366 ( .A(n1242), .B(n1311), .C(n1583), .Y(n2110) );
  NAND2X1 U1367 ( .A(\mem<16><14> ), .B(n1244), .Y(n1584) );
  OAI21X1 U1368 ( .A(n1242), .B(n1313), .C(n1584), .Y(n2109) );
  NAND2X1 U1369 ( .A(\mem<16><15> ), .B(n1244), .Y(n1585) );
  OAI21X1 U1370 ( .A(n1242), .B(n1315), .C(n1585), .Y(n2108) );
  NAND3X1 U1371 ( .A(n1172), .B(n2364), .C(n1324), .Y(n1586) );
  NAND2X1 U1372 ( .A(\mem<15><0> ), .B(n1245), .Y(n1587) );
  OAI21X1 U1373 ( .A(n134), .B(n1285), .C(n1587), .Y(n2107) );
  NAND2X1 U1374 ( .A(\mem<15><1> ), .B(n1245), .Y(n1588) );
  OAI21X1 U1375 ( .A(n134), .B(n1287), .C(n1588), .Y(n2106) );
  NAND2X1 U1376 ( .A(\mem<15><2> ), .B(n1245), .Y(n1589) );
  OAI21X1 U1377 ( .A(n134), .B(n1289), .C(n1589), .Y(n2105) );
  NAND2X1 U1378 ( .A(\mem<15><3> ), .B(n1245), .Y(n1590) );
  OAI21X1 U1379 ( .A(n134), .B(n1291), .C(n1590), .Y(n2104) );
  NAND2X1 U1380 ( .A(\mem<15><4> ), .B(n1245), .Y(n1591) );
  OAI21X1 U1381 ( .A(n134), .B(n1293), .C(n1591), .Y(n2103) );
  NAND2X1 U1382 ( .A(\mem<15><5> ), .B(n1245), .Y(n1592) );
  OAI21X1 U1383 ( .A(n134), .B(n1295), .C(n1592), .Y(n2102) );
  NAND2X1 U1384 ( .A(\mem<15><6> ), .B(n1245), .Y(n1593) );
  OAI21X1 U1385 ( .A(n134), .B(n1297), .C(n1593), .Y(n2101) );
  NAND2X1 U1386 ( .A(\mem<15><7> ), .B(n1245), .Y(n1594) );
  OAI21X1 U1387 ( .A(n134), .B(n1299), .C(n1594), .Y(n2100) );
  NAND2X1 U1388 ( .A(\mem<15><8> ), .B(n1246), .Y(n1595) );
  OAI21X1 U1389 ( .A(n134), .B(n1301), .C(n1595), .Y(n2099) );
  NAND2X1 U1390 ( .A(\mem<15><9> ), .B(n1246), .Y(n1596) );
  OAI21X1 U1391 ( .A(n134), .B(n1303), .C(n1596), .Y(n2098) );
  NAND2X1 U1392 ( .A(\mem<15><10> ), .B(n1246), .Y(n1597) );
  OAI21X1 U1393 ( .A(n134), .B(n1305), .C(n1597), .Y(n2097) );
  NAND2X1 U1394 ( .A(\mem<15><11> ), .B(n1246), .Y(n1598) );
  OAI21X1 U1395 ( .A(n134), .B(n1307), .C(n1598), .Y(n2096) );
  NAND2X1 U1396 ( .A(\mem<15><12> ), .B(n1246), .Y(n1599) );
  OAI21X1 U1397 ( .A(n134), .B(n1309), .C(n1599), .Y(n2095) );
  NAND2X1 U1398 ( .A(\mem<15><13> ), .B(n1246), .Y(n1600) );
  OAI21X1 U1399 ( .A(n134), .B(n1311), .C(n1600), .Y(n2094) );
  NAND2X1 U1400 ( .A(\mem<15><14> ), .B(n1246), .Y(n1601) );
  OAI21X1 U1401 ( .A(n134), .B(n1313), .C(n1601), .Y(n2093) );
  NAND2X1 U1402 ( .A(\mem<15><15> ), .B(n1246), .Y(n1602) );
  OAI21X1 U1403 ( .A(n134), .B(n1315), .C(n1602), .Y(n2092) );
  NAND2X1 U1404 ( .A(\mem<14><0> ), .B(n1247), .Y(n1603) );
  OAI21X1 U1405 ( .A(n136), .B(n1285), .C(n1603), .Y(n2091) );
  NAND2X1 U1406 ( .A(\mem<14><1> ), .B(n1247), .Y(n1604) );
  OAI21X1 U1407 ( .A(n136), .B(n1287), .C(n1604), .Y(n2090) );
  NAND2X1 U1408 ( .A(\mem<14><2> ), .B(n1247), .Y(n1605) );
  OAI21X1 U1409 ( .A(n136), .B(n1289), .C(n1605), .Y(n2089) );
  NAND2X1 U1410 ( .A(\mem<14><3> ), .B(n1247), .Y(n1606) );
  OAI21X1 U1411 ( .A(n136), .B(n1291), .C(n1606), .Y(n2088) );
  NAND2X1 U1412 ( .A(\mem<14><4> ), .B(n1247), .Y(n1607) );
  OAI21X1 U1413 ( .A(n136), .B(n1293), .C(n1607), .Y(n2087) );
  NAND2X1 U1414 ( .A(\mem<14><5> ), .B(n1247), .Y(n1608) );
  OAI21X1 U1415 ( .A(n136), .B(n1295), .C(n1608), .Y(n2086) );
  NAND2X1 U1416 ( .A(\mem<14><6> ), .B(n1247), .Y(n1609) );
  OAI21X1 U1417 ( .A(n136), .B(n1297), .C(n1609), .Y(n2085) );
  NAND2X1 U1418 ( .A(\mem<14><7> ), .B(n1247), .Y(n1610) );
  OAI21X1 U1419 ( .A(n136), .B(n1299), .C(n1610), .Y(n2084) );
  NAND2X1 U1420 ( .A(\mem<14><8> ), .B(n1248), .Y(n1611) );
  OAI21X1 U1421 ( .A(n136), .B(n1301), .C(n1611), .Y(n2083) );
  NAND2X1 U1422 ( .A(\mem<14><9> ), .B(n1248), .Y(n1612) );
  OAI21X1 U1423 ( .A(n136), .B(n1303), .C(n1612), .Y(n2082) );
  NAND2X1 U1424 ( .A(\mem<14><10> ), .B(n1248), .Y(n1613) );
  OAI21X1 U1425 ( .A(n136), .B(n1305), .C(n1613), .Y(n2081) );
  NAND2X1 U1426 ( .A(\mem<14><11> ), .B(n1248), .Y(n1614) );
  OAI21X1 U1427 ( .A(n136), .B(n1307), .C(n1614), .Y(n2080) );
  NAND2X1 U1428 ( .A(\mem<14><12> ), .B(n1248), .Y(n1615) );
  OAI21X1 U1429 ( .A(n136), .B(n1309), .C(n1615), .Y(n2079) );
  NAND2X1 U1430 ( .A(\mem<14><13> ), .B(n1248), .Y(n1616) );
  OAI21X1 U1431 ( .A(n136), .B(n1311), .C(n1616), .Y(n2078) );
  NAND2X1 U1432 ( .A(\mem<14><14> ), .B(n1248), .Y(n1617) );
  OAI21X1 U1433 ( .A(n136), .B(n1313), .C(n1617), .Y(n2077) );
  NAND2X1 U1434 ( .A(\mem<14><15> ), .B(n1248), .Y(n1618) );
  OAI21X1 U1435 ( .A(n136), .B(n1315), .C(n1618), .Y(n2076) );
  NAND2X1 U1436 ( .A(\mem<13><0> ), .B(n1249), .Y(n1619) );
  OAI21X1 U1437 ( .A(n138), .B(n1285), .C(n1619), .Y(n2075) );
  NAND2X1 U1438 ( .A(\mem<13><1> ), .B(n1249), .Y(n1620) );
  OAI21X1 U1439 ( .A(n138), .B(n1287), .C(n1620), .Y(n2074) );
  NAND2X1 U1440 ( .A(\mem<13><2> ), .B(n1249), .Y(n1621) );
  OAI21X1 U1441 ( .A(n138), .B(n1289), .C(n1621), .Y(n2073) );
  NAND2X1 U1442 ( .A(\mem<13><3> ), .B(n1249), .Y(n1622) );
  OAI21X1 U1443 ( .A(n138), .B(n1291), .C(n1622), .Y(n2072) );
  NAND2X1 U1444 ( .A(\mem<13><4> ), .B(n1249), .Y(n1623) );
  OAI21X1 U1445 ( .A(n138), .B(n1293), .C(n1623), .Y(n2071) );
  NAND2X1 U1446 ( .A(\mem<13><5> ), .B(n1249), .Y(n1624) );
  OAI21X1 U1447 ( .A(n138), .B(n1295), .C(n1624), .Y(n2070) );
  NAND2X1 U1448 ( .A(\mem<13><6> ), .B(n1249), .Y(n1625) );
  OAI21X1 U1449 ( .A(n138), .B(n1297), .C(n1625), .Y(n2069) );
  NAND2X1 U1450 ( .A(\mem<13><7> ), .B(n1249), .Y(n1626) );
  OAI21X1 U1451 ( .A(n138), .B(n1299), .C(n1626), .Y(n2068) );
  NAND2X1 U1452 ( .A(\mem<13><8> ), .B(n1250), .Y(n1627) );
  OAI21X1 U1453 ( .A(n138), .B(n1301), .C(n1627), .Y(n2067) );
  NAND2X1 U1454 ( .A(\mem<13><9> ), .B(n1250), .Y(n1628) );
  OAI21X1 U1455 ( .A(n138), .B(n1303), .C(n1628), .Y(n2066) );
  NAND2X1 U1456 ( .A(\mem<13><10> ), .B(n1250), .Y(n1629) );
  OAI21X1 U1457 ( .A(n138), .B(n1305), .C(n1629), .Y(n2065) );
  NAND2X1 U1458 ( .A(\mem<13><11> ), .B(n1250), .Y(n1630) );
  OAI21X1 U1459 ( .A(n138), .B(n1307), .C(n1630), .Y(n2064) );
  NAND2X1 U1460 ( .A(\mem<13><12> ), .B(n1250), .Y(n1631) );
  OAI21X1 U1461 ( .A(n138), .B(n1309), .C(n1631), .Y(n2063) );
  NAND2X1 U1462 ( .A(\mem<13><13> ), .B(n1250), .Y(n1632) );
  OAI21X1 U1463 ( .A(n138), .B(n1311), .C(n1632), .Y(n2062) );
  NAND2X1 U1464 ( .A(\mem<13><14> ), .B(n1250), .Y(n1633) );
  OAI21X1 U1465 ( .A(n138), .B(n1313), .C(n1633), .Y(n2061) );
  NAND2X1 U1466 ( .A(\mem<13><15> ), .B(n1250), .Y(n1634) );
  OAI21X1 U1467 ( .A(n138), .B(n1315), .C(n1634), .Y(n2060) );
  NAND2X1 U1468 ( .A(\mem<12><0> ), .B(n1251), .Y(n1635) );
  OAI21X1 U1469 ( .A(n140), .B(n1285), .C(n1635), .Y(n2059) );
  NAND2X1 U1470 ( .A(\mem<12><1> ), .B(n1251), .Y(n1636) );
  OAI21X1 U1471 ( .A(n140), .B(n1287), .C(n1636), .Y(n2058) );
  NAND2X1 U1472 ( .A(\mem<12><2> ), .B(n1251), .Y(n1637) );
  OAI21X1 U1473 ( .A(n140), .B(n1289), .C(n1637), .Y(n2057) );
  NAND2X1 U1474 ( .A(\mem<12><3> ), .B(n1251), .Y(n1638) );
  OAI21X1 U1475 ( .A(n140), .B(n1291), .C(n1638), .Y(n2056) );
  NAND2X1 U1476 ( .A(\mem<12><4> ), .B(n1251), .Y(n1639) );
  OAI21X1 U1477 ( .A(n140), .B(n1293), .C(n1639), .Y(n2055) );
  NAND2X1 U1478 ( .A(\mem<12><5> ), .B(n1251), .Y(n1640) );
  OAI21X1 U1479 ( .A(n140), .B(n1295), .C(n1640), .Y(n2054) );
  NAND2X1 U1480 ( .A(\mem<12><6> ), .B(n1251), .Y(n1641) );
  OAI21X1 U1481 ( .A(n140), .B(n1297), .C(n1641), .Y(n2053) );
  NAND2X1 U1482 ( .A(\mem<12><7> ), .B(n1251), .Y(n1642) );
  OAI21X1 U1483 ( .A(n140), .B(n1299), .C(n1642), .Y(n2052) );
  NAND2X1 U1484 ( .A(\mem<12><8> ), .B(n1252), .Y(n1643) );
  OAI21X1 U1485 ( .A(n140), .B(n1301), .C(n1643), .Y(n2051) );
  NAND2X1 U1486 ( .A(\mem<12><9> ), .B(n1252), .Y(n1644) );
  OAI21X1 U1487 ( .A(n140), .B(n1303), .C(n1644), .Y(n2050) );
  NAND2X1 U1488 ( .A(\mem<12><10> ), .B(n1252), .Y(n1645) );
  OAI21X1 U1489 ( .A(n140), .B(n1305), .C(n1645), .Y(n2049) );
  NAND2X1 U1490 ( .A(\mem<12><11> ), .B(n1252), .Y(n1646) );
  OAI21X1 U1491 ( .A(n140), .B(n1307), .C(n1646), .Y(n2048) );
  NAND2X1 U1492 ( .A(\mem<12><12> ), .B(n1252), .Y(n1647) );
  OAI21X1 U1493 ( .A(n140), .B(n1309), .C(n1647), .Y(n2047) );
  NAND2X1 U1494 ( .A(\mem<12><13> ), .B(n1252), .Y(n1648) );
  OAI21X1 U1495 ( .A(n140), .B(n1311), .C(n1648), .Y(n2046) );
  NAND2X1 U1496 ( .A(\mem<12><14> ), .B(n1252), .Y(n1649) );
  OAI21X1 U1497 ( .A(n140), .B(n1313), .C(n1649), .Y(n2045) );
  NAND2X1 U1498 ( .A(\mem<12><15> ), .B(n1252), .Y(n1650) );
  OAI21X1 U1499 ( .A(n140), .B(n1315), .C(n1650), .Y(n2044) );
  NAND2X1 U1500 ( .A(\mem<11><0> ), .B(n1253), .Y(n1651) );
  OAI21X1 U1501 ( .A(n142), .B(n1285), .C(n1651), .Y(n2043) );
  NAND2X1 U1502 ( .A(\mem<11><1> ), .B(n1253), .Y(n1652) );
  OAI21X1 U1503 ( .A(n142), .B(n1286), .C(n1652), .Y(n2042) );
  NAND2X1 U1504 ( .A(\mem<11><2> ), .B(n1253), .Y(n1653) );
  OAI21X1 U1505 ( .A(n142), .B(n1288), .C(n1653), .Y(n2041) );
  NAND2X1 U1506 ( .A(\mem<11><3> ), .B(n1253), .Y(n1654) );
  OAI21X1 U1507 ( .A(n142), .B(n1290), .C(n1654), .Y(n2040) );
  NAND2X1 U1508 ( .A(\mem<11><4> ), .B(n1253), .Y(n1655) );
  OAI21X1 U1509 ( .A(n142), .B(n1292), .C(n1655), .Y(n2039) );
  NAND2X1 U1510 ( .A(\mem<11><5> ), .B(n1253), .Y(n1656) );
  OAI21X1 U1511 ( .A(n142), .B(n1294), .C(n1656), .Y(n2038) );
  NAND2X1 U1512 ( .A(\mem<11><6> ), .B(n1253), .Y(n1657) );
  OAI21X1 U1513 ( .A(n142), .B(n1296), .C(n1657), .Y(n2037) );
  NAND2X1 U1514 ( .A(\mem<11><7> ), .B(n1253), .Y(n1658) );
  OAI21X1 U1515 ( .A(n142), .B(n1298), .C(n1658), .Y(n2036) );
  NAND2X1 U1516 ( .A(\mem<11><8> ), .B(n1254), .Y(n1659) );
  OAI21X1 U1517 ( .A(n142), .B(n1300), .C(n1659), .Y(n2035) );
  NAND2X1 U1518 ( .A(\mem<11><9> ), .B(n1254), .Y(n1660) );
  OAI21X1 U1519 ( .A(n142), .B(n1302), .C(n1660), .Y(n2034) );
  NAND2X1 U1520 ( .A(\mem<11><10> ), .B(n1254), .Y(n1661) );
  OAI21X1 U1521 ( .A(n142), .B(n1304), .C(n1661), .Y(n2033) );
  NAND2X1 U1522 ( .A(\mem<11><11> ), .B(n1254), .Y(n1662) );
  OAI21X1 U1523 ( .A(n142), .B(n1306), .C(n1662), .Y(n2032) );
  NAND2X1 U1524 ( .A(\mem<11><12> ), .B(n1254), .Y(n1663) );
  OAI21X1 U1525 ( .A(n142), .B(n1308), .C(n1663), .Y(n2031) );
  NAND2X1 U1526 ( .A(\mem<11><13> ), .B(n1254), .Y(n1664) );
  OAI21X1 U1527 ( .A(n142), .B(n1310), .C(n1664), .Y(n2030) );
  NAND2X1 U1528 ( .A(\mem<11><14> ), .B(n1254), .Y(n1665) );
  OAI21X1 U1529 ( .A(n142), .B(n1312), .C(n1665), .Y(n2029) );
  NAND2X1 U1530 ( .A(\mem<11><15> ), .B(n1254), .Y(n1666) );
  OAI21X1 U1531 ( .A(n142), .B(n1314), .C(n1666), .Y(n2028) );
  NAND2X1 U1532 ( .A(\mem<10><0> ), .B(n1255), .Y(n1667) );
  OAI21X1 U1533 ( .A(n144), .B(n1285), .C(n1667), .Y(n2027) );
  NAND2X1 U1534 ( .A(\mem<10><1> ), .B(n1255), .Y(n1668) );
  OAI21X1 U1535 ( .A(n144), .B(n1286), .C(n1668), .Y(n2026) );
  NAND2X1 U1536 ( .A(\mem<10><2> ), .B(n1255), .Y(n1669) );
  OAI21X1 U1537 ( .A(n144), .B(n1288), .C(n1669), .Y(n2025) );
  NAND2X1 U1538 ( .A(\mem<10><3> ), .B(n1255), .Y(n1670) );
  OAI21X1 U1539 ( .A(n144), .B(n1290), .C(n1670), .Y(n2024) );
  NAND2X1 U1540 ( .A(\mem<10><4> ), .B(n1255), .Y(n1671) );
  OAI21X1 U1541 ( .A(n144), .B(n1292), .C(n1671), .Y(n2023) );
  NAND2X1 U1542 ( .A(\mem<10><5> ), .B(n1255), .Y(n1672) );
  OAI21X1 U1543 ( .A(n144), .B(n1294), .C(n1672), .Y(n2022) );
  NAND2X1 U1544 ( .A(\mem<10><6> ), .B(n1255), .Y(n1673) );
  OAI21X1 U1545 ( .A(n144), .B(n1296), .C(n1673), .Y(n2021) );
  NAND2X1 U1546 ( .A(\mem<10><7> ), .B(n1255), .Y(n1674) );
  OAI21X1 U1547 ( .A(n144), .B(n1298), .C(n1674), .Y(n2020) );
  NAND2X1 U1548 ( .A(\mem<10><8> ), .B(n1256), .Y(n1675) );
  OAI21X1 U1549 ( .A(n144), .B(n1300), .C(n1675), .Y(n2019) );
  NAND2X1 U1550 ( .A(\mem<10><9> ), .B(n1256), .Y(n1676) );
  OAI21X1 U1551 ( .A(n144), .B(n1302), .C(n1676), .Y(n2018) );
  NAND2X1 U1552 ( .A(\mem<10><10> ), .B(n1256), .Y(n1677) );
  OAI21X1 U1553 ( .A(n144), .B(n1304), .C(n1677), .Y(n2017) );
  NAND2X1 U1554 ( .A(\mem<10><11> ), .B(n1256), .Y(n1678) );
  OAI21X1 U1555 ( .A(n144), .B(n1306), .C(n1678), .Y(n2016) );
  NAND2X1 U1556 ( .A(\mem<10><12> ), .B(n1256), .Y(n1679) );
  OAI21X1 U1557 ( .A(n144), .B(n1308), .C(n1679), .Y(n2015) );
  NAND2X1 U1558 ( .A(\mem<10><13> ), .B(n1256), .Y(n1680) );
  OAI21X1 U1559 ( .A(n144), .B(n1310), .C(n1680), .Y(n2014) );
  NAND2X1 U1560 ( .A(\mem<10><14> ), .B(n1256), .Y(n1681) );
  OAI21X1 U1561 ( .A(n144), .B(n1312), .C(n1681), .Y(n2013) );
  NAND2X1 U1562 ( .A(\mem<10><15> ), .B(n1256), .Y(n1682) );
  OAI21X1 U1563 ( .A(n144), .B(n1314), .C(n1682), .Y(n2012) );
  NAND2X1 U1564 ( .A(\mem<9><0> ), .B(n1257), .Y(n1683) );
  OAI21X1 U1565 ( .A(n146), .B(n1285), .C(n1683), .Y(n2011) );
  NAND2X1 U1566 ( .A(\mem<9><1> ), .B(n1257), .Y(n1684) );
  OAI21X1 U1567 ( .A(n146), .B(n1286), .C(n1684), .Y(n2010) );
  NAND2X1 U1568 ( .A(\mem<9><2> ), .B(n1257), .Y(n1685) );
  OAI21X1 U1569 ( .A(n146), .B(n1288), .C(n1685), .Y(n2009) );
  NAND2X1 U1570 ( .A(\mem<9><3> ), .B(n1257), .Y(n1686) );
  OAI21X1 U1571 ( .A(n146), .B(n1290), .C(n1686), .Y(n2008) );
  NAND2X1 U1572 ( .A(\mem<9><4> ), .B(n1257), .Y(n1687) );
  OAI21X1 U1573 ( .A(n146), .B(n1292), .C(n1687), .Y(n2007) );
  NAND2X1 U1574 ( .A(\mem<9><5> ), .B(n1257), .Y(n1688) );
  OAI21X1 U1575 ( .A(n146), .B(n1294), .C(n1688), .Y(n2006) );
  NAND2X1 U1576 ( .A(\mem<9><6> ), .B(n1257), .Y(n1689) );
  OAI21X1 U1577 ( .A(n146), .B(n1296), .C(n1689), .Y(n2005) );
  NAND2X1 U1578 ( .A(\mem<9><7> ), .B(n1257), .Y(n1690) );
  OAI21X1 U1579 ( .A(n146), .B(n1298), .C(n1690), .Y(n2004) );
  NAND2X1 U1580 ( .A(\mem<9><8> ), .B(n1258), .Y(n1691) );
  OAI21X1 U1581 ( .A(n146), .B(n1300), .C(n1691), .Y(n2003) );
  NAND2X1 U1582 ( .A(\mem<9><9> ), .B(n1258), .Y(n1692) );
  OAI21X1 U1583 ( .A(n146), .B(n1302), .C(n1692), .Y(n2002) );
  NAND2X1 U1584 ( .A(\mem<9><10> ), .B(n1258), .Y(n1693) );
  OAI21X1 U1585 ( .A(n146), .B(n1304), .C(n1693), .Y(n2001) );
  NAND2X1 U1586 ( .A(\mem<9><11> ), .B(n1258), .Y(n1694) );
  OAI21X1 U1587 ( .A(n146), .B(n1306), .C(n1694), .Y(n2000) );
  NAND2X1 U1588 ( .A(\mem<9><12> ), .B(n1258), .Y(n1695) );
  OAI21X1 U1589 ( .A(n146), .B(n1308), .C(n1695), .Y(n1999) );
  NAND2X1 U1590 ( .A(\mem<9><13> ), .B(n1258), .Y(n1696) );
  OAI21X1 U1591 ( .A(n146), .B(n1310), .C(n1696), .Y(n1998) );
  NAND2X1 U1592 ( .A(\mem<9><14> ), .B(n1258), .Y(n1697) );
  OAI21X1 U1593 ( .A(n146), .B(n1312), .C(n1697), .Y(n1997) );
  NAND2X1 U1594 ( .A(\mem<9><15> ), .B(n1258), .Y(n1698) );
  OAI21X1 U1595 ( .A(n146), .B(n1314), .C(n1698), .Y(n1996) );
  NAND2X1 U1596 ( .A(\mem<8><0> ), .B(n1260), .Y(n1700) );
  OAI21X1 U1597 ( .A(n1259), .B(n1285), .C(n1700), .Y(n1995) );
  NAND2X1 U1598 ( .A(\mem<8><1> ), .B(n1260), .Y(n1701) );
  OAI21X1 U1599 ( .A(n1259), .B(n1286), .C(n1701), .Y(n1994) );
  NAND2X1 U1600 ( .A(\mem<8><2> ), .B(n1260), .Y(n1702) );
  OAI21X1 U1601 ( .A(n1259), .B(n1288), .C(n1702), .Y(n1993) );
  NAND2X1 U1602 ( .A(\mem<8><3> ), .B(n1260), .Y(n1703) );
  OAI21X1 U1603 ( .A(n1259), .B(n1290), .C(n1703), .Y(n1992) );
  NAND2X1 U1604 ( .A(\mem<8><4> ), .B(n1260), .Y(n1704) );
  OAI21X1 U1605 ( .A(n1259), .B(n1292), .C(n1704), .Y(n1991) );
  NAND2X1 U1606 ( .A(\mem<8><5> ), .B(n1260), .Y(n1705) );
  OAI21X1 U1607 ( .A(n1259), .B(n1294), .C(n1705), .Y(n1990) );
  NAND2X1 U1608 ( .A(\mem<8><6> ), .B(n1260), .Y(n1706) );
  OAI21X1 U1609 ( .A(n1259), .B(n1296), .C(n1706), .Y(n1989) );
  NAND2X1 U1610 ( .A(\mem<8><7> ), .B(n1260), .Y(n1707) );
  OAI21X1 U1611 ( .A(n1259), .B(n1298), .C(n1707), .Y(n1988) );
  NAND2X1 U1612 ( .A(\mem<8><8> ), .B(n1261), .Y(n1708) );
  OAI21X1 U1613 ( .A(n1259), .B(n1300), .C(n1708), .Y(n1987) );
  NAND2X1 U1614 ( .A(\mem<8><9> ), .B(n1261), .Y(n1709) );
  OAI21X1 U1615 ( .A(n1259), .B(n1302), .C(n1709), .Y(n1986) );
  NAND2X1 U1616 ( .A(\mem<8><10> ), .B(n1261), .Y(n1710) );
  OAI21X1 U1617 ( .A(n1259), .B(n1304), .C(n1710), .Y(n1985) );
  NAND2X1 U1618 ( .A(\mem<8><11> ), .B(n1261), .Y(n1711) );
  OAI21X1 U1619 ( .A(n1259), .B(n1306), .C(n1711), .Y(n1984) );
  NAND2X1 U1620 ( .A(\mem<8><12> ), .B(n1261), .Y(n1712) );
  OAI21X1 U1621 ( .A(n1259), .B(n1308), .C(n1712), .Y(n1983) );
  NAND2X1 U1622 ( .A(\mem<8><13> ), .B(n1261), .Y(n1713) );
  OAI21X1 U1623 ( .A(n1259), .B(n1310), .C(n1713), .Y(n1982) );
  NAND2X1 U1624 ( .A(\mem<8><14> ), .B(n1261), .Y(n1714) );
  OAI21X1 U1625 ( .A(n1259), .B(n1312), .C(n1714), .Y(n1981) );
  NAND2X1 U1626 ( .A(\mem<8><15> ), .B(n1261), .Y(n1715) );
  OAI21X1 U1627 ( .A(n1259), .B(n1314), .C(n1715), .Y(n1980) );
  NAND3X1 U1628 ( .A(n1323), .B(n2364), .C(n1324), .Y(n1716) );
  NAND2X1 U1629 ( .A(\mem<7><0> ), .B(n1262), .Y(n1717) );
  OAI21X1 U1630 ( .A(n148), .B(n1284), .C(n1717), .Y(n1979) );
  NAND2X1 U1631 ( .A(\mem<7><1> ), .B(n1262), .Y(n1718) );
  OAI21X1 U1632 ( .A(n148), .B(n1286), .C(n1718), .Y(n1978) );
  NAND2X1 U1633 ( .A(\mem<7><2> ), .B(n1262), .Y(n1719) );
  OAI21X1 U1634 ( .A(n148), .B(n1288), .C(n1719), .Y(n1977) );
  NAND2X1 U1635 ( .A(\mem<7><3> ), .B(n1262), .Y(n1720) );
  OAI21X1 U1636 ( .A(n148), .B(n1290), .C(n1720), .Y(n1976) );
  NAND2X1 U1637 ( .A(\mem<7><4> ), .B(n1262), .Y(n1721) );
  OAI21X1 U1638 ( .A(n148), .B(n1292), .C(n1721), .Y(n1975) );
  NAND2X1 U1639 ( .A(\mem<7><5> ), .B(n1262), .Y(n1722) );
  OAI21X1 U1640 ( .A(n148), .B(n1294), .C(n1722), .Y(n1974) );
  NAND2X1 U1641 ( .A(\mem<7><6> ), .B(n1262), .Y(n1723) );
  OAI21X1 U1642 ( .A(n148), .B(n1296), .C(n1723), .Y(n1973) );
  NAND2X1 U1643 ( .A(\mem<7><7> ), .B(n1262), .Y(n1724) );
  OAI21X1 U1644 ( .A(n148), .B(n1298), .C(n1724), .Y(n1972) );
  NAND2X1 U1645 ( .A(\mem<7><8> ), .B(n1263), .Y(n1725) );
  OAI21X1 U1646 ( .A(n148), .B(n1300), .C(n1725), .Y(n1971) );
  NAND2X1 U1647 ( .A(\mem<7><9> ), .B(n1263), .Y(n1726) );
  OAI21X1 U1648 ( .A(n148), .B(n1302), .C(n1726), .Y(n1970) );
  NAND2X1 U1649 ( .A(\mem<7><10> ), .B(n1263), .Y(n1727) );
  OAI21X1 U1650 ( .A(n148), .B(n1304), .C(n1727), .Y(n1969) );
  NAND2X1 U1651 ( .A(\mem<7><11> ), .B(n1263), .Y(n1728) );
  OAI21X1 U1652 ( .A(n148), .B(n1306), .C(n1728), .Y(n1968) );
  NAND2X1 U1653 ( .A(\mem<7><12> ), .B(n1263), .Y(n1729) );
  OAI21X1 U1654 ( .A(n148), .B(n1308), .C(n1729), .Y(n1967) );
  NAND2X1 U1655 ( .A(\mem<7><13> ), .B(n1263), .Y(n1730) );
  OAI21X1 U1656 ( .A(n148), .B(n1310), .C(n1730), .Y(n1966) );
  NAND2X1 U1657 ( .A(\mem<7><14> ), .B(n1263), .Y(n1731) );
  OAI21X1 U1658 ( .A(n148), .B(n1312), .C(n1731), .Y(n1965) );
  NAND2X1 U1659 ( .A(\mem<7><15> ), .B(n1263), .Y(n1732) );
  OAI21X1 U1660 ( .A(n148), .B(n1314), .C(n1732), .Y(n1964) );
  NAND2X1 U1661 ( .A(\mem<6><0> ), .B(n1264), .Y(n1733) );
  OAI21X1 U1662 ( .A(n150), .B(n1285), .C(n1733), .Y(n1963) );
  NAND2X1 U1663 ( .A(\mem<6><1> ), .B(n1264), .Y(n1734) );
  OAI21X1 U1664 ( .A(n150), .B(n1286), .C(n1734), .Y(n1962) );
  NAND2X1 U1665 ( .A(\mem<6><2> ), .B(n1264), .Y(n1735) );
  OAI21X1 U1666 ( .A(n150), .B(n1288), .C(n1735), .Y(n1961) );
  NAND2X1 U1667 ( .A(\mem<6><3> ), .B(n1264), .Y(n1736) );
  OAI21X1 U1668 ( .A(n150), .B(n1290), .C(n1736), .Y(n1960) );
  NAND2X1 U1669 ( .A(\mem<6><4> ), .B(n1264), .Y(n1737) );
  OAI21X1 U1670 ( .A(n150), .B(n1292), .C(n1737), .Y(n1959) );
  NAND2X1 U1671 ( .A(\mem<6><5> ), .B(n1264), .Y(n1738) );
  OAI21X1 U1672 ( .A(n150), .B(n1294), .C(n1738), .Y(n1958) );
  NAND2X1 U1673 ( .A(\mem<6><6> ), .B(n1264), .Y(n1739) );
  OAI21X1 U1674 ( .A(n150), .B(n1296), .C(n1739), .Y(n1957) );
  NAND2X1 U1675 ( .A(\mem<6><7> ), .B(n1264), .Y(n1740) );
  OAI21X1 U1676 ( .A(n150), .B(n1298), .C(n1740), .Y(n1956) );
  NAND2X1 U1677 ( .A(\mem<6><8> ), .B(n1265), .Y(n1741) );
  OAI21X1 U1678 ( .A(n150), .B(n1300), .C(n1741), .Y(n1955) );
  NAND2X1 U1679 ( .A(\mem<6><9> ), .B(n1265), .Y(n1742) );
  OAI21X1 U1680 ( .A(n150), .B(n1302), .C(n1742), .Y(n1954) );
  NAND2X1 U1681 ( .A(\mem<6><10> ), .B(n1265), .Y(n1743) );
  OAI21X1 U1682 ( .A(n150), .B(n1304), .C(n1743), .Y(n1953) );
  NAND2X1 U1683 ( .A(\mem<6><11> ), .B(n1265), .Y(n1744) );
  OAI21X1 U1684 ( .A(n150), .B(n1306), .C(n1744), .Y(n1952) );
  NAND2X1 U1685 ( .A(\mem<6><12> ), .B(n1265), .Y(n1745) );
  OAI21X1 U1686 ( .A(n150), .B(n1308), .C(n1745), .Y(n1951) );
  NAND2X1 U1687 ( .A(\mem<6><13> ), .B(n1265), .Y(n1746) );
  OAI21X1 U1688 ( .A(n150), .B(n1310), .C(n1746), .Y(n1950) );
  NAND2X1 U1689 ( .A(\mem<6><14> ), .B(n1265), .Y(n1747) );
  OAI21X1 U1690 ( .A(n150), .B(n1312), .C(n1747), .Y(n1949) );
  NAND2X1 U1691 ( .A(\mem<6><15> ), .B(n1265), .Y(n1748) );
  OAI21X1 U1692 ( .A(n150), .B(n1314), .C(n1748), .Y(n1948) );
  NAND2X1 U1693 ( .A(\mem<5><0> ), .B(n1266), .Y(n1750) );
  OAI21X1 U1694 ( .A(n152), .B(n1284), .C(n1750), .Y(n1947) );
  NAND2X1 U1695 ( .A(\mem<5><1> ), .B(n1266), .Y(n1751) );
  OAI21X1 U1696 ( .A(n152), .B(n1286), .C(n1751), .Y(n1946) );
  NAND2X1 U1697 ( .A(\mem<5><2> ), .B(n1266), .Y(n1752) );
  OAI21X1 U1698 ( .A(n152), .B(n1288), .C(n1752), .Y(n1945) );
  NAND2X1 U1699 ( .A(\mem<5><3> ), .B(n1266), .Y(n1753) );
  OAI21X1 U1700 ( .A(n152), .B(n1290), .C(n1753), .Y(n1944) );
  NAND2X1 U1701 ( .A(\mem<5><4> ), .B(n1266), .Y(n1754) );
  OAI21X1 U1702 ( .A(n152), .B(n1292), .C(n1754), .Y(n1943) );
  NAND2X1 U1703 ( .A(\mem<5><5> ), .B(n1266), .Y(n1755) );
  OAI21X1 U1704 ( .A(n152), .B(n1294), .C(n1755), .Y(n1942) );
  NAND2X1 U1705 ( .A(\mem<5><6> ), .B(n1266), .Y(n1756) );
  OAI21X1 U1706 ( .A(n152), .B(n1296), .C(n1756), .Y(n1941) );
  NAND2X1 U1707 ( .A(\mem<5><7> ), .B(n1266), .Y(n1757) );
  OAI21X1 U1708 ( .A(n152), .B(n1298), .C(n1757), .Y(n1940) );
  NAND2X1 U1709 ( .A(\mem<5><8> ), .B(n1267), .Y(n1758) );
  OAI21X1 U1710 ( .A(n152), .B(n1300), .C(n1758), .Y(n1939) );
  NAND2X1 U1711 ( .A(\mem<5><9> ), .B(n1267), .Y(n1759) );
  OAI21X1 U1712 ( .A(n152), .B(n1302), .C(n1759), .Y(n1938) );
  NAND2X1 U1713 ( .A(\mem<5><10> ), .B(n1267), .Y(n1760) );
  OAI21X1 U1714 ( .A(n152), .B(n1304), .C(n1760), .Y(n1937) );
  NAND2X1 U1715 ( .A(\mem<5><11> ), .B(n1267), .Y(n1761) );
  OAI21X1 U1716 ( .A(n152), .B(n1306), .C(n1761), .Y(n1936) );
  NAND2X1 U1717 ( .A(\mem<5><12> ), .B(n1267), .Y(n1762) );
  OAI21X1 U1718 ( .A(n152), .B(n1308), .C(n1762), .Y(n1935) );
  NAND2X1 U1719 ( .A(\mem<5><13> ), .B(n1267), .Y(n1763) );
  OAI21X1 U1720 ( .A(n152), .B(n1310), .C(n1763), .Y(n1934) );
  NAND2X1 U1721 ( .A(\mem<5><14> ), .B(n1267), .Y(n1764) );
  OAI21X1 U1722 ( .A(n152), .B(n1312), .C(n1764), .Y(n1933) );
  NAND2X1 U1723 ( .A(\mem<5><15> ), .B(n1267), .Y(n1765) );
  OAI21X1 U1724 ( .A(n152), .B(n1314), .C(n1765), .Y(n1932) );
  NAND2X1 U1725 ( .A(\mem<4><0> ), .B(n1268), .Y(n1767) );
  OAI21X1 U1726 ( .A(n154), .B(n1285), .C(n1767), .Y(n1931) );
  NAND2X1 U1727 ( .A(\mem<4><1> ), .B(n1268), .Y(n1768) );
  OAI21X1 U1728 ( .A(n154), .B(n1286), .C(n1768), .Y(n1930) );
  NAND2X1 U1729 ( .A(\mem<4><2> ), .B(n1268), .Y(n1769) );
  OAI21X1 U1730 ( .A(n154), .B(n1288), .C(n1769), .Y(n1929) );
  NAND2X1 U1731 ( .A(\mem<4><3> ), .B(n1268), .Y(n1770) );
  OAI21X1 U1732 ( .A(n154), .B(n1290), .C(n1770), .Y(n1928) );
  NAND2X1 U1733 ( .A(\mem<4><4> ), .B(n1268), .Y(n1771) );
  OAI21X1 U1734 ( .A(n154), .B(n1292), .C(n1771), .Y(n1927) );
  NAND2X1 U1735 ( .A(\mem<4><5> ), .B(n1268), .Y(n1772) );
  OAI21X1 U1736 ( .A(n154), .B(n1294), .C(n1772), .Y(n1926) );
  NAND2X1 U1737 ( .A(\mem<4><6> ), .B(n1268), .Y(n1773) );
  OAI21X1 U1738 ( .A(n154), .B(n1296), .C(n1773), .Y(n1925) );
  NAND2X1 U1739 ( .A(\mem<4><7> ), .B(n1268), .Y(n1774) );
  OAI21X1 U1740 ( .A(n154), .B(n1298), .C(n1774), .Y(n1924) );
  NAND2X1 U1741 ( .A(\mem<4><8> ), .B(n1269), .Y(n1775) );
  OAI21X1 U1742 ( .A(n154), .B(n1300), .C(n1775), .Y(n1923) );
  NAND2X1 U1743 ( .A(\mem<4><9> ), .B(n1269), .Y(n1776) );
  OAI21X1 U1744 ( .A(n154), .B(n1302), .C(n1776), .Y(n1922) );
  NAND2X1 U1745 ( .A(\mem<4><10> ), .B(n1269), .Y(n1777) );
  OAI21X1 U1746 ( .A(n154), .B(n1304), .C(n1777), .Y(n1921) );
  NAND2X1 U1747 ( .A(\mem<4><11> ), .B(n1269), .Y(n1778) );
  OAI21X1 U1748 ( .A(n154), .B(n1306), .C(n1778), .Y(n1920) );
  NAND2X1 U1749 ( .A(\mem<4><12> ), .B(n1269), .Y(n1779) );
  OAI21X1 U1750 ( .A(n154), .B(n1308), .C(n1779), .Y(n1919) );
  NAND2X1 U1751 ( .A(\mem<4><13> ), .B(n1269), .Y(n1780) );
  OAI21X1 U1752 ( .A(n154), .B(n1310), .C(n1780), .Y(n1918) );
  NAND2X1 U1753 ( .A(\mem<4><14> ), .B(n1269), .Y(n1781) );
  OAI21X1 U1754 ( .A(n154), .B(n1312), .C(n1781), .Y(n1917) );
  NAND2X1 U1755 ( .A(\mem<4><15> ), .B(n1269), .Y(n1782) );
  OAI21X1 U1756 ( .A(n154), .B(n1314), .C(n1782), .Y(n1916) );
  NAND2X1 U1757 ( .A(\mem<3><0> ), .B(n1270), .Y(n1784) );
  OAI21X1 U1758 ( .A(n156), .B(n1284), .C(n1784), .Y(n1915) );
  NAND2X1 U1759 ( .A(\mem<3><1> ), .B(n1270), .Y(n1785) );
  OAI21X1 U1760 ( .A(n156), .B(n1286), .C(n1785), .Y(n1914) );
  NAND2X1 U1761 ( .A(\mem<3><2> ), .B(n1270), .Y(n1786) );
  OAI21X1 U1762 ( .A(n156), .B(n1288), .C(n1786), .Y(n1913) );
  NAND2X1 U1763 ( .A(\mem<3><3> ), .B(n1270), .Y(n1787) );
  OAI21X1 U1764 ( .A(n156), .B(n1290), .C(n1787), .Y(n1912) );
  NAND2X1 U1765 ( .A(\mem<3><4> ), .B(n1270), .Y(n1788) );
  OAI21X1 U1766 ( .A(n156), .B(n1292), .C(n1788), .Y(n1911) );
  NAND2X1 U1767 ( .A(\mem<3><5> ), .B(n1270), .Y(n1789) );
  OAI21X1 U1768 ( .A(n156), .B(n1294), .C(n1789), .Y(n1910) );
  NAND2X1 U1769 ( .A(\mem<3><6> ), .B(n1270), .Y(n1790) );
  OAI21X1 U1770 ( .A(n156), .B(n1296), .C(n1790), .Y(n1909) );
  NAND2X1 U1771 ( .A(\mem<3><7> ), .B(n1270), .Y(n1791) );
  OAI21X1 U1772 ( .A(n156), .B(n1298), .C(n1791), .Y(n1908) );
  NAND2X1 U1773 ( .A(\mem<3><8> ), .B(n1271), .Y(n1792) );
  OAI21X1 U1774 ( .A(n156), .B(n1300), .C(n1792), .Y(n1907) );
  NAND2X1 U1775 ( .A(\mem<3><9> ), .B(n1271), .Y(n1793) );
  OAI21X1 U1776 ( .A(n156), .B(n1302), .C(n1793), .Y(n1906) );
  NAND2X1 U1777 ( .A(\mem<3><10> ), .B(n1271), .Y(n1794) );
  OAI21X1 U1778 ( .A(n156), .B(n1304), .C(n1794), .Y(n1905) );
  NAND2X1 U1779 ( .A(\mem<3><11> ), .B(n1271), .Y(n1795) );
  OAI21X1 U1780 ( .A(n156), .B(n1306), .C(n1795), .Y(n1904) );
  NAND2X1 U1781 ( .A(\mem<3><12> ), .B(n1271), .Y(n1796) );
  OAI21X1 U1782 ( .A(n156), .B(n1308), .C(n1796), .Y(n1903) );
  NAND2X1 U1783 ( .A(\mem<3><13> ), .B(n1271), .Y(n1797) );
  OAI21X1 U1784 ( .A(n156), .B(n1310), .C(n1797), .Y(n1902) );
  NAND2X1 U1785 ( .A(\mem<3><14> ), .B(n1271), .Y(n1798) );
  OAI21X1 U1786 ( .A(n156), .B(n1312), .C(n1798), .Y(n1901) );
  NAND2X1 U1787 ( .A(\mem<3><15> ), .B(n1271), .Y(n1799) );
  OAI21X1 U1788 ( .A(n156), .B(n1314), .C(n1799), .Y(n1900) );
  NAND2X1 U1789 ( .A(\mem<2><0> ), .B(n1272), .Y(n1801) );
  OAI21X1 U1790 ( .A(n158), .B(n1285), .C(n1801), .Y(n1899) );
  NAND2X1 U1791 ( .A(\mem<2><1> ), .B(n1272), .Y(n1802) );
  OAI21X1 U1792 ( .A(n158), .B(n1286), .C(n1802), .Y(n1898) );
  NAND2X1 U1793 ( .A(\mem<2><2> ), .B(n1272), .Y(n1803) );
  OAI21X1 U1794 ( .A(n158), .B(n1288), .C(n1803), .Y(n1897) );
  NAND2X1 U1795 ( .A(\mem<2><3> ), .B(n1272), .Y(n1804) );
  OAI21X1 U1796 ( .A(n158), .B(n1290), .C(n1804), .Y(n1896) );
  NAND2X1 U1797 ( .A(\mem<2><4> ), .B(n1272), .Y(n1805) );
  OAI21X1 U1798 ( .A(n158), .B(n1292), .C(n1805), .Y(n1895) );
  NAND2X1 U1799 ( .A(\mem<2><5> ), .B(n1272), .Y(n1806) );
  OAI21X1 U1800 ( .A(n158), .B(n1294), .C(n1806), .Y(n1894) );
  NAND2X1 U1801 ( .A(\mem<2><6> ), .B(n1272), .Y(n1807) );
  OAI21X1 U1802 ( .A(n158), .B(n1296), .C(n1807), .Y(n1893) );
  NAND2X1 U1803 ( .A(\mem<2><7> ), .B(n1272), .Y(n1808) );
  OAI21X1 U1804 ( .A(n158), .B(n1298), .C(n1808), .Y(n1892) );
  NAND2X1 U1805 ( .A(\mem<2><8> ), .B(n1273), .Y(n1809) );
  OAI21X1 U1806 ( .A(n158), .B(n1300), .C(n1809), .Y(n1891) );
  NAND2X1 U1807 ( .A(\mem<2><9> ), .B(n1273), .Y(n1810) );
  OAI21X1 U1808 ( .A(n158), .B(n1302), .C(n1810), .Y(n1890) );
  NAND2X1 U1809 ( .A(\mem<2><10> ), .B(n1273), .Y(n1811) );
  OAI21X1 U1810 ( .A(n158), .B(n1304), .C(n1811), .Y(n1889) );
  NAND2X1 U1811 ( .A(\mem<2><11> ), .B(n1273), .Y(n1812) );
  OAI21X1 U1812 ( .A(n158), .B(n1306), .C(n1812), .Y(n1888) );
  NAND2X1 U1813 ( .A(\mem<2><12> ), .B(n1273), .Y(n1813) );
  OAI21X1 U1814 ( .A(n158), .B(n1308), .C(n1813), .Y(n1887) );
  NAND2X1 U1815 ( .A(\mem<2><13> ), .B(n1273), .Y(n1814) );
  OAI21X1 U1816 ( .A(n158), .B(n1310), .C(n1814), .Y(n1886) );
  NAND2X1 U1817 ( .A(\mem<2><14> ), .B(n1273), .Y(n1815) );
  OAI21X1 U1818 ( .A(n158), .B(n1312), .C(n1815), .Y(n1885) );
  NAND2X1 U1819 ( .A(\mem<2><15> ), .B(n1273), .Y(n1816) );
  OAI21X1 U1820 ( .A(n158), .B(n1314), .C(n1816), .Y(n1884) );
  NAND2X1 U1821 ( .A(\mem<1><0> ), .B(n1274), .Y(n1818) );
  OAI21X1 U1822 ( .A(n160), .B(n1284), .C(n1818), .Y(n1883) );
  NAND2X1 U1823 ( .A(\mem<1><1> ), .B(n1274), .Y(n1819) );
  OAI21X1 U1824 ( .A(n160), .B(n1286), .C(n1819), .Y(n1882) );
  NAND2X1 U1825 ( .A(\mem<1><2> ), .B(n1274), .Y(n1820) );
  OAI21X1 U1826 ( .A(n160), .B(n1288), .C(n1820), .Y(n1881) );
  NAND2X1 U1827 ( .A(\mem<1><3> ), .B(n1274), .Y(n1821) );
  OAI21X1 U1828 ( .A(n160), .B(n1290), .C(n1821), .Y(n1880) );
  NAND2X1 U1829 ( .A(\mem<1><4> ), .B(n1274), .Y(n1822) );
  OAI21X1 U1830 ( .A(n160), .B(n1292), .C(n1822), .Y(n1879) );
  NAND2X1 U1831 ( .A(\mem<1><5> ), .B(n1274), .Y(n1823) );
  OAI21X1 U1832 ( .A(n160), .B(n1294), .C(n1823), .Y(n1878) );
  NAND2X1 U1833 ( .A(\mem<1><6> ), .B(n1274), .Y(n1824) );
  OAI21X1 U1834 ( .A(n160), .B(n1296), .C(n1824), .Y(n1877) );
  NAND2X1 U1835 ( .A(\mem<1><7> ), .B(n1274), .Y(n1825) );
  OAI21X1 U1836 ( .A(n160), .B(n1298), .C(n1825), .Y(n1876) );
  NAND2X1 U1837 ( .A(\mem<1><8> ), .B(n1275), .Y(n1826) );
  OAI21X1 U1838 ( .A(n160), .B(n1300), .C(n1826), .Y(n1875) );
  NAND2X1 U1839 ( .A(\mem<1><9> ), .B(n1275), .Y(n1827) );
  OAI21X1 U1840 ( .A(n160), .B(n1302), .C(n1827), .Y(n1874) );
  NAND2X1 U1841 ( .A(\mem<1><10> ), .B(n1275), .Y(n1828) );
  OAI21X1 U1842 ( .A(n160), .B(n1304), .C(n1828), .Y(n1873) );
  NAND2X1 U1843 ( .A(\mem<1><11> ), .B(n1275), .Y(n1829) );
  OAI21X1 U1844 ( .A(n160), .B(n1306), .C(n1829), .Y(n1872) );
  NAND2X1 U1845 ( .A(\mem<1><12> ), .B(n1275), .Y(n1830) );
  OAI21X1 U1846 ( .A(n160), .B(n1308), .C(n1830), .Y(n1871) );
  NAND2X1 U1847 ( .A(\mem<1><13> ), .B(n1275), .Y(n1831) );
  OAI21X1 U1848 ( .A(n160), .B(n1310), .C(n1831), .Y(n1870) );
  NAND2X1 U1849 ( .A(\mem<1><14> ), .B(n1275), .Y(n1832) );
  OAI21X1 U1850 ( .A(n160), .B(n1312), .C(n1832), .Y(n1869) );
  NAND2X1 U1851 ( .A(\mem<1><15> ), .B(n1275), .Y(n1833) );
  OAI21X1 U1852 ( .A(n160), .B(n1314), .C(n1833), .Y(n1868) );
  NAND2X1 U1853 ( .A(\mem<0><0> ), .B(n1277), .Y(n1836) );
  OAI21X1 U1854 ( .A(n1276), .B(n1285), .C(n1836), .Y(n1867) );
  NAND2X1 U1855 ( .A(\mem<0><1> ), .B(n1277), .Y(n1837) );
  OAI21X1 U1856 ( .A(n1276), .B(n1286), .C(n1837), .Y(n1866) );
  NAND2X1 U1857 ( .A(\mem<0><2> ), .B(n1277), .Y(n1838) );
  OAI21X1 U1858 ( .A(n1276), .B(n1288), .C(n1838), .Y(n1865) );
  NAND2X1 U1859 ( .A(\mem<0><3> ), .B(n1277), .Y(n1839) );
  OAI21X1 U1860 ( .A(n1276), .B(n1290), .C(n1839), .Y(n1864) );
  NAND2X1 U1861 ( .A(\mem<0><4> ), .B(n1277), .Y(n1840) );
  OAI21X1 U1862 ( .A(n1276), .B(n1292), .C(n1840), .Y(n1863) );
  NAND2X1 U1863 ( .A(\mem<0><5> ), .B(n1277), .Y(n1841) );
  OAI21X1 U1864 ( .A(n1276), .B(n1294), .C(n1841), .Y(n1862) );
  NAND2X1 U1865 ( .A(\mem<0><6> ), .B(n1277), .Y(n1842) );
  OAI21X1 U1866 ( .A(n1276), .B(n1296), .C(n1842), .Y(n1861) );
  NAND2X1 U1867 ( .A(\mem<0><7> ), .B(n1277), .Y(n1843) );
  OAI21X1 U1868 ( .A(n1276), .B(n1298), .C(n1843), .Y(n1860) );
  NAND2X1 U1869 ( .A(\mem<0><8> ), .B(n1278), .Y(n1844) );
  OAI21X1 U1870 ( .A(n1276), .B(n1300), .C(n1844), .Y(n1859) );
  NAND2X1 U1871 ( .A(\mem<0><9> ), .B(n1278), .Y(n1845) );
  OAI21X1 U1872 ( .A(n1276), .B(n1302), .C(n1845), .Y(n1858) );
  NAND2X1 U1873 ( .A(\mem<0><10> ), .B(n1278), .Y(n1846) );
  OAI21X1 U1874 ( .A(n1276), .B(n1304), .C(n1846), .Y(n1857) );
  NAND2X1 U1875 ( .A(\mem<0><11> ), .B(n1278), .Y(n1847) );
  OAI21X1 U1876 ( .A(n1276), .B(n1306), .C(n1847), .Y(n1856) );
  NAND2X1 U1877 ( .A(\mem<0><12> ), .B(n1278), .Y(n1848) );
  OAI21X1 U1878 ( .A(n1276), .B(n1308), .C(n1848), .Y(n1855) );
  NAND2X1 U1879 ( .A(\mem<0><13> ), .B(n1278), .Y(n1849) );
  OAI21X1 U1880 ( .A(n1276), .B(n1310), .C(n1849), .Y(n1854) );
  NAND2X1 U1881 ( .A(\mem<0><14> ), .B(n1278), .Y(n1850) );
  OAI21X1 U1882 ( .A(n1276), .B(n1312), .C(n1850), .Y(n1853) );
  NAND2X1 U1883 ( .A(\mem<0><15> ), .B(n1278), .Y(n1851) );
  OAI21X1 U1884 ( .A(n1276), .B(n1314), .C(n1851), .Y(n1852) );
endmodule


module memc_Size16_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<15> , \data_in<14> , \data_in<13> ,
         \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> ,
         \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> ,
         \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , write, clk,
         rst, createdump, \file_id<4> , \file_id<3> , \file_id<2> ,
         \file_id<1> , \file_id<0> ;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><15> , \mem<0><14> , \mem<0><13> ,
         \mem<0><12> , \mem<0><11> , \mem<0><10> , \mem<0><9> , \mem<0><8> ,
         \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> , \mem<0><3> ,
         \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><15> , \mem<1><14> ,
         \mem<1><13> , \mem<1><12> , \mem<1><11> , \mem<1><10> , \mem<1><9> ,
         \mem<1><8> , \mem<1><7> , \mem<1><6> , \mem<1><5> , \mem<1><4> ,
         \mem<1><3> , \mem<1><2> , \mem<1><1> , \mem<1><0> , \mem<2><15> ,
         \mem<2><14> , \mem<2><13> , \mem<2><12> , \mem<2><11> , \mem<2><10> ,
         \mem<2><9> , \mem<2><8> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><15> , \mem<3><14> , \mem<3><13> , \mem<3><12> , \mem<3><11> ,
         \mem<3><10> , \mem<3><9> , \mem<3><8> , \mem<3><7> , \mem<3><6> ,
         \mem<3><5> , \mem<3><4> , \mem<3><3> , \mem<3><2> , \mem<3><1> ,
         \mem<3><0> , \mem<4><15> , \mem<4><14> , \mem<4><13> , \mem<4><12> ,
         \mem<4><11> , \mem<4><10> , \mem<4><9> , \mem<4><8> , \mem<4><7> ,
         \mem<4><6> , \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><15> , \mem<5><14> , \mem<5><13> ,
         \mem<5><12> , \mem<5><11> , \mem<5><10> , \mem<5><9> , \mem<5><8> ,
         \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> , \mem<5><3> ,
         \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><15> , \mem<6><14> ,
         \mem<6><13> , \mem<6><12> , \mem<6><11> , \mem<6><10> , \mem<6><9> ,
         \mem<6><8> , \mem<6><7> , \mem<6><6> , \mem<6><5> , \mem<6><4> ,
         \mem<6><3> , \mem<6><2> , \mem<6><1> , \mem<6><0> , \mem<7><15> ,
         \mem<7><14> , \mem<7><13> , \mem<7><12> , \mem<7><11> , \mem<7><10> ,
         \mem<7><9> , \mem<7><8> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><15> , \mem<8><14> , \mem<8><13> , \mem<8><12> , \mem<8><11> ,
         \mem<8><10> , \mem<8><9> , \mem<8><8> , \mem<8><7> , \mem<8><6> ,
         \mem<8><5> , \mem<8><4> , \mem<8><3> , \mem<8><2> , \mem<8><1> ,
         \mem<8><0> , \mem<9><15> , \mem<9><14> , \mem<9><13> , \mem<9><12> ,
         \mem<9><11> , \mem<9><10> , \mem<9><9> , \mem<9><8> , \mem<9><7> ,
         \mem<9><6> , \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><15> , \mem<10><14> , \mem<10><13> ,
         \mem<10><12> , \mem<10><11> , \mem<10><10> , \mem<10><9> ,
         \mem<10><8> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><15> ,
         \mem<11><14> , \mem<11><13> , \mem<11><12> , \mem<11><11> ,
         \mem<11><10> , \mem<11><9> , \mem<11><8> , \mem<11><7> , \mem<11><6> ,
         \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> , \mem<11><1> ,
         \mem<11><0> , \mem<12><15> , \mem<12><14> , \mem<12><13> ,
         \mem<12><12> , \mem<12><11> , \mem<12><10> , \mem<12><9> ,
         \mem<12><8> , \mem<12><7> , \mem<12><6> , \mem<12><5> , \mem<12><4> ,
         \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> , \mem<13><15> ,
         \mem<13><14> , \mem<13><13> , \mem<13><12> , \mem<13><11> ,
         \mem<13><10> , \mem<13><9> , \mem<13><8> , \mem<13><7> , \mem<13><6> ,
         \mem<13><5> , \mem<13><4> , \mem<13><3> , \mem<13><2> , \mem<13><1> ,
         \mem<13><0> , \mem<14><15> , \mem<14><14> , \mem<14><13> ,
         \mem<14><12> , \mem<14><11> , \mem<14><10> , \mem<14><9> ,
         \mem<14><8> , \mem<14><7> , \mem<14><6> , \mem<14><5> , \mem<14><4> ,
         \mem<14><3> , \mem<14><2> , \mem<14><1> , \mem<14><0> , \mem<15><15> ,
         \mem<15><14> , \mem<15><13> , \mem<15><12> , \mem<15><11> ,
         \mem<15><10> , \mem<15><9> , \mem<15><8> , \mem<15><7> , \mem<15><6> ,
         \mem<15><5> , \mem<15><4> , \mem<15><3> , \mem<15><2> , \mem<15><1> ,
         \mem<15><0> , \mem<16><15> , \mem<16><14> , \mem<16><13> ,
         \mem<16><12> , \mem<16><11> , \mem<16><10> , \mem<16><9> ,
         \mem<16><8> , \mem<16><7> , \mem<16><6> , \mem<16><5> , \mem<16><4> ,
         \mem<16><3> , \mem<16><2> , \mem<16><1> , \mem<16><0> , \mem<17><15> ,
         \mem<17><14> , \mem<17><13> , \mem<17><12> , \mem<17><11> ,
         \mem<17><10> , \mem<17><9> , \mem<17><8> , \mem<17><7> , \mem<17><6> ,
         \mem<17><5> , \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> ,
         \mem<17><0> , \mem<18><15> , \mem<18><14> , \mem<18><13> ,
         \mem<18><12> , \mem<18><11> , \mem<18><10> , \mem<18><9> ,
         \mem<18><8> , \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> ,
         \mem<18><3> , \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><15> ,
         \mem<19><14> , \mem<19><13> , \mem<19><12> , \mem<19><11> ,
         \mem<19><10> , \mem<19><9> , \mem<19><8> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><15> , \mem<20><14> , \mem<20><13> ,
         \mem<20><12> , \mem<20><11> , \mem<20><10> , \mem<20><9> ,
         \mem<20><8> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><15> ,
         \mem<21><14> , \mem<21><13> , \mem<21><12> , \mem<21><11> ,
         \mem<21><10> , \mem<21><9> , \mem<21><8> , \mem<21><7> , \mem<21><6> ,
         \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> , \mem<21><1> ,
         \mem<21><0> , \mem<22><15> , \mem<22><14> , \mem<22><13> ,
         \mem<22><12> , \mem<22><11> , \mem<22><10> , \mem<22><9> ,
         \mem<22><8> , \mem<22><7> , \mem<22><6> , \mem<22><5> , \mem<22><4> ,
         \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> , \mem<23><15> ,
         \mem<23><14> , \mem<23><13> , \mem<23><12> , \mem<23><11> ,
         \mem<23><10> , \mem<23><9> , \mem<23><8> , \mem<23><7> , \mem<23><6> ,
         \mem<23><5> , \mem<23><4> , \mem<23><3> , \mem<23><2> , \mem<23><1> ,
         \mem<23><0> , \mem<24><15> , \mem<24><14> , \mem<24><13> ,
         \mem<24><12> , \mem<24><11> , \mem<24><10> , \mem<24><9> ,
         \mem<24><8> , \mem<24><7> , \mem<24><6> , \mem<24><5> , \mem<24><4> ,
         \mem<24><3> , \mem<24><2> , \mem<24><1> , \mem<24><0> , \mem<25><15> ,
         \mem<25><14> , \mem<25><13> , \mem<25><12> , \mem<25><11> ,
         \mem<25><10> , \mem<25><9> , \mem<25><8> , \mem<25><7> , \mem<25><6> ,
         \mem<25><5> , \mem<25><4> , \mem<25><3> , \mem<25><2> , \mem<25><1> ,
         \mem<25><0> , \mem<26><15> , \mem<26><14> , \mem<26><13> ,
         \mem<26><12> , \mem<26><11> , \mem<26><10> , \mem<26><9> ,
         \mem<26><8> , \mem<26><7> , \mem<26><6> , \mem<26><5> , \mem<26><4> ,
         \mem<26><3> , \mem<26><2> , \mem<26><1> , \mem<26><0> , \mem<27><15> ,
         \mem<27><14> , \mem<27><13> , \mem<27><12> , \mem<27><11> ,
         \mem<27><10> , \mem<27><9> , \mem<27><8> , \mem<27><7> , \mem<27><6> ,
         \mem<27><5> , \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> ,
         \mem<27><0> , \mem<28><15> , \mem<28><14> , \mem<28><13> ,
         \mem<28><12> , \mem<28><11> , \mem<28><10> , \mem<28><9> ,
         \mem<28><8> , \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> ,
         \mem<28><3> , \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><15> ,
         \mem<29><14> , \mem<29><13> , \mem<29><12> , \mem<29><11> ,
         \mem<29><10> , \mem<29><9> , \mem<29><8> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><15> , \mem<30><14> , \mem<30><13> ,
         \mem<30><12> , \mem<30><11> , \mem<30><10> , \mem<30><9> ,
         \mem<30><8> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><15> ,
         \mem<31><14> , \mem<31><13> , \mem<31><12> , \mem<31><11> ,
         \mem<31><10> , \mem<31><9> , \mem<31><8> , \mem<31><7> , \mem<31><6> ,
         \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> , \mem<31><1> ,
         \mem<31><0> , N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><15>  ( .D(n2152), .CLK(clk), .Q(\mem<0><15> ) );
  DFFPOSX1 \mem_reg<0><14>  ( .D(n2153), .CLK(clk), .Q(\mem<0><14> ) );
  DFFPOSX1 \mem_reg<0><13>  ( .D(n2154), .CLK(clk), .Q(\mem<0><13> ) );
  DFFPOSX1 \mem_reg<0><12>  ( .D(n2155), .CLK(clk), .Q(\mem<0><12> ) );
  DFFPOSX1 \mem_reg<0><11>  ( .D(n2156), .CLK(clk), .Q(\mem<0><11> ) );
  DFFPOSX1 \mem_reg<0><10>  ( .D(n2157), .CLK(clk), .Q(\mem<0><10> ) );
  DFFPOSX1 \mem_reg<0><9>  ( .D(n2158), .CLK(clk), .Q(\mem<0><9> ) );
  DFFPOSX1 \mem_reg<0><8>  ( .D(n2159), .CLK(clk), .Q(\mem<0><8> ) );
  DFFPOSX1 \mem_reg<0><7>  ( .D(n2160), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n2161), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n2162), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n2163), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n2164), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n2165), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n2166), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n2167), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><15>  ( .D(n2168), .CLK(clk), .Q(\mem<1><15> ) );
  DFFPOSX1 \mem_reg<1><14>  ( .D(n2169), .CLK(clk), .Q(\mem<1><14> ) );
  DFFPOSX1 \mem_reg<1><13>  ( .D(n2170), .CLK(clk), .Q(\mem<1><13> ) );
  DFFPOSX1 \mem_reg<1><12>  ( .D(n2171), .CLK(clk), .Q(\mem<1><12> ) );
  DFFPOSX1 \mem_reg<1><11>  ( .D(n2172), .CLK(clk), .Q(\mem<1><11> ) );
  DFFPOSX1 \mem_reg<1><10>  ( .D(n2173), .CLK(clk), .Q(\mem<1><10> ) );
  DFFPOSX1 \mem_reg<1><9>  ( .D(n2174), .CLK(clk), .Q(\mem<1><9> ) );
  DFFPOSX1 \mem_reg<1><8>  ( .D(n2175), .CLK(clk), .Q(\mem<1><8> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n2176), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n2177), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n2178), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n2179), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n2180), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n2181), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n2182), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n2183), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><15>  ( .D(n2184), .CLK(clk), .Q(\mem<2><15> ) );
  DFFPOSX1 \mem_reg<2><14>  ( .D(n2185), .CLK(clk), .Q(\mem<2><14> ) );
  DFFPOSX1 \mem_reg<2><13>  ( .D(n2186), .CLK(clk), .Q(\mem<2><13> ) );
  DFFPOSX1 \mem_reg<2><12>  ( .D(n2187), .CLK(clk), .Q(\mem<2><12> ) );
  DFFPOSX1 \mem_reg<2><11>  ( .D(n2188), .CLK(clk), .Q(\mem<2><11> ) );
  DFFPOSX1 \mem_reg<2><10>  ( .D(n2189), .CLK(clk), .Q(\mem<2><10> ) );
  DFFPOSX1 \mem_reg<2><9>  ( .D(n2190), .CLK(clk), .Q(\mem<2><9> ) );
  DFFPOSX1 \mem_reg<2><8>  ( .D(n2191), .CLK(clk), .Q(\mem<2><8> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n2192), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n2193), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n2194), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n2195), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n2196), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n2197), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n2198), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n2199), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><15>  ( .D(n2200), .CLK(clk), .Q(\mem<3><15> ) );
  DFFPOSX1 \mem_reg<3><14>  ( .D(n2201), .CLK(clk), .Q(\mem<3><14> ) );
  DFFPOSX1 \mem_reg<3><13>  ( .D(n2202), .CLK(clk), .Q(\mem<3><13> ) );
  DFFPOSX1 \mem_reg<3><12>  ( .D(n2203), .CLK(clk), .Q(\mem<3><12> ) );
  DFFPOSX1 \mem_reg<3><11>  ( .D(n2204), .CLK(clk), .Q(\mem<3><11> ) );
  DFFPOSX1 \mem_reg<3><10>  ( .D(n2205), .CLK(clk), .Q(\mem<3><10> ) );
  DFFPOSX1 \mem_reg<3><9>  ( .D(n2206), .CLK(clk), .Q(\mem<3><9> ) );
  DFFPOSX1 \mem_reg<3><8>  ( .D(n2207), .CLK(clk), .Q(\mem<3><8> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n2208), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n2209), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n2210), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n2211), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n2212), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n2213), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n2214), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n2215), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><15>  ( .D(n2216), .CLK(clk), .Q(\mem<4><15> ) );
  DFFPOSX1 \mem_reg<4><14>  ( .D(n2217), .CLK(clk), .Q(\mem<4><14> ) );
  DFFPOSX1 \mem_reg<4><13>  ( .D(n2218), .CLK(clk), .Q(\mem<4><13> ) );
  DFFPOSX1 \mem_reg<4><12>  ( .D(n2219), .CLK(clk), .Q(\mem<4><12> ) );
  DFFPOSX1 \mem_reg<4><11>  ( .D(n2220), .CLK(clk), .Q(\mem<4><11> ) );
  DFFPOSX1 \mem_reg<4><10>  ( .D(n2221), .CLK(clk), .Q(\mem<4><10> ) );
  DFFPOSX1 \mem_reg<4><9>  ( .D(n2222), .CLK(clk), .Q(\mem<4><9> ) );
  DFFPOSX1 \mem_reg<4><8>  ( .D(n2223), .CLK(clk), .Q(\mem<4><8> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n2224), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n2225), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n2226), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n2227), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n2228), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n2229), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n2230), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n2231), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><15>  ( .D(n2232), .CLK(clk), .Q(\mem<5><15> ) );
  DFFPOSX1 \mem_reg<5><14>  ( .D(n2233), .CLK(clk), .Q(\mem<5><14> ) );
  DFFPOSX1 \mem_reg<5><13>  ( .D(n2234), .CLK(clk), .Q(\mem<5><13> ) );
  DFFPOSX1 \mem_reg<5><12>  ( .D(n2235), .CLK(clk), .Q(\mem<5><12> ) );
  DFFPOSX1 \mem_reg<5><11>  ( .D(n2236), .CLK(clk), .Q(\mem<5><11> ) );
  DFFPOSX1 \mem_reg<5><10>  ( .D(n2237), .CLK(clk), .Q(\mem<5><10> ) );
  DFFPOSX1 \mem_reg<5><9>  ( .D(n2238), .CLK(clk), .Q(\mem<5><9> ) );
  DFFPOSX1 \mem_reg<5><8>  ( .D(n2239), .CLK(clk), .Q(\mem<5><8> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n2240), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n2241), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n2242), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n2243), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n2244), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n2245), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n2246), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n2247), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><15>  ( .D(n2248), .CLK(clk), .Q(\mem<6><15> ) );
  DFFPOSX1 \mem_reg<6><14>  ( .D(n2249), .CLK(clk), .Q(\mem<6><14> ) );
  DFFPOSX1 \mem_reg<6><13>  ( .D(n2250), .CLK(clk), .Q(\mem<6><13> ) );
  DFFPOSX1 \mem_reg<6><12>  ( .D(n2251), .CLK(clk), .Q(\mem<6><12> ) );
  DFFPOSX1 \mem_reg<6><11>  ( .D(n2252), .CLK(clk), .Q(\mem<6><11> ) );
  DFFPOSX1 \mem_reg<6><10>  ( .D(n2253), .CLK(clk), .Q(\mem<6><10> ) );
  DFFPOSX1 \mem_reg<6><9>  ( .D(n2254), .CLK(clk), .Q(\mem<6><9> ) );
  DFFPOSX1 \mem_reg<6><8>  ( .D(n2255), .CLK(clk), .Q(\mem<6><8> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n2256), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n2257), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n2258), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n2259), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n2260), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n2261), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n2262), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n2263), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><15>  ( .D(n2264), .CLK(clk), .Q(\mem<7><15> ) );
  DFFPOSX1 \mem_reg<7><14>  ( .D(n2265), .CLK(clk), .Q(\mem<7><14> ) );
  DFFPOSX1 \mem_reg<7><13>  ( .D(n2266), .CLK(clk), .Q(\mem<7><13> ) );
  DFFPOSX1 \mem_reg<7><12>  ( .D(n2267), .CLK(clk), .Q(\mem<7><12> ) );
  DFFPOSX1 \mem_reg<7><11>  ( .D(n2268), .CLK(clk), .Q(\mem<7><11> ) );
  DFFPOSX1 \mem_reg<7><10>  ( .D(n2269), .CLK(clk), .Q(\mem<7><10> ) );
  DFFPOSX1 \mem_reg<7><9>  ( .D(n2270), .CLK(clk), .Q(\mem<7><9> ) );
  DFFPOSX1 \mem_reg<7><8>  ( .D(n2271), .CLK(clk), .Q(\mem<7><8> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n2272), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n2273), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n2274), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n2275), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n2276), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n2277), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n2278), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n2279), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><15>  ( .D(n2280), .CLK(clk), .Q(\mem<8><15> ) );
  DFFPOSX1 \mem_reg<8><14>  ( .D(n2281), .CLK(clk), .Q(\mem<8><14> ) );
  DFFPOSX1 \mem_reg<8><13>  ( .D(n2282), .CLK(clk), .Q(\mem<8><13> ) );
  DFFPOSX1 \mem_reg<8><12>  ( .D(n2283), .CLK(clk), .Q(\mem<8><12> ) );
  DFFPOSX1 \mem_reg<8><11>  ( .D(n2284), .CLK(clk), .Q(\mem<8><11> ) );
  DFFPOSX1 \mem_reg<8><10>  ( .D(n2285), .CLK(clk), .Q(\mem<8><10> ) );
  DFFPOSX1 \mem_reg<8><9>  ( .D(n2286), .CLK(clk), .Q(\mem<8><9> ) );
  DFFPOSX1 \mem_reg<8><8>  ( .D(n2287), .CLK(clk), .Q(\mem<8><8> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n2288), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n2289), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n2290), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n2291), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n2292), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n2293), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n2294), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n2295), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><15>  ( .D(n2296), .CLK(clk), .Q(\mem<9><15> ) );
  DFFPOSX1 \mem_reg<9><14>  ( .D(n2297), .CLK(clk), .Q(\mem<9><14> ) );
  DFFPOSX1 \mem_reg<9><13>  ( .D(n2298), .CLK(clk), .Q(\mem<9><13> ) );
  DFFPOSX1 \mem_reg<9><12>  ( .D(n2299), .CLK(clk), .Q(\mem<9><12> ) );
  DFFPOSX1 \mem_reg<9><11>  ( .D(n2300), .CLK(clk), .Q(\mem<9><11> ) );
  DFFPOSX1 \mem_reg<9><10>  ( .D(n2301), .CLK(clk), .Q(\mem<9><10> ) );
  DFFPOSX1 \mem_reg<9><9>  ( .D(n2302), .CLK(clk), .Q(\mem<9><9> ) );
  DFFPOSX1 \mem_reg<9><8>  ( .D(n2303), .CLK(clk), .Q(\mem<9><8> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n2304), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n2305), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n2306), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n2307), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n2308), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n2309), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n2310), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n2311), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><15>  ( .D(n2312), .CLK(clk), .Q(\mem<10><15> ) );
  DFFPOSX1 \mem_reg<10><14>  ( .D(n2313), .CLK(clk), .Q(\mem<10><14> ) );
  DFFPOSX1 \mem_reg<10><13>  ( .D(n2314), .CLK(clk), .Q(\mem<10><13> ) );
  DFFPOSX1 \mem_reg<10><12>  ( .D(n2315), .CLK(clk), .Q(\mem<10><12> ) );
  DFFPOSX1 \mem_reg<10><11>  ( .D(n2316), .CLK(clk), .Q(\mem<10><11> ) );
  DFFPOSX1 \mem_reg<10><10>  ( .D(n2317), .CLK(clk), .Q(\mem<10><10> ) );
  DFFPOSX1 \mem_reg<10><9>  ( .D(n2318), .CLK(clk), .Q(\mem<10><9> ) );
  DFFPOSX1 \mem_reg<10><8>  ( .D(n2319), .CLK(clk), .Q(\mem<10><8> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n2320), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n2321), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n2322), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n2323), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n2324), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n2325), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n2326), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n2327), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><15>  ( .D(n2328), .CLK(clk), .Q(\mem<11><15> ) );
  DFFPOSX1 \mem_reg<11><14>  ( .D(n2329), .CLK(clk), .Q(\mem<11><14> ) );
  DFFPOSX1 \mem_reg<11><13>  ( .D(n2330), .CLK(clk), .Q(\mem<11><13> ) );
  DFFPOSX1 \mem_reg<11><12>  ( .D(n2331), .CLK(clk), .Q(\mem<11><12> ) );
  DFFPOSX1 \mem_reg<11><11>  ( .D(n2332), .CLK(clk), .Q(\mem<11><11> ) );
  DFFPOSX1 \mem_reg<11><10>  ( .D(n2333), .CLK(clk), .Q(\mem<11><10> ) );
  DFFPOSX1 \mem_reg<11><9>  ( .D(n2334), .CLK(clk), .Q(\mem<11><9> ) );
  DFFPOSX1 \mem_reg<11><8>  ( .D(n2335), .CLK(clk), .Q(\mem<11><8> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n2336), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n2337), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n2338), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n2339), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n2340), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n2341), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n2342), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n2343), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><15>  ( .D(n2344), .CLK(clk), .Q(\mem<12><15> ) );
  DFFPOSX1 \mem_reg<12><14>  ( .D(n2345), .CLK(clk), .Q(\mem<12><14> ) );
  DFFPOSX1 \mem_reg<12><13>  ( .D(n2346), .CLK(clk), .Q(\mem<12><13> ) );
  DFFPOSX1 \mem_reg<12><12>  ( .D(n2347), .CLK(clk), .Q(\mem<12><12> ) );
  DFFPOSX1 \mem_reg<12><11>  ( .D(n2348), .CLK(clk), .Q(\mem<12><11> ) );
  DFFPOSX1 \mem_reg<12><10>  ( .D(n2349), .CLK(clk), .Q(\mem<12><10> ) );
  DFFPOSX1 \mem_reg<12><9>  ( .D(n2350), .CLK(clk), .Q(\mem<12><9> ) );
  DFFPOSX1 \mem_reg<12><8>  ( .D(n2351), .CLK(clk), .Q(\mem<12><8> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n2352), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n2353), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n2354), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n2355), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n2356), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n2357), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n2358), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n2359), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><15>  ( .D(n2360), .CLK(clk), .Q(\mem<13><15> ) );
  DFFPOSX1 \mem_reg<13><14>  ( .D(n2361), .CLK(clk), .Q(\mem<13><14> ) );
  DFFPOSX1 \mem_reg<13><13>  ( .D(n2362), .CLK(clk), .Q(\mem<13><13> ) );
  DFFPOSX1 \mem_reg<13><12>  ( .D(n2363), .CLK(clk), .Q(\mem<13><12> ) );
  DFFPOSX1 \mem_reg<13><11>  ( .D(n2364), .CLK(clk), .Q(\mem<13><11> ) );
  DFFPOSX1 \mem_reg<13><10>  ( .D(n2365), .CLK(clk), .Q(\mem<13><10> ) );
  DFFPOSX1 \mem_reg<13><9>  ( .D(n2366), .CLK(clk), .Q(\mem<13><9> ) );
  DFFPOSX1 \mem_reg<13><8>  ( .D(n2367), .CLK(clk), .Q(\mem<13><8> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n2368), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n2369), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n2370), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n2371), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n2372), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n2373), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n2374), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n2375), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><15>  ( .D(n2376), .CLK(clk), .Q(\mem<14><15> ) );
  DFFPOSX1 \mem_reg<14><14>  ( .D(n2377), .CLK(clk), .Q(\mem<14><14> ) );
  DFFPOSX1 \mem_reg<14><13>  ( .D(n2378), .CLK(clk), .Q(\mem<14><13> ) );
  DFFPOSX1 \mem_reg<14><12>  ( .D(n2379), .CLK(clk), .Q(\mem<14><12> ) );
  DFFPOSX1 \mem_reg<14><11>  ( .D(n2380), .CLK(clk), .Q(\mem<14><11> ) );
  DFFPOSX1 \mem_reg<14><10>  ( .D(n2381), .CLK(clk), .Q(\mem<14><10> ) );
  DFFPOSX1 \mem_reg<14><9>  ( .D(n2382), .CLK(clk), .Q(\mem<14><9> ) );
  DFFPOSX1 \mem_reg<14><8>  ( .D(n2383), .CLK(clk), .Q(\mem<14><8> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n2384), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n2385), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n2386), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n2387), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n2388), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n2389), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n2390), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n2391), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><15>  ( .D(n2392), .CLK(clk), .Q(\mem<15><15> ) );
  DFFPOSX1 \mem_reg<15><14>  ( .D(n2393), .CLK(clk), .Q(\mem<15><14> ) );
  DFFPOSX1 \mem_reg<15><13>  ( .D(n2394), .CLK(clk), .Q(\mem<15><13> ) );
  DFFPOSX1 \mem_reg<15><12>  ( .D(n2395), .CLK(clk), .Q(\mem<15><12> ) );
  DFFPOSX1 \mem_reg<15><11>  ( .D(n2396), .CLK(clk), .Q(\mem<15><11> ) );
  DFFPOSX1 \mem_reg<15><10>  ( .D(n2397), .CLK(clk), .Q(\mem<15><10> ) );
  DFFPOSX1 \mem_reg<15><9>  ( .D(n2398), .CLK(clk), .Q(\mem<15><9> ) );
  DFFPOSX1 \mem_reg<15><8>  ( .D(n2399), .CLK(clk), .Q(\mem<15><8> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n2400), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n2401), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n2402), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n2403), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n2404), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n2405), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n2406), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n2407), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><15>  ( .D(n2408), .CLK(clk), .Q(\mem<16><15> ) );
  DFFPOSX1 \mem_reg<16><14>  ( .D(n2409), .CLK(clk), .Q(\mem<16><14> ) );
  DFFPOSX1 \mem_reg<16><13>  ( .D(n2410), .CLK(clk), .Q(\mem<16><13> ) );
  DFFPOSX1 \mem_reg<16><12>  ( .D(n2411), .CLK(clk), .Q(\mem<16><12> ) );
  DFFPOSX1 \mem_reg<16><11>  ( .D(n2412), .CLK(clk), .Q(\mem<16><11> ) );
  DFFPOSX1 \mem_reg<16><10>  ( .D(n2413), .CLK(clk), .Q(\mem<16><10> ) );
  DFFPOSX1 \mem_reg<16><9>  ( .D(n2414), .CLK(clk), .Q(\mem<16><9> ) );
  DFFPOSX1 \mem_reg<16><8>  ( .D(n2415), .CLK(clk), .Q(\mem<16><8> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n2416), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n2417), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n2418), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n2419), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n2420), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n2421), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n2422), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n2423), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><15>  ( .D(n2424), .CLK(clk), .Q(\mem<17><15> ) );
  DFFPOSX1 \mem_reg<17><14>  ( .D(n2425), .CLK(clk), .Q(\mem<17><14> ) );
  DFFPOSX1 \mem_reg<17><13>  ( .D(n2426), .CLK(clk), .Q(\mem<17><13> ) );
  DFFPOSX1 \mem_reg<17><12>  ( .D(n2427), .CLK(clk), .Q(\mem<17><12> ) );
  DFFPOSX1 \mem_reg<17><11>  ( .D(n2428), .CLK(clk), .Q(\mem<17><11> ) );
  DFFPOSX1 \mem_reg<17><10>  ( .D(n2429), .CLK(clk), .Q(\mem<17><10> ) );
  DFFPOSX1 \mem_reg<17><9>  ( .D(n2430), .CLK(clk), .Q(\mem<17><9> ) );
  DFFPOSX1 \mem_reg<17><8>  ( .D(n2431), .CLK(clk), .Q(\mem<17><8> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n2432), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n2433), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n2434), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n2435), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n2436), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n2437), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n2438), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n2439), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><15>  ( .D(n2440), .CLK(clk), .Q(\mem<18><15> ) );
  DFFPOSX1 \mem_reg<18><14>  ( .D(n2441), .CLK(clk), .Q(\mem<18><14> ) );
  DFFPOSX1 \mem_reg<18><13>  ( .D(n2442), .CLK(clk), .Q(\mem<18><13> ) );
  DFFPOSX1 \mem_reg<18><12>  ( .D(n2443), .CLK(clk), .Q(\mem<18><12> ) );
  DFFPOSX1 \mem_reg<18><11>  ( .D(n2444), .CLK(clk), .Q(\mem<18><11> ) );
  DFFPOSX1 \mem_reg<18><10>  ( .D(n2445), .CLK(clk), .Q(\mem<18><10> ) );
  DFFPOSX1 \mem_reg<18><9>  ( .D(n2446), .CLK(clk), .Q(\mem<18><9> ) );
  DFFPOSX1 \mem_reg<18><8>  ( .D(n2447), .CLK(clk), .Q(\mem<18><8> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n2448), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n2449), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n2450), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n2451), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n2452), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n2453), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n2454), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n2455), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><15>  ( .D(n2456), .CLK(clk), .Q(\mem<19><15> ) );
  DFFPOSX1 \mem_reg<19><14>  ( .D(n2457), .CLK(clk), .Q(\mem<19><14> ) );
  DFFPOSX1 \mem_reg<19><13>  ( .D(n2458), .CLK(clk), .Q(\mem<19><13> ) );
  DFFPOSX1 \mem_reg<19><12>  ( .D(n2459), .CLK(clk), .Q(\mem<19><12> ) );
  DFFPOSX1 \mem_reg<19><11>  ( .D(n2460), .CLK(clk), .Q(\mem<19><11> ) );
  DFFPOSX1 \mem_reg<19><10>  ( .D(n2461), .CLK(clk), .Q(\mem<19><10> ) );
  DFFPOSX1 \mem_reg<19><9>  ( .D(n2462), .CLK(clk), .Q(\mem<19><9> ) );
  DFFPOSX1 \mem_reg<19><8>  ( .D(n2463), .CLK(clk), .Q(\mem<19><8> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n2464), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n2465), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n2466), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n2467), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n2468), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n2469), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n2470), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n2471), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><15>  ( .D(n2472), .CLK(clk), .Q(\mem<20><15> ) );
  DFFPOSX1 \mem_reg<20><14>  ( .D(n2473), .CLK(clk), .Q(\mem<20><14> ) );
  DFFPOSX1 \mem_reg<20><13>  ( .D(n2474), .CLK(clk), .Q(\mem<20><13> ) );
  DFFPOSX1 \mem_reg<20><12>  ( .D(n2475), .CLK(clk), .Q(\mem<20><12> ) );
  DFFPOSX1 \mem_reg<20><11>  ( .D(n2476), .CLK(clk), .Q(\mem<20><11> ) );
  DFFPOSX1 \mem_reg<20><10>  ( .D(n2477), .CLK(clk), .Q(\mem<20><10> ) );
  DFFPOSX1 \mem_reg<20><9>  ( .D(n2478), .CLK(clk), .Q(\mem<20><9> ) );
  DFFPOSX1 \mem_reg<20><8>  ( .D(n2479), .CLK(clk), .Q(\mem<20><8> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n2480), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n2481), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n2482), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n2483), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n2484), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n2485), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n2486), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n2487), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><15>  ( .D(n2488), .CLK(clk), .Q(\mem<21><15> ) );
  DFFPOSX1 \mem_reg<21><14>  ( .D(n2489), .CLK(clk), .Q(\mem<21><14> ) );
  DFFPOSX1 \mem_reg<21><13>  ( .D(n2490), .CLK(clk), .Q(\mem<21><13> ) );
  DFFPOSX1 \mem_reg<21><12>  ( .D(n2491), .CLK(clk), .Q(\mem<21><12> ) );
  DFFPOSX1 \mem_reg<21><11>  ( .D(n2492), .CLK(clk), .Q(\mem<21><11> ) );
  DFFPOSX1 \mem_reg<21><10>  ( .D(n2493), .CLK(clk), .Q(\mem<21><10> ) );
  DFFPOSX1 \mem_reg<21><9>  ( .D(n2494), .CLK(clk), .Q(\mem<21><9> ) );
  DFFPOSX1 \mem_reg<21><8>  ( .D(n2495), .CLK(clk), .Q(\mem<21><8> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n2496), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n2497), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n2498), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n2499), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n2500), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n2501), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n2502), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n2503), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><15>  ( .D(n2504), .CLK(clk), .Q(\mem<22><15> ) );
  DFFPOSX1 \mem_reg<22><14>  ( .D(n2505), .CLK(clk), .Q(\mem<22><14> ) );
  DFFPOSX1 \mem_reg<22><13>  ( .D(n2506), .CLK(clk), .Q(\mem<22><13> ) );
  DFFPOSX1 \mem_reg<22><12>  ( .D(n2507), .CLK(clk), .Q(\mem<22><12> ) );
  DFFPOSX1 \mem_reg<22><11>  ( .D(n2508), .CLK(clk), .Q(\mem<22><11> ) );
  DFFPOSX1 \mem_reg<22><10>  ( .D(n2509), .CLK(clk), .Q(\mem<22><10> ) );
  DFFPOSX1 \mem_reg<22><9>  ( .D(n2510), .CLK(clk), .Q(\mem<22><9> ) );
  DFFPOSX1 \mem_reg<22><8>  ( .D(n2511), .CLK(clk), .Q(\mem<22><8> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n2512), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n2513), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n2514), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n2515), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n2516), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n2517), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n2518), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n2519), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><15>  ( .D(n2520), .CLK(clk), .Q(\mem<23><15> ) );
  DFFPOSX1 \mem_reg<23><14>  ( .D(n2521), .CLK(clk), .Q(\mem<23><14> ) );
  DFFPOSX1 \mem_reg<23><13>  ( .D(n2522), .CLK(clk), .Q(\mem<23><13> ) );
  DFFPOSX1 \mem_reg<23><12>  ( .D(n2523), .CLK(clk), .Q(\mem<23><12> ) );
  DFFPOSX1 \mem_reg<23><11>  ( .D(n2524), .CLK(clk), .Q(\mem<23><11> ) );
  DFFPOSX1 \mem_reg<23><10>  ( .D(n2525), .CLK(clk), .Q(\mem<23><10> ) );
  DFFPOSX1 \mem_reg<23><9>  ( .D(n2526), .CLK(clk), .Q(\mem<23><9> ) );
  DFFPOSX1 \mem_reg<23><8>  ( .D(n2527), .CLK(clk), .Q(\mem<23><8> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n2528), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n2529), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n2530), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n2531), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n2532), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n2533), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n2534), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n2535), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><15>  ( .D(n2536), .CLK(clk), .Q(\mem<24><15> ) );
  DFFPOSX1 \mem_reg<24><14>  ( .D(n2537), .CLK(clk), .Q(\mem<24><14> ) );
  DFFPOSX1 \mem_reg<24><13>  ( .D(n2538), .CLK(clk), .Q(\mem<24><13> ) );
  DFFPOSX1 \mem_reg<24><12>  ( .D(n2539), .CLK(clk), .Q(\mem<24><12> ) );
  DFFPOSX1 \mem_reg<24><11>  ( .D(n2540), .CLK(clk), .Q(\mem<24><11> ) );
  DFFPOSX1 \mem_reg<24><10>  ( .D(n2541), .CLK(clk), .Q(\mem<24><10> ) );
  DFFPOSX1 \mem_reg<24><9>  ( .D(n2542), .CLK(clk), .Q(\mem<24><9> ) );
  DFFPOSX1 \mem_reg<24><8>  ( .D(n2543), .CLK(clk), .Q(\mem<24><8> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n2544), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n2545), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n2546), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n2547), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n2548), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n2549), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n2550), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n2551), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><15>  ( .D(n2552), .CLK(clk), .Q(\mem<25><15> ) );
  DFFPOSX1 \mem_reg<25><14>  ( .D(n2553), .CLK(clk), .Q(\mem<25><14> ) );
  DFFPOSX1 \mem_reg<25><13>  ( .D(n2554), .CLK(clk), .Q(\mem<25><13> ) );
  DFFPOSX1 \mem_reg<25><12>  ( .D(n2555), .CLK(clk), .Q(\mem<25><12> ) );
  DFFPOSX1 \mem_reg<25><11>  ( .D(n2556), .CLK(clk), .Q(\mem<25><11> ) );
  DFFPOSX1 \mem_reg<25><10>  ( .D(n2557), .CLK(clk), .Q(\mem<25><10> ) );
  DFFPOSX1 \mem_reg<25><9>  ( .D(n2558), .CLK(clk), .Q(\mem<25><9> ) );
  DFFPOSX1 \mem_reg<25><8>  ( .D(n2559), .CLK(clk), .Q(\mem<25><8> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n2560), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n2561), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n2562), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n2563), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n2564), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n2565), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n2566), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n2567), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><15>  ( .D(n2568), .CLK(clk), .Q(\mem<26><15> ) );
  DFFPOSX1 \mem_reg<26><14>  ( .D(n2569), .CLK(clk), .Q(\mem<26><14> ) );
  DFFPOSX1 \mem_reg<26><13>  ( .D(n2570), .CLK(clk), .Q(\mem<26><13> ) );
  DFFPOSX1 \mem_reg<26><12>  ( .D(n2571), .CLK(clk), .Q(\mem<26><12> ) );
  DFFPOSX1 \mem_reg<26><11>  ( .D(n2572), .CLK(clk), .Q(\mem<26><11> ) );
  DFFPOSX1 \mem_reg<26><10>  ( .D(n2573), .CLK(clk), .Q(\mem<26><10> ) );
  DFFPOSX1 \mem_reg<26><9>  ( .D(n2574), .CLK(clk), .Q(\mem<26><9> ) );
  DFFPOSX1 \mem_reg<26><8>  ( .D(n2575), .CLK(clk), .Q(\mem<26><8> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n2576), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n2577), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n2578), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n2579), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n2580), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n2581), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n2582), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n2583), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><15>  ( .D(n2584), .CLK(clk), .Q(\mem<27><15> ) );
  DFFPOSX1 \mem_reg<27><14>  ( .D(n2585), .CLK(clk), .Q(\mem<27><14> ) );
  DFFPOSX1 \mem_reg<27><13>  ( .D(n2586), .CLK(clk), .Q(\mem<27><13> ) );
  DFFPOSX1 \mem_reg<27><12>  ( .D(n2587), .CLK(clk), .Q(\mem<27><12> ) );
  DFFPOSX1 \mem_reg<27><11>  ( .D(n2588), .CLK(clk), .Q(\mem<27><11> ) );
  DFFPOSX1 \mem_reg<27><10>  ( .D(n2589), .CLK(clk), .Q(\mem<27><10> ) );
  DFFPOSX1 \mem_reg<27><9>  ( .D(n2590), .CLK(clk), .Q(\mem<27><9> ) );
  DFFPOSX1 \mem_reg<27><8>  ( .D(n2591), .CLK(clk), .Q(\mem<27><8> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n2592), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n2593), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n2594), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n2595), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n2596), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n2597), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n2598), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n2599), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><15>  ( .D(n2600), .CLK(clk), .Q(\mem<28><15> ) );
  DFFPOSX1 \mem_reg<28><14>  ( .D(n2601), .CLK(clk), .Q(\mem<28><14> ) );
  DFFPOSX1 \mem_reg<28><13>  ( .D(n2602), .CLK(clk), .Q(\mem<28><13> ) );
  DFFPOSX1 \mem_reg<28><12>  ( .D(n2603), .CLK(clk), .Q(\mem<28><12> ) );
  DFFPOSX1 \mem_reg<28><11>  ( .D(n2604), .CLK(clk), .Q(\mem<28><11> ) );
  DFFPOSX1 \mem_reg<28><10>  ( .D(n2605), .CLK(clk), .Q(\mem<28><10> ) );
  DFFPOSX1 \mem_reg<28><9>  ( .D(n2606), .CLK(clk), .Q(\mem<28><9> ) );
  DFFPOSX1 \mem_reg<28><8>  ( .D(n2607), .CLK(clk), .Q(\mem<28><8> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n2608), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n2609), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n2610), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n2611), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n2612), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n2613), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n2614), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n2615), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><15>  ( .D(n2616), .CLK(clk), .Q(\mem<29><15> ) );
  DFFPOSX1 \mem_reg<29><14>  ( .D(n2617), .CLK(clk), .Q(\mem<29><14> ) );
  DFFPOSX1 \mem_reg<29><13>  ( .D(n2618), .CLK(clk), .Q(\mem<29><13> ) );
  DFFPOSX1 \mem_reg<29><12>  ( .D(n2619), .CLK(clk), .Q(\mem<29><12> ) );
  DFFPOSX1 \mem_reg<29><11>  ( .D(n2620), .CLK(clk), .Q(\mem<29><11> ) );
  DFFPOSX1 \mem_reg<29><10>  ( .D(n2621), .CLK(clk), .Q(\mem<29><10> ) );
  DFFPOSX1 \mem_reg<29><9>  ( .D(n2622), .CLK(clk), .Q(\mem<29><9> ) );
  DFFPOSX1 \mem_reg<29><8>  ( .D(n2623), .CLK(clk), .Q(\mem<29><8> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n2624), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n2625), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n2626), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n2627), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n2628), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n2629), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n2630), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n2631), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><15>  ( .D(n2632), .CLK(clk), .Q(\mem<30><15> ) );
  DFFPOSX1 \mem_reg<30><14>  ( .D(n2633), .CLK(clk), .Q(\mem<30><14> ) );
  DFFPOSX1 \mem_reg<30><13>  ( .D(n2634), .CLK(clk), .Q(\mem<30><13> ) );
  DFFPOSX1 \mem_reg<30><12>  ( .D(n2635), .CLK(clk), .Q(\mem<30><12> ) );
  DFFPOSX1 \mem_reg<30><11>  ( .D(n2636), .CLK(clk), .Q(\mem<30><11> ) );
  DFFPOSX1 \mem_reg<30><10>  ( .D(n2637), .CLK(clk), .Q(\mem<30><10> ) );
  DFFPOSX1 \mem_reg<30><9>  ( .D(n2638), .CLK(clk), .Q(\mem<30><9> ) );
  DFFPOSX1 \mem_reg<30><8>  ( .D(n2639), .CLK(clk), .Q(\mem<30><8> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n2640), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n2641), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n2642), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n2643), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n2644), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n2645), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n2646), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n2647), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><15>  ( .D(n2648), .CLK(clk), .Q(\mem<31><15> ) );
  DFFPOSX1 \mem_reg<31><14>  ( .D(n2649), .CLK(clk), .Q(\mem<31><14> ) );
  DFFPOSX1 \mem_reg<31><13>  ( .D(n2650), .CLK(clk), .Q(\mem<31><13> ) );
  DFFPOSX1 \mem_reg<31><12>  ( .D(n2651), .CLK(clk), .Q(\mem<31><12> ) );
  DFFPOSX1 \mem_reg<31><11>  ( .D(n2652), .CLK(clk), .Q(\mem<31><11> ) );
  DFFPOSX1 \mem_reg<31><10>  ( .D(n2653), .CLK(clk), .Q(\mem<31><10> ) );
  DFFPOSX1 \mem_reg<31><9>  ( .D(n2654), .CLK(clk), .Q(\mem<31><9> ) );
  DFFPOSX1 \mem_reg<31><8>  ( .D(n2655), .CLK(clk), .Q(\mem<31><8> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n2656), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n2657), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n2658), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n2659), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n2660), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n2661), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n2662), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n2663), .CLK(clk), .Q(\mem<31><0> ) );
  NOR3X1 U1176 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n2664) );
  INVX2 U2 ( .A(n1839), .Y(n1847) );
  INVX2 U3 ( .A(n1839), .Y(n1845) );
  INVX2 U4 ( .A(n1839), .Y(n1846) );
  INVX1 U5 ( .A(n1838), .Y(n1852) );
  INVX1 U6 ( .A(n1837), .Y(n1854) );
  INVX1 U7 ( .A(n1837), .Y(n1853) );
  INVX4 U8 ( .A(n21), .Y(n1247) );
  INVX4 U9 ( .A(n5), .Y(n1244) );
  INVX1 U10 ( .A(n1856), .Y(n1839) );
  INVX1 U11 ( .A(n1855), .Y(n1837) );
  INVX1 U12 ( .A(n1856), .Y(n1838) );
  INVX1 U13 ( .A(n1824), .Y(n1825) );
  INVX1 U14 ( .A(n1824), .Y(n1826) );
  INVX1 U15 ( .A(n1824), .Y(n1827) );
  INVX1 U16 ( .A(n1823), .Y(n1828) );
  INVX2 U17 ( .A(n1839), .Y(n1848) );
  INVX1 U18 ( .A(n1823), .Y(n1829) );
  INVX2 U19 ( .A(n1839), .Y(n1849) );
  INVX1 U20 ( .A(n1823), .Y(n1830) );
  INVX1 U21 ( .A(n1836), .Y(n1831) );
  INVX1 U22 ( .A(n1836), .Y(n1832) );
  INVX1 U23 ( .A(n1836), .Y(n1833) );
  INVX2 U24 ( .A(n1823), .Y(n1834) );
  INVX2 U25 ( .A(n1824), .Y(n1835) );
  INVX1 U26 ( .A(n1800), .Y(N32) );
  INVX1 U27 ( .A(n1801), .Y(N31) );
  INVX1 U28 ( .A(n1802), .Y(N30) );
  INVX1 U29 ( .A(n1803), .Y(N29) );
  INVX1 U30 ( .A(n1804), .Y(N28) );
  INVX1 U31 ( .A(n1805), .Y(N27) );
  INVX1 U32 ( .A(n1806), .Y(N26) );
  INVX1 U33 ( .A(n1807), .Y(N25) );
  INVX1 U34 ( .A(n1808), .Y(N24) );
  INVX1 U35 ( .A(n1809), .Y(N23) );
  INVX1 U36 ( .A(n1810), .Y(N22) );
  INVX1 U37 ( .A(n1811), .Y(N21) );
  INVX1 U38 ( .A(n1812), .Y(N20) );
  INVX1 U39 ( .A(n1813), .Y(N19) );
  INVX1 U40 ( .A(n1814), .Y(N18) );
  INVX1 U41 ( .A(n1815), .Y(N17) );
  INVX2 U42 ( .A(n1942), .Y(n1822) );
  INVX1 U43 ( .A(N13), .Y(n1943) );
  INVX1 U44 ( .A(n1943), .Y(n1817) );
  INVX1 U45 ( .A(n1943), .Y(n1818) );
  INVX1 U46 ( .A(n1939), .Y(n1836) );
  INVX1 U47 ( .A(n1942), .Y(n1821) );
  INVX1 U48 ( .A(n1942), .Y(n1819) );
  INVX1 U49 ( .A(n1942), .Y(n1820) );
  INVX1 U50 ( .A(n1938), .Y(n1855) );
  INVX2 U51 ( .A(n1838), .Y(n1851) );
  INVX1 U52 ( .A(n1944), .Y(n1816) );
  INVX1 U53 ( .A(n1855), .Y(n1840) );
  INVX1 U54 ( .A(rst), .Y(n1937) );
  INVX1 U55 ( .A(n1939), .Y(n1824) );
  INVX1 U56 ( .A(n1939), .Y(n1823) );
  INVX1 U57 ( .A(n1238), .Y(n1857) );
  INVX1 U58 ( .A(n1239), .Y(n1864) );
  INVX1 U59 ( .A(n1240), .Y(n1881) );
  INVX1 U60 ( .A(n1241), .Y(n1898) );
  INVX4 U61 ( .A(n1), .Y(n2) );
  OR2X2 U62 ( .A(write), .B(rst), .Y(n1) );
  AND2X2 U63 ( .A(write), .B(n1937), .Y(n3) );
  AND2X2 U64 ( .A(\data_in<0> ), .B(n1903), .Y(n4) );
  AND2X2 U65 ( .A(n1903), .B(n1242), .Y(n5) );
  AND2X2 U66 ( .A(\data_in<1> ), .B(n1903), .Y(n6) );
  AND2X2 U67 ( .A(\data_in<2> ), .B(n1903), .Y(n7) );
  AND2X2 U68 ( .A(\data_in<3> ), .B(n1903), .Y(n8) );
  AND2X2 U69 ( .A(\data_in<4> ), .B(n1903), .Y(n9) );
  AND2X2 U70 ( .A(\data_in<5> ), .B(n1903), .Y(n10) );
  AND2X2 U71 ( .A(\data_in<6> ), .B(n1903), .Y(n11) );
  AND2X2 U72 ( .A(\data_in<7> ), .B(n1903), .Y(n12) );
  AND2X2 U73 ( .A(\data_in<8> ), .B(n1903), .Y(n13) );
  AND2X2 U74 ( .A(\data_in<9> ), .B(n1903), .Y(n14) );
  AND2X2 U75 ( .A(\data_in<10> ), .B(n1903), .Y(n15) );
  AND2X2 U76 ( .A(\data_in<11> ), .B(n1902), .Y(n16) );
  AND2X2 U77 ( .A(\data_in<12> ), .B(n1902), .Y(n17) );
  AND2X2 U78 ( .A(\data_in<13> ), .B(n1902), .Y(n18) );
  AND2X2 U79 ( .A(\data_in<14> ), .B(n1902), .Y(n19) );
  AND2X2 U80 ( .A(\data_in<15> ), .B(n1902), .Y(n20) );
  AND2X2 U81 ( .A(n1903), .B(n1245), .Y(n21) );
  AND2X2 U82 ( .A(n1903), .B(n1248), .Y(n22) );
  AND2X2 U83 ( .A(n1903), .B(n1252), .Y(n23) );
  AND2X2 U84 ( .A(n1903), .B(n1256), .Y(n24) );
  AND2X2 U85 ( .A(n1903), .B(n1260), .Y(n25) );
  AND2X2 U86 ( .A(n1903), .B(n1264), .Y(n26) );
  AND2X2 U87 ( .A(n1903), .B(n1238), .Y(n27) );
  AND2X2 U88 ( .A(n1903), .B(n1270), .Y(n28) );
  AND2X2 U89 ( .A(n1903), .B(n1274), .Y(n29) );
  AND2X2 U90 ( .A(n1903), .B(n1278), .Y(n30) );
  AND2X2 U91 ( .A(n1903), .B(n1282), .Y(n31) );
  AND2X2 U92 ( .A(n1901), .B(n1286), .Y(n32) );
  INVX1 U93 ( .A(n32), .Y(n33) );
  AND2X2 U94 ( .A(n1901), .B(n1288), .Y(n34) );
  INVX1 U95 ( .A(n34), .Y(n35) );
  AND2X2 U96 ( .A(n1901), .B(n1290), .Y(n36) );
  INVX1 U97 ( .A(n36), .Y(n37) );
  AND2X2 U98 ( .A(n1901), .B(n1239), .Y(n38) );
  INVX1 U99 ( .A(n38), .Y(n39) );
  AND2X2 U100 ( .A(n1901), .B(n1292), .Y(n40) );
  INVX1 U101 ( .A(n40), .Y(n41) );
  AND2X2 U102 ( .A(n1901), .B(n1294), .Y(n42) );
  INVX1 U103 ( .A(n42), .Y(n43) );
  AND2X2 U104 ( .A(n1901), .B(n1296), .Y(n44) );
  INVX1 U105 ( .A(n44), .Y(n45) );
  AND2X2 U106 ( .A(n1901), .B(n1298), .Y(n46) );
  INVX1 U107 ( .A(n46), .Y(n47) );
  AND2X2 U108 ( .A(n1901), .B(n1300), .Y(n48) );
  INVX1 U109 ( .A(n48), .Y(n49) );
  AND2X2 U110 ( .A(n1901), .B(n1302), .Y(n50) );
  INVX1 U111 ( .A(n50), .Y(n51) );
  AND2X2 U112 ( .A(n1901), .B(n1304), .Y(n52) );
  INVX1 U113 ( .A(n52), .Y(n53) );
  AND2X2 U114 ( .A(n1902), .B(n1240), .Y(n54) );
  INVX1 U115 ( .A(n54), .Y(n55) );
  AND2X2 U116 ( .A(n1902), .B(n1306), .Y(n56) );
  INVX1 U117 ( .A(n56), .Y(n57) );
  AND2X2 U118 ( .A(n1902), .B(n1308), .Y(n58) );
  INVX1 U119 ( .A(n58), .Y(n59) );
  AND2X2 U120 ( .A(n1902), .B(n1310), .Y(n60) );
  INVX1 U121 ( .A(n60), .Y(n61) );
  AND2X2 U122 ( .A(n1902), .B(n1312), .Y(n62) );
  INVX1 U123 ( .A(n62), .Y(n63) );
  AND2X2 U124 ( .A(n1902), .B(n1314), .Y(n64) );
  INVX1 U125 ( .A(n64), .Y(n65) );
  AND2X2 U126 ( .A(n1902), .B(n1316), .Y(n66) );
  INVX1 U127 ( .A(n66), .Y(n67) );
  AND2X2 U128 ( .A(n1902), .B(n1318), .Y(n68) );
  INVX1 U129 ( .A(n68), .Y(n69) );
  AND2X2 U130 ( .A(n1901), .B(n1241), .Y(n70) );
  INVX1 U131 ( .A(n70), .Y(n71) );
  AND2X2 U132 ( .A(\mem<19><0> ), .B(n1858), .Y(n72) );
  INVX1 U133 ( .A(n72), .Y(n73) );
  AND2X2 U134 ( .A(\mem<19><1> ), .B(n1858), .Y(n74) );
  INVX1 U135 ( .A(n74), .Y(n75) );
  AND2X2 U136 ( .A(\mem<19><2> ), .B(n1858), .Y(n76) );
  INVX1 U137 ( .A(n76), .Y(n77) );
  AND2X2 U138 ( .A(\mem<19><3> ), .B(n1858), .Y(n78) );
  INVX1 U139 ( .A(n78), .Y(n79) );
  AND2X2 U140 ( .A(\mem<19><4> ), .B(n1858), .Y(n80) );
  INVX1 U141 ( .A(n80), .Y(n81) );
  AND2X2 U142 ( .A(\mem<19><5> ), .B(n1858), .Y(n82) );
  INVX1 U143 ( .A(n82), .Y(n83) );
  AND2X2 U144 ( .A(\mem<19><6> ), .B(n1858), .Y(n84) );
  INVX1 U145 ( .A(n84), .Y(n85) );
  AND2X2 U146 ( .A(\mem<19><7> ), .B(n1858), .Y(n86) );
  INVX1 U147 ( .A(n86), .Y(n87) );
  AND2X2 U148 ( .A(\mem<19><8> ), .B(n1859), .Y(n88) );
  INVX1 U149 ( .A(n88), .Y(n89) );
  AND2X2 U150 ( .A(\mem<19><9> ), .B(n1859), .Y(n90) );
  INVX1 U151 ( .A(n90), .Y(n91) );
  AND2X2 U152 ( .A(\mem<19><10> ), .B(n1859), .Y(n92) );
  INVX1 U153 ( .A(n92), .Y(n93) );
  AND2X2 U154 ( .A(\mem<19><11> ), .B(n1859), .Y(n94) );
  INVX1 U155 ( .A(n94), .Y(n95) );
  AND2X2 U156 ( .A(\mem<19><12> ), .B(n1859), .Y(n96) );
  INVX1 U157 ( .A(n96), .Y(n97) );
  AND2X2 U158 ( .A(\mem<19><13> ), .B(n1859), .Y(n98) );
  INVX1 U159 ( .A(n98), .Y(n99) );
  AND2X2 U160 ( .A(\mem<19><14> ), .B(n1859), .Y(n100) );
  INVX1 U161 ( .A(n100), .Y(n101) );
  AND2X2 U162 ( .A(\mem<19><15> ), .B(n1859), .Y(n102) );
  INVX1 U163 ( .A(n102), .Y(n103) );
  AND2X2 U164 ( .A(\mem<18><0> ), .B(n1860), .Y(n104) );
  INVX1 U165 ( .A(n104), .Y(n105) );
  AND2X2 U166 ( .A(\mem<18><1> ), .B(n1860), .Y(n106) );
  INVX1 U167 ( .A(n106), .Y(n107) );
  AND2X2 U168 ( .A(\mem<18><2> ), .B(n1860), .Y(n108) );
  INVX1 U169 ( .A(n108), .Y(n109) );
  AND2X2 U170 ( .A(\mem<18><3> ), .B(n1860), .Y(n110) );
  INVX1 U171 ( .A(n110), .Y(n111) );
  AND2X2 U172 ( .A(\mem<18><4> ), .B(n1860), .Y(n112) );
  INVX1 U173 ( .A(n112), .Y(n113) );
  AND2X2 U174 ( .A(\mem<18><5> ), .B(n1860), .Y(n114) );
  INVX1 U175 ( .A(n114), .Y(n115) );
  AND2X2 U176 ( .A(\mem<18><6> ), .B(n1860), .Y(n116) );
  INVX1 U177 ( .A(n116), .Y(n117) );
  AND2X2 U178 ( .A(\mem<18><7> ), .B(n1860), .Y(n118) );
  INVX1 U179 ( .A(n118), .Y(n119) );
  AND2X2 U180 ( .A(\mem<18><8> ), .B(n1861), .Y(n120) );
  INVX1 U181 ( .A(n120), .Y(n121) );
  AND2X2 U182 ( .A(\mem<18><9> ), .B(n1861), .Y(n122) );
  INVX1 U183 ( .A(n122), .Y(n123) );
  AND2X2 U184 ( .A(\mem<18><10> ), .B(n1861), .Y(n124) );
  INVX1 U185 ( .A(n124), .Y(n125) );
  AND2X2 U186 ( .A(\mem<18><11> ), .B(n1861), .Y(n126) );
  INVX1 U187 ( .A(n126), .Y(n127) );
  AND2X2 U188 ( .A(\mem<18><12> ), .B(n1861), .Y(n128) );
  INVX1 U189 ( .A(n128), .Y(n129) );
  AND2X2 U190 ( .A(\mem<18><13> ), .B(n1861), .Y(n130) );
  INVX1 U191 ( .A(n130), .Y(n131) );
  AND2X2 U192 ( .A(\mem<18><14> ), .B(n1861), .Y(n132) );
  INVX1 U193 ( .A(n132), .Y(n133) );
  AND2X2 U194 ( .A(\mem<18><15> ), .B(n1861), .Y(n134) );
  INVX1 U195 ( .A(n134), .Y(n135) );
  AND2X2 U196 ( .A(\mem<17><0> ), .B(n1862), .Y(n136) );
  INVX1 U197 ( .A(n136), .Y(n137) );
  AND2X2 U198 ( .A(\mem<17><1> ), .B(n1862), .Y(n138) );
  INVX1 U199 ( .A(n138), .Y(n139) );
  AND2X2 U200 ( .A(\mem<17><2> ), .B(n1862), .Y(n140) );
  INVX1 U201 ( .A(n140), .Y(n141) );
  AND2X2 U202 ( .A(\mem<17><3> ), .B(n1862), .Y(n142) );
  INVX1 U203 ( .A(n142), .Y(n143) );
  AND2X2 U204 ( .A(\mem<17><4> ), .B(n1862), .Y(n144) );
  INVX1 U205 ( .A(n144), .Y(n145) );
  AND2X2 U206 ( .A(\mem<17><5> ), .B(n1862), .Y(n146) );
  INVX1 U207 ( .A(n146), .Y(n147) );
  AND2X2 U208 ( .A(\mem<17><6> ), .B(n1862), .Y(n148) );
  INVX1 U209 ( .A(n148), .Y(n149) );
  AND2X2 U210 ( .A(\mem<17><7> ), .B(n1862), .Y(n150) );
  INVX1 U211 ( .A(n150), .Y(n151) );
  AND2X2 U212 ( .A(\mem<17><8> ), .B(n1863), .Y(n152) );
  INVX1 U213 ( .A(n152), .Y(n153) );
  AND2X2 U214 ( .A(\mem<17><9> ), .B(n1863), .Y(n154) );
  INVX1 U215 ( .A(n154), .Y(n155) );
  AND2X2 U216 ( .A(\mem<17><10> ), .B(n1863), .Y(n156) );
  INVX1 U217 ( .A(n156), .Y(n157) );
  AND2X2 U218 ( .A(\mem<17><11> ), .B(n1863), .Y(n158) );
  INVX1 U219 ( .A(n158), .Y(n159) );
  AND2X2 U220 ( .A(\mem<17><12> ), .B(n1863), .Y(n160) );
  INVX1 U221 ( .A(n160), .Y(n161) );
  AND2X2 U222 ( .A(\mem<17><13> ), .B(n1863), .Y(n162) );
  INVX1 U223 ( .A(n162), .Y(n163) );
  AND2X2 U224 ( .A(\mem<17><14> ), .B(n1863), .Y(n164) );
  INVX1 U225 ( .A(n164), .Y(n165) );
  AND2X2 U226 ( .A(\mem<17><15> ), .B(n1863), .Y(n166) );
  INVX1 U227 ( .A(n166), .Y(n167) );
  AND2X2 U228 ( .A(\mem<16><0> ), .B(n1865), .Y(n168) );
  INVX1 U229 ( .A(n168), .Y(n169) );
  AND2X2 U230 ( .A(\mem<16><1> ), .B(n1865), .Y(n170) );
  INVX1 U231 ( .A(n170), .Y(n171) );
  AND2X2 U232 ( .A(\mem<16><2> ), .B(n1865), .Y(n172) );
  INVX1 U233 ( .A(n172), .Y(n173) );
  AND2X2 U234 ( .A(\mem<16><3> ), .B(n1865), .Y(n174) );
  INVX1 U235 ( .A(n174), .Y(n175) );
  AND2X2 U236 ( .A(\mem<16><4> ), .B(n1865), .Y(n176) );
  INVX1 U237 ( .A(n176), .Y(n177) );
  AND2X2 U238 ( .A(\mem<16><5> ), .B(n1865), .Y(n178) );
  INVX1 U239 ( .A(n178), .Y(n179) );
  AND2X2 U240 ( .A(\mem<16><6> ), .B(n1865), .Y(n180) );
  INVX1 U241 ( .A(n180), .Y(n181) );
  AND2X2 U242 ( .A(\mem<16><7> ), .B(n1865), .Y(n182) );
  INVX1 U243 ( .A(n182), .Y(n183) );
  AND2X2 U244 ( .A(\mem<16><8> ), .B(n1866), .Y(n184) );
  INVX1 U245 ( .A(n184), .Y(n185) );
  AND2X2 U246 ( .A(\mem<16><9> ), .B(n1866), .Y(n186) );
  INVX1 U247 ( .A(n186), .Y(n187) );
  AND2X2 U248 ( .A(\mem<16><10> ), .B(n1866), .Y(n188) );
  INVX1 U249 ( .A(n188), .Y(n189) );
  AND2X2 U250 ( .A(\mem<16><11> ), .B(n1866), .Y(n190) );
  INVX1 U251 ( .A(n190), .Y(n191) );
  AND2X2 U252 ( .A(\mem<16><12> ), .B(n1866), .Y(n192) );
  INVX1 U253 ( .A(n192), .Y(n193) );
  AND2X2 U254 ( .A(\mem<16><13> ), .B(n1866), .Y(n194) );
  INVX1 U255 ( .A(n194), .Y(n195) );
  AND2X2 U256 ( .A(\mem<16><14> ), .B(n1866), .Y(n196) );
  INVX1 U257 ( .A(n196), .Y(n197) );
  AND2X2 U258 ( .A(\mem<16><15> ), .B(n1866), .Y(n198) );
  INVX1 U259 ( .A(n198), .Y(n199) );
  AND2X2 U260 ( .A(\mem<15><0> ), .B(n1867), .Y(n200) );
  INVX1 U261 ( .A(n200), .Y(n201) );
  AND2X2 U262 ( .A(\mem<15><1> ), .B(n1867), .Y(n202) );
  INVX1 U263 ( .A(n202), .Y(n203) );
  AND2X2 U264 ( .A(\mem<15><2> ), .B(n1867), .Y(n204) );
  INVX1 U265 ( .A(n204), .Y(n205) );
  AND2X2 U266 ( .A(\mem<15><3> ), .B(n1867), .Y(n206) );
  INVX1 U267 ( .A(n206), .Y(n207) );
  AND2X2 U268 ( .A(\mem<15><4> ), .B(n1867), .Y(n208) );
  INVX1 U269 ( .A(n208), .Y(n209) );
  AND2X2 U270 ( .A(\mem<15><5> ), .B(n1867), .Y(n210) );
  INVX1 U271 ( .A(n210), .Y(n211) );
  AND2X2 U272 ( .A(\mem<15><6> ), .B(n1867), .Y(n212) );
  INVX1 U273 ( .A(n212), .Y(n213) );
  AND2X2 U274 ( .A(\mem<15><7> ), .B(n1867), .Y(n215) );
  INVX1 U275 ( .A(n215), .Y(n216) );
  AND2X2 U276 ( .A(\mem<15><8> ), .B(n1868), .Y(n217) );
  INVX1 U277 ( .A(n217), .Y(n218) );
  AND2X2 U278 ( .A(\mem<15><9> ), .B(n1868), .Y(n219) );
  INVX1 U279 ( .A(n219), .Y(n220) );
  AND2X2 U280 ( .A(\mem<15><10> ), .B(n1868), .Y(n221) );
  INVX1 U281 ( .A(n221), .Y(n222) );
  AND2X2 U282 ( .A(\mem<15><11> ), .B(n1868), .Y(n223) );
  INVX1 U283 ( .A(n223), .Y(n224) );
  AND2X2 U284 ( .A(\mem<15><12> ), .B(n1868), .Y(n225) );
  INVX1 U285 ( .A(n225), .Y(n226) );
  AND2X2 U286 ( .A(\mem<15><13> ), .B(n1868), .Y(n227) );
  INVX1 U287 ( .A(n227), .Y(n228) );
  AND2X2 U288 ( .A(\mem<15><14> ), .B(n1868), .Y(n229) );
  INVX1 U289 ( .A(n229), .Y(n230) );
  AND2X2 U290 ( .A(\mem<15><15> ), .B(n1868), .Y(n231) );
  INVX1 U291 ( .A(n231), .Y(n232) );
  AND2X2 U292 ( .A(\mem<14><0> ), .B(n1869), .Y(n233) );
  INVX1 U293 ( .A(n233), .Y(n234) );
  AND2X2 U294 ( .A(\mem<14><1> ), .B(n1869), .Y(n235) );
  INVX1 U295 ( .A(n235), .Y(n236) );
  AND2X2 U296 ( .A(\mem<14><2> ), .B(n1869), .Y(n237) );
  INVX1 U297 ( .A(n237), .Y(n238) );
  AND2X2 U298 ( .A(\mem<14><3> ), .B(n1869), .Y(n239) );
  INVX1 U299 ( .A(n239), .Y(n240) );
  AND2X2 U300 ( .A(\mem<14><4> ), .B(n1869), .Y(n241) );
  INVX1 U301 ( .A(n241), .Y(n242) );
  AND2X2 U302 ( .A(\mem<14><5> ), .B(n1869), .Y(n243) );
  INVX1 U303 ( .A(n243), .Y(n244) );
  AND2X2 U304 ( .A(\mem<14><6> ), .B(n1869), .Y(n245) );
  INVX1 U305 ( .A(n245), .Y(n246) );
  AND2X2 U306 ( .A(\mem<14><7> ), .B(n1869), .Y(n247) );
  INVX1 U307 ( .A(n247), .Y(n248) );
  AND2X2 U308 ( .A(\mem<14><8> ), .B(n1870), .Y(n249) );
  INVX1 U309 ( .A(n249), .Y(n250) );
  AND2X2 U310 ( .A(\mem<14><9> ), .B(n1870), .Y(n251) );
  INVX1 U311 ( .A(n251), .Y(n252) );
  AND2X2 U312 ( .A(\mem<14><10> ), .B(n1870), .Y(n253) );
  INVX1 U313 ( .A(n253), .Y(n254) );
  AND2X2 U314 ( .A(\mem<14><11> ), .B(n1870), .Y(n255) );
  INVX1 U315 ( .A(n255), .Y(n256) );
  AND2X2 U316 ( .A(\mem<14><12> ), .B(n1870), .Y(n257) );
  INVX1 U317 ( .A(n257), .Y(n258) );
  AND2X2 U318 ( .A(\mem<14><13> ), .B(n1870), .Y(n259) );
  INVX1 U319 ( .A(n259), .Y(n260) );
  AND2X2 U320 ( .A(\mem<14><14> ), .B(n1870), .Y(n261) );
  INVX1 U321 ( .A(n261), .Y(n262) );
  AND2X2 U322 ( .A(\mem<14><15> ), .B(n1870), .Y(n263) );
  INVX1 U323 ( .A(n263), .Y(n264) );
  AND2X2 U324 ( .A(\mem<13><0> ), .B(n1871), .Y(n265) );
  INVX1 U325 ( .A(n265), .Y(n266) );
  AND2X2 U326 ( .A(\mem<13><1> ), .B(n1871), .Y(n267) );
  INVX1 U327 ( .A(n267), .Y(n268) );
  AND2X2 U328 ( .A(\mem<13><2> ), .B(n1871), .Y(n269) );
  INVX1 U329 ( .A(n269), .Y(n270) );
  AND2X2 U330 ( .A(\mem<13><3> ), .B(n1871), .Y(n271) );
  INVX1 U331 ( .A(n271), .Y(n272) );
  AND2X2 U332 ( .A(\mem<13><4> ), .B(n1871), .Y(n273) );
  INVX1 U333 ( .A(n273), .Y(n274) );
  AND2X2 U334 ( .A(\mem<13><5> ), .B(n1871), .Y(n275) );
  INVX1 U335 ( .A(n275), .Y(n276) );
  AND2X2 U336 ( .A(\mem<13><6> ), .B(n1871), .Y(n277) );
  INVX1 U337 ( .A(n277), .Y(n278) );
  AND2X2 U338 ( .A(\mem<13><7> ), .B(n1871), .Y(n279) );
  INVX1 U339 ( .A(n279), .Y(n280) );
  AND2X2 U340 ( .A(\mem<13><8> ), .B(n1872), .Y(n281) );
  INVX1 U341 ( .A(n281), .Y(n282) );
  AND2X2 U342 ( .A(\mem<13><9> ), .B(n1872), .Y(n283) );
  INVX1 U343 ( .A(n283), .Y(n284) );
  AND2X2 U344 ( .A(\mem<13><10> ), .B(n1872), .Y(n285) );
  INVX1 U345 ( .A(n285), .Y(n286) );
  AND2X2 U346 ( .A(\mem<13><11> ), .B(n1872), .Y(n287) );
  INVX1 U347 ( .A(n287), .Y(n288) );
  AND2X2 U348 ( .A(\mem<13><12> ), .B(n1872), .Y(n289) );
  INVX1 U349 ( .A(n289), .Y(n290) );
  AND2X2 U350 ( .A(\mem<13><13> ), .B(n1872), .Y(n291) );
  INVX1 U351 ( .A(n291), .Y(n292) );
  AND2X2 U352 ( .A(\mem<13><14> ), .B(n1872), .Y(n293) );
  INVX1 U353 ( .A(n293), .Y(n294) );
  AND2X2 U354 ( .A(\mem<13><15> ), .B(n1872), .Y(n295) );
  INVX1 U355 ( .A(n295), .Y(n296) );
  AND2X2 U356 ( .A(\mem<12><0> ), .B(n1873), .Y(n297) );
  INVX1 U357 ( .A(n297), .Y(n298) );
  AND2X2 U358 ( .A(\mem<12><1> ), .B(n1873), .Y(n299) );
  INVX1 U359 ( .A(n299), .Y(n300) );
  AND2X2 U360 ( .A(\mem<12><2> ), .B(n1873), .Y(n301) );
  INVX1 U361 ( .A(n301), .Y(n302) );
  AND2X2 U362 ( .A(\mem<12><3> ), .B(n1873), .Y(n303) );
  INVX1 U363 ( .A(n303), .Y(n304) );
  AND2X2 U364 ( .A(\mem<12><4> ), .B(n1873), .Y(n305) );
  INVX1 U365 ( .A(n305), .Y(n306) );
  AND2X2 U366 ( .A(\mem<12><5> ), .B(n1873), .Y(n307) );
  INVX1 U367 ( .A(n307), .Y(n308) );
  AND2X2 U368 ( .A(\mem<12><6> ), .B(n1873), .Y(n309) );
  INVX1 U369 ( .A(n309), .Y(n310) );
  AND2X2 U370 ( .A(\mem<12><7> ), .B(n1873), .Y(n311) );
  INVX1 U371 ( .A(n311), .Y(n312) );
  AND2X2 U372 ( .A(\mem<12><8> ), .B(n1874), .Y(n313) );
  INVX1 U373 ( .A(n313), .Y(n314) );
  AND2X2 U374 ( .A(\mem<12><9> ), .B(n1874), .Y(n315) );
  INVX1 U375 ( .A(n315), .Y(n316) );
  AND2X2 U376 ( .A(\mem<12><10> ), .B(n1874), .Y(n317) );
  INVX1 U377 ( .A(n317), .Y(n318) );
  AND2X2 U378 ( .A(\mem<12><11> ), .B(n1874), .Y(n319) );
  INVX1 U379 ( .A(n319), .Y(n320) );
  AND2X2 U380 ( .A(\mem<12><12> ), .B(n1874), .Y(n321) );
  INVX1 U381 ( .A(n321), .Y(n322) );
  AND2X2 U382 ( .A(\mem<12><13> ), .B(n1874), .Y(n323) );
  INVX1 U383 ( .A(n323), .Y(n324) );
  AND2X2 U384 ( .A(\mem<12><14> ), .B(n1874), .Y(n325) );
  INVX1 U385 ( .A(n325), .Y(n326) );
  AND2X2 U386 ( .A(\mem<12><15> ), .B(n1874), .Y(n327) );
  INVX1 U387 ( .A(n327), .Y(n328) );
  AND2X2 U388 ( .A(\mem<11><0> ), .B(n1875), .Y(n329) );
  INVX1 U389 ( .A(n329), .Y(n330) );
  AND2X2 U390 ( .A(\mem<11><1> ), .B(n1875), .Y(n331) );
  INVX1 U391 ( .A(n331), .Y(n332) );
  AND2X2 U392 ( .A(\mem<11><2> ), .B(n1875), .Y(n333) );
  INVX1 U393 ( .A(n333), .Y(n334) );
  AND2X2 U394 ( .A(\mem<11><3> ), .B(n1875), .Y(n335) );
  INVX1 U395 ( .A(n335), .Y(n336) );
  AND2X2 U396 ( .A(\mem<11><4> ), .B(n1875), .Y(n337) );
  INVX1 U397 ( .A(n337), .Y(n338) );
  AND2X2 U398 ( .A(\mem<11><5> ), .B(n1875), .Y(n339) );
  INVX1 U399 ( .A(n339), .Y(n340) );
  AND2X2 U400 ( .A(\mem<11><6> ), .B(n1875), .Y(n341) );
  INVX1 U401 ( .A(n341), .Y(n342) );
  AND2X2 U402 ( .A(\mem<11><7> ), .B(n1875), .Y(n343) );
  INVX1 U403 ( .A(n343), .Y(n344) );
  AND2X2 U404 ( .A(\mem<11><8> ), .B(n1876), .Y(n345) );
  INVX1 U405 ( .A(n345), .Y(n346) );
  AND2X2 U406 ( .A(\mem<11><9> ), .B(n1876), .Y(n347) );
  INVX1 U407 ( .A(n347), .Y(n348) );
  AND2X2 U408 ( .A(\mem<11><10> ), .B(n1876), .Y(n349) );
  INVX1 U409 ( .A(n349), .Y(n350) );
  AND2X2 U410 ( .A(\mem<11><11> ), .B(n1876), .Y(n351) );
  INVX1 U411 ( .A(n351), .Y(n352) );
  AND2X2 U412 ( .A(\mem<11><12> ), .B(n1876), .Y(n353) );
  INVX1 U413 ( .A(n353), .Y(n354) );
  AND2X2 U414 ( .A(\mem<11><13> ), .B(n1876), .Y(n355) );
  INVX1 U415 ( .A(n355), .Y(n356) );
  AND2X2 U416 ( .A(\mem<11><14> ), .B(n1876), .Y(n357) );
  INVX1 U417 ( .A(n357), .Y(n358) );
  AND2X2 U418 ( .A(\mem<11><15> ), .B(n1876), .Y(n359) );
  INVX1 U419 ( .A(n359), .Y(n360) );
  AND2X2 U420 ( .A(\mem<10><0> ), .B(n1877), .Y(n361) );
  INVX1 U421 ( .A(n361), .Y(n362) );
  AND2X2 U422 ( .A(\mem<10><1> ), .B(n1877), .Y(n363) );
  INVX1 U423 ( .A(n363), .Y(n364) );
  AND2X2 U424 ( .A(\mem<10><2> ), .B(n1877), .Y(n365) );
  INVX1 U425 ( .A(n365), .Y(n366) );
  AND2X2 U426 ( .A(\mem<10><3> ), .B(n1877), .Y(n367) );
  INVX1 U427 ( .A(n367), .Y(n368) );
  AND2X2 U428 ( .A(\mem<10><4> ), .B(n1877), .Y(n369) );
  INVX1 U429 ( .A(n369), .Y(n370) );
  AND2X2 U430 ( .A(\mem<10><5> ), .B(n1877), .Y(n371) );
  INVX1 U431 ( .A(n371), .Y(n372) );
  AND2X2 U432 ( .A(\mem<10><6> ), .B(n1877), .Y(n373) );
  INVX1 U433 ( .A(n373), .Y(n374) );
  AND2X2 U434 ( .A(\mem<10><7> ), .B(n1877), .Y(n375) );
  INVX1 U435 ( .A(n375), .Y(n376) );
  AND2X2 U436 ( .A(\mem<10><8> ), .B(n1878), .Y(n377) );
  INVX1 U437 ( .A(n377), .Y(n378) );
  AND2X2 U438 ( .A(\mem<10><9> ), .B(n1878), .Y(n379) );
  INVX1 U439 ( .A(n379), .Y(n380) );
  AND2X2 U440 ( .A(\mem<10><10> ), .B(n1878), .Y(n381) );
  INVX1 U441 ( .A(n381), .Y(n382) );
  AND2X2 U442 ( .A(\mem<10><11> ), .B(n1878), .Y(n383) );
  INVX1 U443 ( .A(n383), .Y(n384) );
  AND2X2 U444 ( .A(\mem<10><12> ), .B(n1878), .Y(n385) );
  INVX1 U445 ( .A(n385), .Y(n386) );
  AND2X2 U446 ( .A(\mem<10><13> ), .B(n1878), .Y(n387) );
  INVX1 U447 ( .A(n387), .Y(n388) );
  AND2X2 U448 ( .A(\mem<10><14> ), .B(n1878), .Y(n389) );
  INVX1 U449 ( .A(n389), .Y(n390) );
  AND2X2 U450 ( .A(\mem<10><15> ), .B(n1878), .Y(n391) );
  INVX1 U451 ( .A(n391), .Y(n392) );
  AND2X2 U452 ( .A(\mem<9><0> ), .B(n1879), .Y(n393) );
  INVX1 U453 ( .A(n393), .Y(n394) );
  AND2X2 U454 ( .A(\mem<9><1> ), .B(n1879), .Y(n395) );
  INVX1 U455 ( .A(n395), .Y(n396) );
  AND2X2 U456 ( .A(\mem<9><2> ), .B(n1879), .Y(n397) );
  INVX1 U457 ( .A(n397), .Y(n398) );
  AND2X2 U458 ( .A(\mem<9><3> ), .B(n1879), .Y(n399) );
  INVX1 U459 ( .A(n399), .Y(n400) );
  AND2X2 U460 ( .A(\mem<9><4> ), .B(n1879), .Y(n401) );
  INVX1 U461 ( .A(n401), .Y(n402) );
  AND2X2 U462 ( .A(\mem<9><5> ), .B(n1879), .Y(n403) );
  INVX1 U463 ( .A(n403), .Y(n404) );
  AND2X2 U464 ( .A(\mem<9><6> ), .B(n1879), .Y(n405) );
  INVX1 U465 ( .A(n405), .Y(n406) );
  AND2X2 U466 ( .A(\mem<9><7> ), .B(n1879), .Y(n407) );
  INVX1 U467 ( .A(n407), .Y(n408) );
  AND2X2 U468 ( .A(\mem<9><8> ), .B(n1880), .Y(n409) );
  INVX1 U469 ( .A(n409), .Y(n410) );
  AND2X2 U470 ( .A(\mem<9><9> ), .B(n1880), .Y(n411) );
  INVX1 U471 ( .A(n411), .Y(n412) );
  AND2X2 U472 ( .A(\mem<9><10> ), .B(n1880), .Y(n413) );
  INVX1 U473 ( .A(n413), .Y(n414) );
  AND2X2 U474 ( .A(\mem<9><11> ), .B(n1880), .Y(n415) );
  INVX1 U475 ( .A(n415), .Y(n416) );
  AND2X2 U476 ( .A(\mem<9><12> ), .B(n1880), .Y(n417) );
  INVX1 U477 ( .A(n417), .Y(n418) );
  AND2X2 U478 ( .A(\mem<9><13> ), .B(n1880), .Y(n419) );
  INVX1 U479 ( .A(n419), .Y(n420) );
  AND2X2 U480 ( .A(\mem<9><14> ), .B(n1880), .Y(n421) );
  INVX1 U481 ( .A(n421), .Y(n422) );
  AND2X2 U482 ( .A(\mem<9><15> ), .B(n1880), .Y(n423) );
  INVX1 U483 ( .A(n423), .Y(n424) );
  AND2X2 U484 ( .A(\mem<8><0> ), .B(n1882), .Y(n425) );
  INVX1 U485 ( .A(n425), .Y(n426) );
  AND2X2 U486 ( .A(\mem<8><1> ), .B(n1882), .Y(n427) );
  INVX1 U487 ( .A(n427), .Y(n428) );
  AND2X2 U488 ( .A(\mem<8><2> ), .B(n1882), .Y(n429) );
  INVX1 U489 ( .A(n429), .Y(n430) );
  AND2X2 U490 ( .A(\mem<8><3> ), .B(n1882), .Y(n431) );
  INVX1 U491 ( .A(n431), .Y(n432) );
  AND2X2 U492 ( .A(\mem<8><4> ), .B(n1882), .Y(n433) );
  INVX1 U493 ( .A(n433), .Y(n434) );
  AND2X2 U494 ( .A(\mem<8><5> ), .B(n1882), .Y(n435) );
  INVX1 U495 ( .A(n435), .Y(n436) );
  AND2X2 U496 ( .A(\mem<8><6> ), .B(n1882), .Y(n437) );
  INVX1 U497 ( .A(n437), .Y(n438) );
  AND2X2 U498 ( .A(\mem<8><7> ), .B(n1882), .Y(n439) );
  INVX1 U499 ( .A(n439), .Y(n440) );
  AND2X2 U500 ( .A(\mem<8><8> ), .B(n1883), .Y(n441) );
  INVX1 U501 ( .A(n441), .Y(n442) );
  AND2X2 U502 ( .A(\mem<8><9> ), .B(n1883), .Y(n443) );
  INVX1 U503 ( .A(n443), .Y(n444) );
  AND2X2 U504 ( .A(\mem<8><10> ), .B(n1883), .Y(n445) );
  INVX1 U505 ( .A(n445), .Y(n446) );
  AND2X2 U506 ( .A(\mem<8><11> ), .B(n1883), .Y(n447) );
  INVX1 U507 ( .A(n447), .Y(n448) );
  AND2X2 U508 ( .A(\mem<8><12> ), .B(n1883), .Y(n449) );
  INVX1 U509 ( .A(n449), .Y(n450) );
  AND2X2 U510 ( .A(\mem<8><13> ), .B(n1883), .Y(n451) );
  INVX1 U511 ( .A(n451), .Y(n452) );
  AND2X2 U512 ( .A(\mem<8><14> ), .B(n1883), .Y(n453) );
  INVX1 U513 ( .A(n453), .Y(n454) );
  AND2X2 U514 ( .A(\mem<8><15> ), .B(n1883), .Y(n455) );
  INVX1 U515 ( .A(n455), .Y(n456) );
  AND2X2 U516 ( .A(\mem<7><0> ), .B(n1884), .Y(n457) );
  INVX1 U517 ( .A(n457), .Y(n458) );
  AND2X2 U518 ( .A(\mem<7><1> ), .B(n1884), .Y(n459) );
  INVX1 U519 ( .A(n459), .Y(n460) );
  AND2X2 U520 ( .A(\mem<7><2> ), .B(n1884), .Y(n461) );
  INVX1 U521 ( .A(n461), .Y(n462) );
  AND2X2 U522 ( .A(\mem<7><3> ), .B(n1884), .Y(n463) );
  INVX1 U523 ( .A(n463), .Y(n464) );
  AND2X2 U524 ( .A(\mem<7><4> ), .B(n1884), .Y(n465) );
  INVX1 U525 ( .A(n465), .Y(n466) );
  AND2X2 U526 ( .A(\mem<7><5> ), .B(n1884), .Y(n467) );
  INVX1 U527 ( .A(n467), .Y(n468) );
  AND2X2 U528 ( .A(\mem<7><6> ), .B(n1884), .Y(n469) );
  INVX1 U529 ( .A(n469), .Y(n470) );
  AND2X2 U530 ( .A(\mem<7><7> ), .B(n1884), .Y(n471) );
  INVX1 U531 ( .A(n471), .Y(n472) );
  AND2X2 U532 ( .A(\mem<7><8> ), .B(n1885), .Y(n473) );
  INVX1 U533 ( .A(n473), .Y(n474) );
  AND2X2 U534 ( .A(\mem<7><9> ), .B(n1885), .Y(n475) );
  INVX1 U535 ( .A(n475), .Y(n476) );
  AND2X2 U536 ( .A(\mem<7><10> ), .B(n1885), .Y(n477) );
  INVX1 U537 ( .A(n477), .Y(n478) );
  AND2X2 U538 ( .A(\mem<7><11> ), .B(n1885), .Y(n479) );
  INVX1 U539 ( .A(n479), .Y(n480) );
  AND2X2 U540 ( .A(\mem<7><12> ), .B(n1885), .Y(n481) );
  INVX1 U541 ( .A(n481), .Y(n482) );
  AND2X2 U542 ( .A(\mem<7><13> ), .B(n1885), .Y(n483) );
  INVX1 U543 ( .A(n483), .Y(n484) );
  AND2X2 U544 ( .A(\mem<7><14> ), .B(n1885), .Y(n485) );
  INVX1 U545 ( .A(n485), .Y(n486) );
  AND2X2 U546 ( .A(\mem<7><15> ), .B(n1885), .Y(n487) );
  INVX1 U547 ( .A(n487), .Y(n488) );
  AND2X2 U548 ( .A(\mem<6><0> ), .B(n1886), .Y(n489) );
  INVX1 U549 ( .A(n489), .Y(n490) );
  AND2X2 U550 ( .A(\mem<6><1> ), .B(n1886), .Y(n491) );
  INVX1 U551 ( .A(n491), .Y(n492) );
  AND2X2 U552 ( .A(\mem<6><2> ), .B(n1886), .Y(n493) );
  INVX1 U553 ( .A(n493), .Y(n494) );
  AND2X2 U554 ( .A(\mem<6><3> ), .B(n1886), .Y(n495) );
  INVX1 U555 ( .A(n495), .Y(n496) );
  AND2X2 U556 ( .A(\mem<6><4> ), .B(n1886), .Y(n497) );
  INVX1 U557 ( .A(n497), .Y(n498) );
  AND2X2 U558 ( .A(\mem<6><5> ), .B(n1886), .Y(n499) );
  INVX1 U559 ( .A(n499), .Y(n500) );
  AND2X2 U560 ( .A(\mem<6><6> ), .B(n1886), .Y(n501) );
  INVX1 U561 ( .A(n501), .Y(n502) );
  AND2X2 U562 ( .A(\mem<6><7> ), .B(n1886), .Y(n503) );
  INVX1 U563 ( .A(n503), .Y(n504) );
  AND2X2 U564 ( .A(\mem<6><8> ), .B(n1887), .Y(n505) );
  INVX1 U565 ( .A(n505), .Y(n506) );
  AND2X2 U566 ( .A(\mem<6><9> ), .B(n1887), .Y(n507) );
  INVX1 U567 ( .A(n507), .Y(n508) );
  AND2X2 U568 ( .A(\mem<6><10> ), .B(n1887), .Y(n509) );
  INVX1 U569 ( .A(n509), .Y(n510) );
  AND2X2 U570 ( .A(\mem<6><11> ), .B(n1887), .Y(n511) );
  INVX1 U571 ( .A(n511), .Y(n512) );
  AND2X2 U572 ( .A(\mem<6><12> ), .B(n1887), .Y(n513) );
  INVX1 U573 ( .A(n513), .Y(n514) );
  AND2X2 U574 ( .A(\mem<6><13> ), .B(n1887), .Y(n515) );
  INVX1 U575 ( .A(n515), .Y(n516) );
  AND2X2 U576 ( .A(\mem<6><14> ), .B(n1887), .Y(n517) );
  INVX1 U577 ( .A(n517), .Y(n518) );
  AND2X2 U578 ( .A(\mem<6><15> ), .B(n1887), .Y(n519) );
  INVX1 U579 ( .A(n519), .Y(n520) );
  AND2X2 U580 ( .A(\mem<5><0> ), .B(n1888), .Y(n521) );
  INVX1 U581 ( .A(n521), .Y(n522) );
  AND2X2 U582 ( .A(\mem<5><1> ), .B(n1888), .Y(n523) );
  INVX1 U583 ( .A(n523), .Y(n524) );
  AND2X2 U584 ( .A(\mem<5><2> ), .B(n1888), .Y(n525) );
  INVX1 U585 ( .A(n525), .Y(n526) );
  AND2X2 U586 ( .A(\mem<5><3> ), .B(n1888), .Y(n527) );
  INVX1 U587 ( .A(n527), .Y(n528) );
  AND2X2 U588 ( .A(\mem<5><4> ), .B(n1888), .Y(n529) );
  INVX1 U589 ( .A(n529), .Y(n530) );
  AND2X2 U590 ( .A(\mem<5><5> ), .B(n1888), .Y(n531) );
  INVX1 U591 ( .A(n531), .Y(n532) );
  AND2X2 U592 ( .A(\mem<5><6> ), .B(n1888), .Y(n533) );
  INVX1 U593 ( .A(n533), .Y(n534) );
  AND2X2 U594 ( .A(\mem<5><7> ), .B(n1888), .Y(n535) );
  INVX1 U595 ( .A(n535), .Y(n536) );
  AND2X2 U596 ( .A(\mem<5><8> ), .B(n1889), .Y(n537) );
  INVX1 U597 ( .A(n537), .Y(n538) );
  AND2X2 U598 ( .A(\mem<5><9> ), .B(n1889), .Y(n539) );
  INVX1 U599 ( .A(n539), .Y(n540) );
  AND2X2 U600 ( .A(\mem<5><10> ), .B(n1889), .Y(n541) );
  INVX1 U601 ( .A(n541), .Y(n542) );
  AND2X2 U602 ( .A(\mem<5><11> ), .B(n1889), .Y(n543) );
  INVX1 U603 ( .A(n543), .Y(n544) );
  AND2X2 U604 ( .A(\mem<5><12> ), .B(n1889), .Y(n545) );
  INVX1 U605 ( .A(n545), .Y(n546) );
  AND2X2 U606 ( .A(\mem<5><13> ), .B(n1889), .Y(n547) );
  INVX1 U607 ( .A(n547), .Y(n548) );
  AND2X2 U608 ( .A(\mem<5><14> ), .B(n1889), .Y(n549) );
  INVX1 U609 ( .A(n549), .Y(n550) );
  AND2X2 U610 ( .A(\mem<5><15> ), .B(n1889), .Y(n551) );
  INVX1 U611 ( .A(n551), .Y(n552) );
  AND2X2 U612 ( .A(\mem<4><0> ), .B(n1890), .Y(n553) );
  INVX1 U613 ( .A(n553), .Y(n554) );
  AND2X2 U614 ( .A(\mem<4><1> ), .B(n1890), .Y(n555) );
  INVX1 U615 ( .A(n555), .Y(n556) );
  AND2X2 U616 ( .A(\mem<4><2> ), .B(n1890), .Y(n557) );
  INVX1 U617 ( .A(n557), .Y(n558) );
  AND2X2 U618 ( .A(\mem<4><3> ), .B(n1890), .Y(n559) );
  INVX1 U619 ( .A(n559), .Y(n560) );
  AND2X2 U620 ( .A(\mem<4><4> ), .B(n1890), .Y(n561) );
  INVX1 U621 ( .A(n561), .Y(n562) );
  AND2X2 U622 ( .A(\mem<4><5> ), .B(n1890), .Y(n563) );
  INVX1 U623 ( .A(n563), .Y(n564) );
  AND2X2 U624 ( .A(\mem<4><6> ), .B(n1890), .Y(n565) );
  INVX1 U625 ( .A(n565), .Y(n566) );
  AND2X2 U626 ( .A(\mem<4><7> ), .B(n1890), .Y(n567) );
  INVX1 U627 ( .A(n567), .Y(n568) );
  AND2X2 U628 ( .A(\mem<4><8> ), .B(n1891), .Y(n569) );
  INVX1 U629 ( .A(n569), .Y(n570) );
  AND2X2 U630 ( .A(\mem<4><9> ), .B(n1891), .Y(n571) );
  INVX1 U631 ( .A(n571), .Y(n572) );
  AND2X2 U632 ( .A(\mem<4><10> ), .B(n1891), .Y(n573) );
  INVX1 U633 ( .A(n573), .Y(n574) );
  AND2X2 U634 ( .A(\mem<4><11> ), .B(n1891), .Y(n575) );
  INVX1 U635 ( .A(n575), .Y(n576) );
  AND2X2 U636 ( .A(\mem<4><12> ), .B(n1891), .Y(n577) );
  INVX1 U637 ( .A(n577), .Y(n578) );
  AND2X2 U638 ( .A(\mem<4><13> ), .B(n1891), .Y(n579) );
  INVX1 U639 ( .A(n579), .Y(n580) );
  AND2X2 U640 ( .A(\mem<4><14> ), .B(n1891), .Y(n581) );
  INVX1 U641 ( .A(n581), .Y(n582) );
  AND2X2 U642 ( .A(\mem<4><15> ), .B(n1891), .Y(n583) );
  INVX1 U643 ( .A(n583), .Y(n584) );
  AND2X2 U644 ( .A(\mem<3><0> ), .B(n1892), .Y(n585) );
  INVX1 U645 ( .A(n585), .Y(n586) );
  AND2X2 U646 ( .A(\mem<3><1> ), .B(n1892), .Y(n587) );
  INVX1 U647 ( .A(n587), .Y(n588) );
  AND2X2 U648 ( .A(\mem<3><2> ), .B(n1892), .Y(n589) );
  INVX1 U649 ( .A(n589), .Y(n590) );
  AND2X2 U650 ( .A(\mem<3><3> ), .B(n1892), .Y(n591) );
  INVX1 U651 ( .A(n591), .Y(n592) );
  AND2X2 U652 ( .A(\mem<3><4> ), .B(n1892), .Y(n593) );
  INVX1 U653 ( .A(n593), .Y(n594) );
  AND2X2 U654 ( .A(\mem<3><5> ), .B(n1892), .Y(n595) );
  INVX1 U655 ( .A(n595), .Y(n596) );
  AND2X2 U656 ( .A(\mem<3><6> ), .B(n1892), .Y(n597) );
  INVX1 U657 ( .A(n597), .Y(n598) );
  AND2X2 U658 ( .A(\mem<3><7> ), .B(n1892), .Y(n599) );
  INVX1 U659 ( .A(n599), .Y(n600) );
  AND2X2 U660 ( .A(\mem<3><8> ), .B(n1893), .Y(n601) );
  INVX1 U661 ( .A(n601), .Y(n602) );
  AND2X2 U662 ( .A(\mem<3><9> ), .B(n1893), .Y(n603) );
  INVX1 U663 ( .A(n603), .Y(n604) );
  AND2X2 U664 ( .A(\mem<3><10> ), .B(n1893), .Y(n605) );
  INVX1 U665 ( .A(n605), .Y(n606) );
  AND2X2 U666 ( .A(\mem<3><11> ), .B(n1893), .Y(n607) );
  INVX1 U667 ( .A(n607), .Y(n608) );
  AND2X2 U668 ( .A(\mem<3><12> ), .B(n1893), .Y(n609) );
  INVX1 U669 ( .A(n609), .Y(n610) );
  AND2X2 U670 ( .A(\mem<3><13> ), .B(n1893), .Y(n611) );
  INVX1 U671 ( .A(n611), .Y(n612) );
  AND2X2 U672 ( .A(\mem<3><14> ), .B(n1893), .Y(n613) );
  INVX1 U673 ( .A(n613), .Y(n614) );
  AND2X2 U674 ( .A(\mem<3><15> ), .B(n1893), .Y(n615) );
  INVX1 U675 ( .A(n615), .Y(n616) );
  AND2X2 U676 ( .A(\mem<2><0> ), .B(n1894), .Y(n617) );
  INVX1 U677 ( .A(n617), .Y(n618) );
  AND2X2 U678 ( .A(\mem<2><1> ), .B(n1894), .Y(n619) );
  INVX1 U679 ( .A(n619), .Y(n620) );
  AND2X2 U680 ( .A(\mem<2><2> ), .B(n1894), .Y(n621) );
  INVX1 U681 ( .A(n621), .Y(n622) );
  AND2X2 U682 ( .A(\mem<2><3> ), .B(n1894), .Y(n623) );
  INVX1 U683 ( .A(n623), .Y(n624) );
  AND2X2 U684 ( .A(\mem<2><4> ), .B(n1894), .Y(n625) );
  INVX1 U685 ( .A(n625), .Y(n626) );
  AND2X2 U686 ( .A(\mem<2><5> ), .B(n1894), .Y(n627) );
  INVX1 U687 ( .A(n627), .Y(n628) );
  AND2X2 U688 ( .A(\mem<2><6> ), .B(n1894), .Y(n629) );
  INVX1 U689 ( .A(n629), .Y(n630) );
  AND2X2 U690 ( .A(\mem<2><7> ), .B(n1894), .Y(n631) );
  INVX1 U691 ( .A(n631), .Y(n632) );
  AND2X2 U692 ( .A(\mem<2><8> ), .B(n1895), .Y(n633) );
  INVX1 U693 ( .A(n633), .Y(n634) );
  AND2X2 U694 ( .A(\mem<2><9> ), .B(n1895), .Y(n635) );
  INVX1 U695 ( .A(n635), .Y(n636) );
  AND2X2 U696 ( .A(\mem<2><10> ), .B(n1895), .Y(n637) );
  INVX1 U697 ( .A(n637), .Y(n638) );
  AND2X2 U698 ( .A(\mem<2><11> ), .B(n1895), .Y(n639) );
  INVX1 U699 ( .A(n639), .Y(n640) );
  AND2X2 U700 ( .A(\mem<2><12> ), .B(n1895), .Y(n641) );
  INVX1 U701 ( .A(n641), .Y(n642) );
  AND2X2 U702 ( .A(\mem<2><13> ), .B(n1895), .Y(n643) );
  INVX1 U703 ( .A(n643), .Y(n644) );
  AND2X2 U704 ( .A(\mem<2><14> ), .B(n1895), .Y(n645) );
  INVX1 U705 ( .A(n645), .Y(n646) );
  AND2X2 U706 ( .A(\mem<2><15> ), .B(n1895), .Y(n647) );
  INVX1 U707 ( .A(n647), .Y(n648) );
  AND2X2 U708 ( .A(\mem<1><0> ), .B(n1896), .Y(n649) );
  INVX1 U709 ( .A(n649), .Y(n650) );
  AND2X2 U710 ( .A(\mem<1><1> ), .B(n1896), .Y(n1163) );
  INVX1 U711 ( .A(n1163), .Y(n1164) );
  AND2X2 U712 ( .A(\mem<1><2> ), .B(n1896), .Y(n1165) );
  INVX1 U713 ( .A(n1165), .Y(n1166) );
  AND2X2 U714 ( .A(\mem<1><3> ), .B(n1896), .Y(n1167) );
  INVX1 U715 ( .A(n1167), .Y(n1168) );
  AND2X2 U716 ( .A(\mem<1><4> ), .B(n1896), .Y(n1169) );
  INVX1 U717 ( .A(n1169), .Y(n1170) );
  AND2X2 U718 ( .A(\mem<1><5> ), .B(n1896), .Y(n1171) );
  INVX1 U719 ( .A(n1171), .Y(n1172) );
  AND2X2 U720 ( .A(\mem<1><6> ), .B(n1896), .Y(n1173) );
  INVX1 U721 ( .A(n1173), .Y(n1174) );
  AND2X2 U722 ( .A(\mem<1><7> ), .B(n1896), .Y(n1175) );
  INVX1 U723 ( .A(n1175), .Y(n1176) );
  AND2X2 U724 ( .A(\mem<1><8> ), .B(n1897), .Y(n1177) );
  INVX1 U725 ( .A(n1177), .Y(n1178) );
  AND2X2 U726 ( .A(\mem<1><9> ), .B(n1897), .Y(n1179) );
  INVX1 U727 ( .A(n1179), .Y(n1180) );
  AND2X2 U728 ( .A(\mem<1><10> ), .B(n1897), .Y(n1181) );
  INVX1 U729 ( .A(n1181), .Y(n1182) );
  AND2X2 U730 ( .A(\mem<1><11> ), .B(n1897), .Y(n1183) );
  INVX1 U731 ( .A(n1183), .Y(n1184) );
  AND2X2 U732 ( .A(\mem<1><12> ), .B(n1897), .Y(n1185) );
  INVX1 U733 ( .A(n1185), .Y(n1186) );
  AND2X2 U734 ( .A(\mem<1><13> ), .B(n1897), .Y(n1187) );
  INVX1 U735 ( .A(n1187), .Y(n1188) );
  AND2X2 U736 ( .A(\mem<1><14> ), .B(n1897), .Y(n1189) );
  INVX1 U737 ( .A(n1189), .Y(n1190) );
  AND2X2 U738 ( .A(\mem<1><15> ), .B(n1897), .Y(n1191) );
  INVX1 U739 ( .A(n1191), .Y(n1192) );
  AND2X2 U740 ( .A(\mem<0><0> ), .B(n1899), .Y(n1193) );
  INVX1 U741 ( .A(n1193), .Y(n1194) );
  AND2X2 U742 ( .A(\mem<0><1> ), .B(n1899), .Y(n1195) );
  INVX1 U743 ( .A(n1195), .Y(n1196) );
  AND2X2 U744 ( .A(\mem<0><2> ), .B(n1899), .Y(n1197) );
  INVX1 U745 ( .A(n1197), .Y(n1198) );
  AND2X2 U746 ( .A(\mem<0><3> ), .B(n1899), .Y(n1199) );
  INVX1 U747 ( .A(n1199), .Y(n1200) );
  AND2X2 U748 ( .A(\mem<0><4> ), .B(n1899), .Y(n1201) );
  INVX1 U749 ( .A(n1201), .Y(n1202) );
  AND2X2 U750 ( .A(\mem<0><5> ), .B(n1899), .Y(n1203) );
  INVX1 U751 ( .A(n1203), .Y(n1204) );
  AND2X2 U752 ( .A(\mem<0><6> ), .B(n1899), .Y(n1205) );
  INVX1 U753 ( .A(n1205), .Y(n1206) );
  AND2X2 U754 ( .A(\mem<0><7> ), .B(n1899), .Y(n1207) );
  INVX1 U755 ( .A(n1207), .Y(n1208) );
  AND2X2 U756 ( .A(\mem<0><8> ), .B(n1900), .Y(n1209) );
  INVX1 U757 ( .A(n1209), .Y(n1210) );
  AND2X2 U758 ( .A(\mem<0><9> ), .B(n1900), .Y(n1211) );
  INVX1 U759 ( .A(n1211), .Y(n1212) );
  AND2X2 U760 ( .A(\mem<0><10> ), .B(n1900), .Y(n1213) );
  INVX1 U761 ( .A(n1213), .Y(n1214) );
  AND2X2 U762 ( .A(\mem<0><11> ), .B(n1900), .Y(n1215) );
  INVX1 U763 ( .A(n1215), .Y(n1216) );
  AND2X2 U764 ( .A(\mem<0><12> ), .B(n1900), .Y(n1217) );
  INVX1 U765 ( .A(n1217), .Y(n1218) );
  AND2X2 U766 ( .A(\mem<0><13> ), .B(n1900), .Y(n1219) );
  INVX1 U767 ( .A(n1219), .Y(n1220) );
  AND2X2 U768 ( .A(\mem<0><14> ), .B(n1900), .Y(n1221) );
  INVX1 U769 ( .A(n1221), .Y(n1222) );
  AND2X2 U770 ( .A(\mem<0><15> ), .B(n1900), .Y(n1223) );
  INVX1 U771 ( .A(n1223), .Y(n1224) );
  INVX1 U772 ( .A(n1940), .Y(n1939) );
  INVX1 U773 ( .A(N14), .Y(n1944) );
  AND2X1 U774 ( .A(n1941), .B(n1939), .Y(n1225) );
  INVX1 U775 ( .A(n1942), .Y(n1941) );
  AND2X1 U776 ( .A(n2664), .B(N14), .Y(n1226) );
  BUFX2 U777 ( .A(n33), .Y(n1858) );
  BUFX2 U778 ( .A(n33), .Y(n1859) );
  BUFX2 U779 ( .A(n35), .Y(n1860) );
  BUFX2 U780 ( .A(n35), .Y(n1861) );
  BUFX2 U781 ( .A(n37), .Y(n1862) );
  BUFX2 U782 ( .A(n37), .Y(n1863) );
  BUFX2 U783 ( .A(n39), .Y(n1865) );
  BUFX2 U784 ( .A(n39), .Y(n1866) );
  BUFX2 U785 ( .A(n41), .Y(n1867) );
  BUFX2 U786 ( .A(n41), .Y(n1868) );
  BUFX2 U787 ( .A(n43), .Y(n1869) );
  BUFX2 U788 ( .A(n43), .Y(n1870) );
  BUFX2 U789 ( .A(n45), .Y(n1871) );
  BUFX2 U790 ( .A(n45), .Y(n1872) );
  BUFX2 U791 ( .A(n47), .Y(n1873) );
  BUFX2 U792 ( .A(n47), .Y(n1874) );
  BUFX2 U793 ( .A(n49), .Y(n1875) );
  BUFX2 U794 ( .A(n49), .Y(n1876) );
  BUFX2 U795 ( .A(n51), .Y(n1877) );
  BUFX2 U796 ( .A(n51), .Y(n1878) );
  BUFX2 U797 ( .A(n53), .Y(n1879) );
  BUFX2 U798 ( .A(n53), .Y(n1880) );
  BUFX2 U799 ( .A(n55), .Y(n1882) );
  BUFX2 U800 ( .A(n55), .Y(n1883) );
  BUFX2 U801 ( .A(n57), .Y(n1884) );
  BUFX2 U802 ( .A(n57), .Y(n1885) );
  BUFX2 U803 ( .A(n59), .Y(n1886) );
  BUFX2 U804 ( .A(n59), .Y(n1887) );
  BUFX2 U805 ( .A(n61), .Y(n1888) );
  BUFX2 U806 ( .A(n61), .Y(n1889) );
  BUFX2 U807 ( .A(n63), .Y(n1890) );
  BUFX2 U808 ( .A(n63), .Y(n1891) );
  BUFX2 U809 ( .A(n65), .Y(n1892) );
  BUFX2 U810 ( .A(n65), .Y(n1893) );
  BUFX2 U811 ( .A(n67), .Y(n1894) );
  BUFX2 U812 ( .A(n67), .Y(n1895) );
  BUFX2 U813 ( .A(n69), .Y(n1896) );
  BUFX2 U814 ( .A(n69), .Y(n1897) );
  BUFX2 U815 ( .A(n71), .Y(n1899) );
  BUFX2 U816 ( .A(n71), .Y(n1900) );
  BUFX2 U817 ( .A(n1977), .Y(n1227) );
  INVX1 U818 ( .A(n1227), .Y(n2145) );
  BUFX2 U819 ( .A(n1994), .Y(n1228) );
  INVX1 U820 ( .A(n1228), .Y(n2146) );
  BUFX2 U821 ( .A(n2011), .Y(n1229) );
  INVX1 U822 ( .A(n1229), .Y(n2147) );
  BUFX2 U823 ( .A(n2028), .Y(n1230) );
  INVX1 U824 ( .A(n1230), .Y(n2148) );
  BUFX2 U825 ( .A(n2045), .Y(n1231) );
  INVX1 U826 ( .A(n1231), .Y(n2149) );
  BUFX2 U827 ( .A(n2142), .Y(n1232) );
  INVX1 U828 ( .A(n1232), .Y(n2143) );
  BUFX2 U829 ( .A(n2144), .Y(n1233) );
  INVX1 U830 ( .A(n1233), .Y(n2150) );
  AND2X1 U831 ( .A(n1852), .B(n1225), .Y(n1234) );
  AND2X1 U832 ( .A(n1817), .B(n1226), .Y(n1235) );
  INVX4 U833 ( .A(n3), .Y(n1904) );
  AND2X1 U834 ( .A(n1938), .B(n1225), .Y(n1236) );
  AND2X1 U835 ( .A(n1943), .B(n1226), .Y(n1237) );
  AND2X1 U836 ( .A(n1235), .B(n2151), .Y(n1238) );
  AND2X1 U837 ( .A(n2151), .B(n1237), .Y(n1239) );
  AND2X1 U838 ( .A(n2151), .B(n2143), .Y(n1240) );
  AND2X1 U839 ( .A(n2151), .B(n2150), .Y(n1241) );
  AND2X1 U840 ( .A(n1234), .B(n1235), .Y(n1242) );
  INVX1 U841 ( .A(n1242), .Y(n1243) );
  AND2X1 U842 ( .A(n1235), .B(n1236), .Y(n1245) );
  INVX1 U843 ( .A(n1245), .Y(n1246) );
  AND2X1 U844 ( .A(n1235), .B(n2145), .Y(n1248) );
  INVX1 U845 ( .A(n1248), .Y(n1249) );
  INVX1 U846 ( .A(n22), .Y(n1250) );
  INVX1 U847 ( .A(n22), .Y(n1251) );
  AND2X1 U848 ( .A(n1235), .B(n2146), .Y(n1252) );
  INVX1 U849 ( .A(n1252), .Y(n1253) );
  INVX1 U850 ( .A(n23), .Y(n1254) );
  INVX1 U851 ( .A(n23), .Y(n1255) );
  AND2X1 U852 ( .A(n1235), .B(n2147), .Y(n1256) );
  INVX1 U853 ( .A(n1256), .Y(n1257) );
  INVX1 U854 ( .A(n24), .Y(n1258) );
  INVX1 U855 ( .A(n24), .Y(n1259) );
  AND2X1 U856 ( .A(n1235), .B(n2148), .Y(n1260) );
  INVX1 U857 ( .A(n1260), .Y(n1261) );
  INVX1 U858 ( .A(n25), .Y(n1262) );
  INVX1 U859 ( .A(n25), .Y(n1263) );
  AND2X1 U860 ( .A(n1235), .B(n2149), .Y(n1264) );
  INVX1 U861 ( .A(n1264), .Y(n1265) );
  INVX1 U862 ( .A(n26), .Y(n1266) );
  INVX1 U863 ( .A(n26), .Y(n1267) );
  INVX1 U864 ( .A(n27), .Y(n1268) );
  INVX1 U865 ( .A(n27), .Y(n1269) );
  AND2X1 U866 ( .A(n1234), .B(n1237), .Y(n1270) );
  INVX1 U867 ( .A(n1270), .Y(n1271) );
  INVX1 U868 ( .A(n28), .Y(n1272) );
  INVX1 U869 ( .A(n28), .Y(n1273) );
  AND2X1 U870 ( .A(n1236), .B(n1237), .Y(n1274) );
  INVX1 U871 ( .A(n1274), .Y(n1275) );
  INVX1 U872 ( .A(n29), .Y(n1276) );
  INVX1 U873 ( .A(n29), .Y(n1277) );
  AND2X1 U874 ( .A(n2145), .B(n1237), .Y(n1278) );
  INVX1 U875 ( .A(n1278), .Y(n1279) );
  INVX1 U876 ( .A(n30), .Y(n1280) );
  INVX1 U877 ( .A(n30), .Y(n1281) );
  AND2X1 U878 ( .A(n2146), .B(n1237), .Y(n1282) );
  INVX1 U879 ( .A(n1282), .Y(n1283) );
  INVX1 U880 ( .A(n31), .Y(n1284) );
  INVX1 U881 ( .A(n31), .Y(n1285) );
  AND2X1 U882 ( .A(n2147), .B(n1237), .Y(n1286) );
  INVX1 U883 ( .A(n1286), .Y(n1287) );
  AND2X1 U884 ( .A(n2148), .B(n1237), .Y(n1288) );
  INVX1 U885 ( .A(n1288), .Y(n1289) );
  AND2X1 U886 ( .A(n2149), .B(n1237), .Y(n1290) );
  INVX1 U887 ( .A(n1290), .Y(n1291) );
  AND2X1 U888 ( .A(n1234), .B(n2143), .Y(n1292) );
  INVX1 U889 ( .A(n1292), .Y(n1293) );
  AND2X1 U890 ( .A(n1236), .B(n2143), .Y(n1294) );
  INVX1 U891 ( .A(n1294), .Y(n1295) );
  AND2X1 U892 ( .A(n2145), .B(n2143), .Y(n1296) );
  INVX1 U893 ( .A(n1296), .Y(n1297) );
  AND2X1 U894 ( .A(n2146), .B(n2143), .Y(n1298) );
  INVX1 U895 ( .A(n1298), .Y(n1299) );
  AND2X1 U896 ( .A(n2147), .B(n2143), .Y(n1300) );
  INVX1 U897 ( .A(n1300), .Y(n1301) );
  AND2X1 U898 ( .A(n2148), .B(n2143), .Y(n1302) );
  INVX1 U899 ( .A(n1302), .Y(n1303) );
  AND2X1 U900 ( .A(n2149), .B(n2143), .Y(n1304) );
  INVX1 U901 ( .A(n1304), .Y(n1305) );
  AND2X1 U902 ( .A(n1234), .B(n2150), .Y(n1306) );
  INVX1 U903 ( .A(n1306), .Y(n1307) );
  AND2X1 U904 ( .A(n1236), .B(n2150), .Y(n1308) );
  INVX1 U905 ( .A(n1308), .Y(n1309) );
  AND2X1 U906 ( .A(n2145), .B(n2150), .Y(n1310) );
  INVX1 U907 ( .A(n1310), .Y(n1311) );
  AND2X1 U908 ( .A(n2146), .B(n2150), .Y(n1312) );
  INVX1 U909 ( .A(n1312), .Y(n1313) );
  AND2X1 U910 ( .A(n2147), .B(n2150), .Y(n1314) );
  INVX1 U911 ( .A(n1314), .Y(n1315) );
  AND2X1 U912 ( .A(n2148), .B(n2150), .Y(n1316) );
  INVX1 U913 ( .A(n1316), .Y(n1317) );
  AND2X1 U914 ( .A(n2149), .B(n2150), .Y(n1318) );
  INVX1 U915 ( .A(n1318), .Y(n1319) );
  MUX2X1 U916 ( .B(n1321), .A(n1322), .S(n1825), .Y(n1320) );
  MUX2X1 U917 ( .B(n1324), .A(n1325), .S(n1825), .Y(n1323) );
  MUX2X1 U918 ( .B(n1327), .A(n1328), .S(n1825), .Y(n1326) );
  MUX2X1 U919 ( .B(n1330), .A(n1331), .S(n1825), .Y(n1329) );
  MUX2X1 U920 ( .B(n1333), .A(n1334), .S(n1818), .Y(n1332) );
  MUX2X1 U921 ( .B(n1336), .A(n1337), .S(n1825), .Y(n1335) );
  MUX2X1 U922 ( .B(n1339), .A(n1340), .S(n1825), .Y(n1338) );
  MUX2X1 U923 ( .B(n1342), .A(n1343), .S(n1825), .Y(n1341) );
  MUX2X1 U924 ( .B(n1345), .A(n1346), .S(n1825), .Y(n1344) );
  MUX2X1 U925 ( .B(n1348), .A(n1349), .S(n1818), .Y(n1347) );
  MUX2X1 U926 ( .B(n1351), .A(n1352), .S(n1826), .Y(n1350) );
  MUX2X1 U927 ( .B(n1354), .A(n1355), .S(n1826), .Y(n1353) );
  MUX2X1 U928 ( .B(n1357), .A(n1358), .S(n1826), .Y(n1356) );
  MUX2X1 U929 ( .B(n1360), .A(n1361), .S(n1826), .Y(n1359) );
  MUX2X1 U930 ( .B(n1363), .A(n1364), .S(n1818), .Y(n1362) );
  MUX2X1 U931 ( .B(n1366), .A(n1367), .S(n1826), .Y(n1365) );
  MUX2X1 U932 ( .B(n1369), .A(n1370), .S(n1826), .Y(n1368) );
  MUX2X1 U933 ( .B(n1372), .A(n1373), .S(n1826), .Y(n1371) );
  MUX2X1 U934 ( .B(n1375), .A(n1376), .S(n1826), .Y(n1374) );
  MUX2X1 U935 ( .B(n1378), .A(n1379), .S(n1818), .Y(n1377) );
  MUX2X1 U936 ( .B(n1381), .A(n1382), .S(n1826), .Y(n1380) );
  MUX2X1 U937 ( .B(n1384), .A(n1385), .S(n1826), .Y(n1383) );
  MUX2X1 U938 ( .B(n1387), .A(n1388), .S(n1826), .Y(n1386) );
  MUX2X1 U939 ( .B(n1390), .A(n1391), .S(n1826), .Y(n1389) );
  MUX2X1 U940 ( .B(n1393), .A(n1394), .S(n1818), .Y(n1392) );
  MUX2X1 U941 ( .B(n1396), .A(n1397), .S(n1827), .Y(n1395) );
  MUX2X1 U942 ( .B(n1399), .A(n1400), .S(n1827), .Y(n1398) );
  MUX2X1 U943 ( .B(n1402), .A(n1403), .S(n1827), .Y(n1401) );
  MUX2X1 U944 ( .B(n1405), .A(n1406), .S(n1827), .Y(n1404) );
  MUX2X1 U945 ( .B(n1408), .A(n1409), .S(n1818), .Y(n1407) );
  MUX2X1 U946 ( .B(n1411), .A(n1412), .S(n1827), .Y(n1410) );
  MUX2X1 U947 ( .B(n1414), .A(n1415), .S(n1827), .Y(n1413) );
  MUX2X1 U948 ( .B(n1417), .A(n1418), .S(n1827), .Y(n1416) );
  MUX2X1 U949 ( .B(n1420), .A(n1421), .S(n1827), .Y(n1419) );
  MUX2X1 U950 ( .B(n1423), .A(n1424), .S(n1818), .Y(n1422) );
  MUX2X1 U951 ( .B(n1426), .A(n1427), .S(n1827), .Y(n1425) );
  MUX2X1 U952 ( .B(n1429), .A(n1430), .S(n1827), .Y(n1428) );
  MUX2X1 U953 ( .B(n1432), .A(n1433), .S(n1827), .Y(n1431) );
  MUX2X1 U954 ( .B(n1435), .A(n1436), .S(n1827), .Y(n1434) );
  MUX2X1 U955 ( .B(n1438), .A(n1439), .S(n1818), .Y(n1437) );
  MUX2X1 U956 ( .B(n1441), .A(n1442), .S(n1828), .Y(n1440) );
  MUX2X1 U957 ( .B(n1444), .A(n1445), .S(n1828), .Y(n1443) );
  MUX2X1 U958 ( .B(n1447), .A(n1448), .S(n1828), .Y(n1446) );
  MUX2X1 U959 ( .B(n1450), .A(n1451), .S(n1828), .Y(n1449) );
  MUX2X1 U960 ( .B(n1453), .A(n1454), .S(n1818), .Y(n1452) );
  MUX2X1 U961 ( .B(n1456), .A(n1457), .S(n1828), .Y(n1455) );
  MUX2X1 U962 ( .B(n1459), .A(n1460), .S(n1828), .Y(n1458) );
  MUX2X1 U963 ( .B(n1462), .A(n1463), .S(n1828), .Y(n1461) );
  MUX2X1 U964 ( .B(n1465), .A(n1466), .S(n1828), .Y(n1464) );
  MUX2X1 U965 ( .B(n1468), .A(n1469), .S(n1818), .Y(n1467) );
  MUX2X1 U966 ( .B(n1471), .A(n1472), .S(n1828), .Y(n1470) );
  MUX2X1 U967 ( .B(n1474), .A(n1475), .S(n1828), .Y(n1473) );
  MUX2X1 U968 ( .B(n1477), .A(n1478), .S(n1828), .Y(n1476) );
  MUX2X1 U969 ( .B(n1480), .A(n1481), .S(n1828), .Y(n1479) );
  MUX2X1 U970 ( .B(n1483), .A(n1484), .S(n1818), .Y(n1482) );
  MUX2X1 U971 ( .B(n1486), .A(n1487), .S(n1829), .Y(n1485) );
  MUX2X1 U972 ( .B(n1489), .A(n1490), .S(n1829), .Y(n1488) );
  MUX2X1 U973 ( .B(n1492), .A(n1493), .S(n1829), .Y(n1491) );
  MUX2X1 U974 ( .B(n1495), .A(n1496), .S(n1829), .Y(n1494) );
  MUX2X1 U975 ( .B(n1498), .A(n1499), .S(n1818), .Y(n1497) );
  MUX2X1 U976 ( .B(n1501), .A(n1502), .S(n1829), .Y(n1500) );
  MUX2X1 U977 ( .B(n1504), .A(n1505), .S(n1829), .Y(n1503) );
  MUX2X1 U978 ( .B(n1507), .A(n1508), .S(n1829), .Y(n1506) );
  MUX2X1 U979 ( .B(n1510), .A(n1511), .S(n1829), .Y(n1509) );
  MUX2X1 U980 ( .B(n1513), .A(n1514), .S(n1818), .Y(n1512) );
  MUX2X1 U981 ( .B(n1516), .A(n1517), .S(n1829), .Y(n1515) );
  MUX2X1 U982 ( .B(n1519), .A(n1520), .S(n1829), .Y(n1518) );
  MUX2X1 U983 ( .B(n1522), .A(n1523), .S(n1829), .Y(n1521) );
  MUX2X1 U984 ( .B(n1525), .A(n1526), .S(n1829), .Y(n1524) );
  MUX2X1 U985 ( .B(n1528), .A(n1529), .S(n1818), .Y(n1527) );
  MUX2X1 U986 ( .B(n1531), .A(n1532), .S(n1830), .Y(n1530) );
  MUX2X1 U987 ( .B(n1534), .A(n1535), .S(n1830), .Y(n1533) );
  MUX2X1 U988 ( .B(n1537), .A(n1538), .S(n1830), .Y(n1536) );
  MUX2X1 U989 ( .B(n1540), .A(n1541), .S(n1830), .Y(n1539) );
  MUX2X1 U990 ( .B(n1543), .A(n1544), .S(n1817), .Y(n1542) );
  MUX2X1 U991 ( .B(n1546), .A(n1547), .S(n1830), .Y(n1545) );
  MUX2X1 U992 ( .B(n1549), .A(n1550), .S(n1830), .Y(n1548) );
  MUX2X1 U993 ( .B(n1552), .A(n1553), .S(n1830), .Y(n1551) );
  MUX2X1 U994 ( .B(n1555), .A(n1556), .S(n1830), .Y(n1554) );
  MUX2X1 U995 ( .B(n1558), .A(n1559), .S(n1817), .Y(n1557) );
  MUX2X1 U996 ( .B(n1561), .A(n1562), .S(n1830), .Y(n1560) );
  MUX2X1 U997 ( .B(n1564), .A(n1565), .S(n1830), .Y(n1563) );
  MUX2X1 U998 ( .B(n1567), .A(n1568), .S(n1830), .Y(n1566) );
  MUX2X1 U999 ( .B(n1570), .A(n1571), .S(n1830), .Y(n1569) );
  MUX2X1 U1000 ( .B(n1573), .A(n1574), .S(n1817), .Y(n1572) );
  MUX2X1 U1001 ( .B(n1576), .A(n1577), .S(n1831), .Y(n1575) );
  MUX2X1 U1002 ( .B(n1579), .A(n1580), .S(n1831), .Y(n1578) );
  MUX2X1 U1003 ( .B(n1582), .A(n1583), .S(n1831), .Y(n1581) );
  MUX2X1 U1004 ( .B(n1585), .A(n1586), .S(n1831), .Y(n1584) );
  MUX2X1 U1005 ( .B(n1588), .A(n1589), .S(n1817), .Y(n1587) );
  MUX2X1 U1006 ( .B(n1591), .A(n1592), .S(n1831), .Y(n1590) );
  MUX2X1 U1007 ( .B(n1594), .A(n1595), .S(n1831), .Y(n1593) );
  MUX2X1 U1008 ( .B(n1597), .A(n1598), .S(n1831), .Y(n1596) );
  MUX2X1 U1009 ( .B(n1600), .A(n1601), .S(n1831), .Y(n1599) );
  MUX2X1 U1010 ( .B(n1603), .A(n1604), .S(n1818), .Y(n1602) );
  MUX2X1 U1011 ( .B(n1606), .A(n1607), .S(n1831), .Y(n1605) );
  MUX2X1 U1012 ( .B(n1609), .A(n1610), .S(n1831), .Y(n1608) );
  MUX2X1 U1013 ( .B(n1612), .A(n1613), .S(n1831), .Y(n1611) );
  MUX2X1 U1014 ( .B(n1615), .A(n1616), .S(n1831), .Y(n1614) );
  MUX2X1 U1015 ( .B(n1618), .A(n1619), .S(n1817), .Y(n1617) );
  MUX2X1 U1016 ( .B(n1621), .A(n1622), .S(n1832), .Y(n1620) );
  MUX2X1 U1017 ( .B(n1624), .A(n1625), .S(n1832), .Y(n1623) );
  MUX2X1 U1018 ( .B(n1627), .A(n1628), .S(n1832), .Y(n1626) );
  MUX2X1 U1019 ( .B(n1630), .A(n1631), .S(n1832), .Y(n1629) );
  MUX2X1 U1020 ( .B(n1633), .A(n1634), .S(n1817), .Y(n1632) );
  MUX2X1 U1021 ( .B(n1636), .A(n1637), .S(n1832), .Y(n1635) );
  MUX2X1 U1022 ( .B(n1639), .A(n1640), .S(n1832), .Y(n1638) );
  MUX2X1 U1023 ( .B(n1642), .A(n1643), .S(n1832), .Y(n1641) );
  MUX2X1 U1024 ( .B(n1645), .A(n1646), .S(n1832), .Y(n1644) );
  MUX2X1 U1025 ( .B(n1648), .A(n1649), .S(n1817), .Y(n1647) );
  MUX2X1 U1026 ( .B(n1651), .A(n1652), .S(n1832), .Y(n1650) );
  MUX2X1 U1027 ( .B(n1654), .A(n1655), .S(n1832), .Y(n1653) );
  MUX2X1 U1028 ( .B(n1657), .A(n1658), .S(n1832), .Y(n1656) );
  MUX2X1 U1029 ( .B(n1660), .A(n1661), .S(n1832), .Y(n1659) );
  MUX2X1 U1030 ( .B(n1663), .A(n1664), .S(n1818), .Y(n1662) );
  MUX2X1 U1031 ( .B(n1666), .A(n1667), .S(n1833), .Y(n1665) );
  MUX2X1 U1032 ( .B(n1669), .A(n1670), .S(n1833), .Y(n1668) );
  MUX2X1 U1033 ( .B(n1672), .A(n1673), .S(n1833), .Y(n1671) );
  MUX2X1 U1034 ( .B(n1675), .A(n1676), .S(n1833), .Y(n1674) );
  MUX2X1 U1035 ( .B(n1678), .A(n1679), .S(n1818), .Y(n1677) );
  MUX2X1 U1036 ( .B(n1681), .A(n1682), .S(n1833), .Y(n1680) );
  MUX2X1 U1037 ( .B(n1684), .A(n1685), .S(n1833), .Y(n1683) );
  MUX2X1 U1038 ( .B(n1687), .A(n1688), .S(n1833), .Y(n1686) );
  MUX2X1 U1039 ( .B(n1690), .A(n1691), .S(n1833), .Y(n1689) );
  MUX2X1 U1040 ( .B(n1693), .A(n1694), .S(n1817), .Y(n1692) );
  MUX2X1 U1041 ( .B(n1696), .A(n1697), .S(n1833), .Y(n1695) );
  MUX2X1 U1042 ( .B(n1699), .A(n1700), .S(n1833), .Y(n1698) );
  MUX2X1 U1043 ( .B(n1702), .A(n1703), .S(n1833), .Y(n1701) );
  MUX2X1 U1044 ( .B(n1705), .A(n1706), .S(n1833), .Y(n1704) );
  MUX2X1 U1045 ( .B(n1708), .A(n1709), .S(n1817), .Y(n1707) );
  MUX2X1 U1046 ( .B(n1711), .A(n1712), .S(n1834), .Y(n1710) );
  MUX2X1 U1047 ( .B(n1714), .A(n1715), .S(n1834), .Y(n1713) );
  MUX2X1 U1048 ( .B(n1717), .A(n1718), .S(n1834), .Y(n1716) );
  MUX2X1 U1049 ( .B(n1720), .A(n1721), .S(n1834), .Y(n1719) );
  MUX2X1 U1050 ( .B(n1723), .A(n1724), .S(n1817), .Y(n1722) );
  MUX2X1 U1051 ( .B(n1726), .A(n1727), .S(n1834), .Y(n1725) );
  MUX2X1 U1052 ( .B(n1729), .A(n1730), .S(n1834), .Y(n1728) );
  MUX2X1 U1053 ( .B(n1732), .A(n1733), .S(n1834), .Y(n1731) );
  MUX2X1 U1054 ( .B(n1735), .A(n1736), .S(n1834), .Y(n1734) );
  MUX2X1 U1055 ( .B(n1738), .A(n1739), .S(n1817), .Y(n1737) );
  MUX2X1 U1056 ( .B(n1741), .A(n1742), .S(n1834), .Y(n1740) );
  MUX2X1 U1057 ( .B(n1744), .A(n1745), .S(n1834), .Y(n1743) );
  MUX2X1 U1058 ( .B(n1747), .A(n1748), .S(n1834), .Y(n1746) );
  MUX2X1 U1059 ( .B(n1750), .A(n1751), .S(n1834), .Y(n1749) );
  MUX2X1 U1060 ( .B(n1753), .A(n1754), .S(n1817), .Y(n1752) );
  MUX2X1 U1061 ( .B(n1756), .A(n1757), .S(n1835), .Y(n1755) );
  MUX2X1 U1062 ( .B(n1759), .A(n1760), .S(n1835), .Y(n1758) );
  MUX2X1 U1063 ( .B(n1762), .A(n1763), .S(n1835), .Y(n1761) );
  MUX2X1 U1064 ( .B(n1765), .A(n1766), .S(n1835), .Y(n1764) );
  MUX2X1 U1065 ( .B(n1768), .A(n1769), .S(n1817), .Y(n1767) );
  MUX2X1 U1066 ( .B(n1771), .A(n1772), .S(n1835), .Y(n1770) );
  MUX2X1 U1067 ( .B(n1774), .A(n1775), .S(n1835), .Y(n1773) );
  MUX2X1 U1068 ( .B(n1777), .A(n1778), .S(n1835), .Y(n1776) );
  MUX2X1 U1069 ( .B(n1780), .A(n1781), .S(n1835), .Y(n1779) );
  MUX2X1 U1070 ( .B(n1783), .A(n1784), .S(n1817), .Y(n1782) );
  MUX2X1 U1071 ( .B(n1786), .A(n1787), .S(n1835), .Y(n1785) );
  MUX2X1 U1072 ( .B(n1789), .A(n1790), .S(n1835), .Y(n1788) );
  MUX2X1 U1073 ( .B(n1792), .A(n1793), .S(n1835), .Y(n1791) );
  MUX2X1 U1074 ( .B(n1795), .A(n1796), .S(n1835), .Y(n1794) );
  MUX2X1 U1075 ( .B(n1798), .A(n1799), .S(n1817), .Y(n1797) );
  MUX2X1 U1076 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n1853), .Y(n1322) );
  MUX2X1 U1077 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1851), .Y(n1321) );
  MUX2X1 U1078 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n1844), .Y(n1325) );
  MUX2X1 U1079 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n1843), .Y(n1324) );
  MUX2X1 U1080 ( .B(n1323), .A(n1320), .S(n1822), .Y(n1334) );
  MUX2X1 U1081 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1841), .Y(n1328) );
  MUX2X1 U1082 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1841), .Y(n1327) );
  MUX2X1 U1083 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n1841), .Y(n1331) );
  MUX2X1 U1084 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n1841), .Y(n1330) );
  MUX2X1 U1085 ( .B(n1329), .A(n1326), .S(n1822), .Y(n1333) );
  MUX2X1 U1086 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n1841), .Y(n1337) );
  MUX2X1 U1087 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n1841), .Y(n1336) );
  MUX2X1 U1088 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n1841), .Y(n1340) );
  MUX2X1 U1089 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n1841), .Y(n1339) );
  MUX2X1 U1090 ( .B(n1338), .A(n1335), .S(n1822), .Y(n1349) );
  MUX2X1 U1091 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n1841), .Y(n1343) );
  MUX2X1 U1092 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n1841), .Y(n1342) );
  MUX2X1 U1093 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n1841), .Y(n1346) );
  MUX2X1 U1094 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n1841), .Y(n1345) );
  MUX2X1 U1095 ( .B(n1344), .A(n1341), .S(n1822), .Y(n1348) );
  MUX2X1 U1096 ( .B(n1347), .A(n1332), .S(n1816), .Y(n1800) );
  MUX2X1 U1097 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n1842), .Y(n1352) );
  MUX2X1 U1098 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n1842), .Y(n1351) );
  MUX2X1 U1099 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n1842), .Y(n1355) );
  MUX2X1 U1100 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n1842), .Y(n1354) );
  MUX2X1 U1101 ( .B(n1353), .A(n1350), .S(n1822), .Y(n1364) );
  MUX2X1 U1102 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n1842), .Y(n1358) );
  MUX2X1 U1103 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n1842), .Y(n1357) );
  MUX2X1 U1104 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n1842), .Y(n1361) );
  MUX2X1 U1105 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n1842), .Y(n1360) );
  MUX2X1 U1106 ( .B(n1359), .A(n1356), .S(n1822), .Y(n1363) );
  MUX2X1 U1107 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n1842), .Y(n1367) );
  MUX2X1 U1108 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n1842), .Y(n1366) );
  MUX2X1 U1109 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n1842), .Y(n1370) );
  MUX2X1 U1110 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n1842), .Y(n1369) );
  MUX2X1 U1111 ( .B(n1368), .A(n1365), .S(n1822), .Y(n1379) );
  MUX2X1 U1112 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n1843), .Y(n1373) );
  MUX2X1 U1113 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n1843), .Y(n1372) );
  MUX2X1 U1114 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n1843), .Y(n1376) );
  MUX2X1 U1115 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n1843), .Y(n1375) );
  MUX2X1 U1116 ( .B(n1374), .A(n1371), .S(n1822), .Y(n1378) );
  MUX2X1 U1117 ( .B(n1377), .A(n1362), .S(n1816), .Y(n1801) );
  MUX2X1 U1118 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n1843), .Y(n1382) );
  MUX2X1 U1119 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n1843), .Y(n1381) );
  MUX2X1 U1120 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n1843), .Y(n1385) );
  MUX2X1 U1121 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n1843), .Y(n1384) );
  MUX2X1 U1122 ( .B(n1383), .A(n1380), .S(n1822), .Y(n1394) );
  MUX2X1 U1123 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n1843), .Y(n1388) );
  MUX2X1 U1124 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n1843), .Y(n1387) );
  MUX2X1 U1125 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n1843), .Y(n1391) );
  MUX2X1 U1126 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n1843), .Y(n1390) );
  MUX2X1 U1127 ( .B(n1389), .A(n1386), .S(n1822), .Y(n1393) );
  MUX2X1 U1128 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n1844), .Y(n1397) );
  MUX2X1 U1129 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n1844), .Y(n1396) );
  MUX2X1 U1130 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n1844), .Y(n1400) );
  MUX2X1 U1131 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n1844), .Y(n1399) );
  MUX2X1 U1132 ( .B(n1398), .A(n1395), .S(n1822), .Y(n1409) );
  MUX2X1 U1133 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n1844), .Y(n1403) );
  MUX2X1 U1134 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n1844), .Y(n1402) );
  MUX2X1 U1135 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n1844), .Y(n1406) );
  MUX2X1 U1136 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n1844), .Y(n1405) );
  MUX2X1 U1137 ( .B(n1404), .A(n1401), .S(n1822), .Y(n1408) );
  MUX2X1 U1138 ( .B(n1407), .A(n1392), .S(n1816), .Y(n1802) );
  MUX2X1 U1139 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n1844), .Y(n1412) );
  MUX2X1 U1140 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n1844), .Y(n1411) );
  MUX2X1 U1141 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n1844), .Y(n1415) );
  MUX2X1 U1142 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n1844), .Y(n1414) );
  MUX2X1 U1143 ( .B(n1413), .A(n1410), .S(n1821), .Y(n1424) );
  MUX2X1 U1144 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n1845), .Y(n1418) );
  MUX2X1 U1145 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n1845), .Y(n1417) );
  MUX2X1 U1146 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n1845), .Y(n1421) );
  MUX2X1 U1147 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n1845), .Y(n1420) );
  MUX2X1 U1148 ( .B(n1419), .A(n1416), .S(n1821), .Y(n1423) );
  MUX2X1 U1149 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n1845), .Y(n1427) );
  MUX2X1 U1150 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n1845), .Y(n1426) );
  MUX2X1 U1151 ( .B(\mem<10><3> ), .A(\mem<11><3> ), .S(n1845), .Y(n1430) );
  MUX2X1 U1152 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n1845), .Y(n1429) );
  MUX2X1 U1153 ( .B(n1428), .A(n1425), .S(n1821), .Y(n1439) );
  MUX2X1 U1154 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n1845), .Y(n1433) );
  MUX2X1 U1155 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n1845), .Y(n1432) );
  MUX2X1 U1156 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n1845), .Y(n1436) );
  MUX2X1 U1157 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n1845), .Y(n1435) );
  MUX2X1 U1158 ( .B(n1434), .A(n1431), .S(n1821), .Y(n1438) );
  MUX2X1 U1159 ( .B(n1437), .A(n1422), .S(n1816), .Y(n1803) );
  MUX2X1 U1160 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n1846), .Y(n1442) );
  MUX2X1 U1161 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n1846), .Y(n1441) );
  MUX2X1 U1162 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n1846), .Y(n1445) );
  MUX2X1 U1163 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n1846), .Y(n1444) );
  MUX2X1 U1164 ( .B(n1443), .A(n1440), .S(n1821), .Y(n1454) );
  MUX2X1 U1165 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n1846), .Y(n1448) );
  MUX2X1 U1166 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n1846), .Y(n1447) );
  MUX2X1 U1167 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n1846), .Y(n1451) );
  MUX2X1 U1168 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n1846), .Y(n1450) );
  MUX2X1 U1169 ( .B(n1449), .A(n1446), .S(n1821), .Y(n1453) );
  MUX2X1 U1170 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n1846), .Y(n1457) );
  MUX2X1 U1171 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n1846), .Y(n1456) );
  MUX2X1 U1172 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n1846), .Y(n1460) );
  MUX2X1 U1173 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n1846), .Y(n1459) );
  MUX2X1 U1174 ( .B(n1458), .A(n1455), .S(n1821), .Y(n1469) );
  MUX2X1 U1175 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n1847), .Y(n1463) );
  MUX2X1 U1177 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n1847), .Y(n1462) );
  MUX2X1 U1178 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n1847), .Y(n1466) );
  MUX2X1 U1179 ( .B(\mem<0><4> ), .A(\mem<1><4> ), .S(n1847), .Y(n1465) );
  MUX2X1 U1180 ( .B(n1464), .A(n1461), .S(n1821), .Y(n1468) );
  MUX2X1 U1181 ( .B(n1467), .A(n1452), .S(n1816), .Y(n1804) );
  MUX2X1 U1182 ( .B(\mem<30><5> ), .A(\mem<31><5> ), .S(n1847), .Y(n1472) );
  MUX2X1 U1183 ( .B(\mem<28><5> ), .A(\mem<29><5> ), .S(n1847), .Y(n1471) );
  MUX2X1 U1184 ( .B(\mem<26><5> ), .A(\mem<27><5> ), .S(n1847), .Y(n1475) );
  MUX2X1 U1185 ( .B(\mem<24><5> ), .A(\mem<25><5> ), .S(n1847), .Y(n1474) );
  MUX2X1 U1186 ( .B(n1473), .A(n1470), .S(n1821), .Y(n1484) );
  MUX2X1 U1187 ( .B(\mem<22><5> ), .A(\mem<23><5> ), .S(n1847), .Y(n1478) );
  MUX2X1 U1188 ( .B(\mem<20><5> ), .A(\mem<21><5> ), .S(n1847), .Y(n1477) );
  MUX2X1 U1189 ( .B(\mem<18><5> ), .A(\mem<19><5> ), .S(n1847), .Y(n1481) );
  MUX2X1 U1190 ( .B(\mem<16><5> ), .A(\mem<17><5> ), .S(n1847), .Y(n1480) );
  MUX2X1 U1191 ( .B(n1479), .A(n1476), .S(n1821), .Y(n1483) );
  MUX2X1 U1192 ( .B(\mem<14><5> ), .A(\mem<15><5> ), .S(n1847), .Y(n1487) );
  MUX2X1 U1193 ( .B(\mem<12><5> ), .A(\mem<13><5> ), .S(n1846), .Y(n1486) );
  MUX2X1 U1194 ( .B(\mem<10><5> ), .A(\mem<11><5> ), .S(n1851), .Y(n1490) );
  MUX2X1 U1195 ( .B(\mem<8><5> ), .A(\mem<9><5> ), .S(n1851), .Y(n1489) );
  MUX2X1 U1196 ( .B(n1488), .A(n1485), .S(n1821), .Y(n1499) );
  MUX2X1 U1197 ( .B(\mem<6><5> ), .A(\mem<7><5> ), .S(n1845), .Y(n1493) );
  MUX2X1 U1198 ( .B(\mem<4><5> ), .A(\mem<5><5> ), .S(n1844), .Y(n1492) );
  MUX2X1 U1199 ( .B(\mem<2><5> ), .A(\mem<3><5> ), .S(n1850), .Y(n1496) );
  MUX2X1 U1200 ( .B(\mem<0><5> ), .A(\mem<1><5> ), .S(n1841), .Y(n1495) );
  MUX2X1 U1201 ( .B(n1494), .A(n1491), .S(n1821), .Y(n1498) );
  MUX2X1 U1202 ( .B(n1497), .A(n1482), .S(n1816), .Y(n1805) );
  MUX2X1 U1203 ( .B(\mem<30><6> ), .A(\mem<31><6> ), .S(n1846), .Y(n1502) );
  MUX2X1 U1204 ( .B(\mem<28><6> ), .A(\mem<29><6> ), .S(n1847), .Y(n1501) );
  MUX2X1 U1205 ( .B(\mem<26><6> ), .A(\mem<27><6> ), .S(n1843), .Y(n1505) );
  MUX2X1 U1206 ( .B(\mem<24><6> ), .A(\mem<25><6> ), .S(n1847), .Y(n1504) );
  MUX2X1 U1207 ( .B(n1503), .A(n1500), .S(n1820), .Y(n1514) );
  MUX2X1 U1208 ( .B(\mem<22><6> ), .A(\mem<23><6> ), .S(n1848), .Y(n1508) );
  MUX2X1 U1209 ( .B(\mem<20><6> ), .A(\mem<21><6> ), .S(n1848), .Y(n1507) );
  MUX2X1 U1210 ( .B(\mem<18><6> ), .A(\mem<19><6> ), .S(n1848), .Y(n1511) );
  MUX2X1 U1211 ( .B(\mem<16><6> ), .A(\mem<17><6> ), .S(n1848), .Y(n1510) );
  MUX2X1 U1212 ( .B(n1509), .A(n1506), .S(n1820), .Y(n1513) );
  MUX2X1 U1213 ( .B(\mem<14><6> ), .A(\mem<15><6> ), .S(n1848), .Y(n1517) );
  MUX2X1 U1214 ( .B(\mem<12><6> ), .A(\mem<13><6> ), .S(n1848), .Y(n1516) );
  MUX2X1 U1215 ( .B(\mem<10><6> ), .A(\mem<11><6> ), .S(n1848), .Y(n1520) );
  MUX2X1 U1216 ( .B(\mem<8><6> ), .A(\mem<9><6> ), .S(n1848), .Y(n1519) );
  MUX2X1 U1217 ( .B(n1518), .A(n1515), .S(n1820), .Y(n1529) );
  MUX2X1 U1218 ( .B(\mem<6><6> ), .A(\mem<7><6> ), .S(n1848), .Y(n1523) );
  MUX2X1 U1219 ( .B(\mem<4><6> ), .A(\mem<5><6> ), .S(n1848), .Y(n1522) );
  MUX2X1 U1220 ( .B(\mem<2><6> ), .A(\mem<3><6> ), .S(n1848), .Y(n1526) );
  MUX2X1 U1221 ( .B(\mem<0><6> ), .A(\mem<1><6> ), .S(n1848), .Y(n1525) );
  MUX2X1 U1222 ( .B(n1524), .A(n1521), .S(n1820), .Y(n1528) );
  MUX2X1 U1223 ( .B(n1527), .A(n1512), .S(n1816), .Y(n1806) );
  MUX2X1 U1224 ( .B(\mem<30><7> ), .A(\mem<31><7> ), .S(n1849), .Y(n1532) );
  MUX2X1 U1225 ( .B(\mem<28><7> ), .A(\mem<29><7> ), .S(n1849), .Y(n1531) );
  MUX2X1 U1226 ( .B(\mem<26><7> ), .A(\mem<27><7> ), .S(n1849), .Y(n1535) );
  MUX2X1 U1227 ( .B(\mem<24><7> ), .A(\mem<25><7> ), .S(n1849), .Y(n1534) );
  MUX2X1 U1228 ( .B(n1533), .A(n1530), .S(n1820), .Y(n1544) );
  MUX2X1 U1229 ( .B(\mem<22><7> ), .A(\mem<23><7> ), .S(n1849), .Y(n1538) );
  MUX2X1 U1230 ( .B(\mem<20><7> ), .A(\mem<21><7> ), .S(n1849), .Y(n1537) );
  MUX2X1 U1231 ( .B(\mem<18><7> ), .A(\mem<19><7> ), .S(n1849), .Y(n1541) );
  MUX2X1 U1232 ( .B(\mem<16><7> ), .A(\mem<17><7> ), .S(n1849), .Y(n1540) );
  MUX2X1 U1233 ( .B(n1539), .A(n1536), .S(n1820), .Y(n1543) );
  MUX2X1 U1234 ( .B(\mem<14><7> ), .A(\mem<15><7> ), .S(n1849), .Y(n1547) );
  MUX2X1 U1235 ( .B(\mem<12><7> ), .A(\mem<13><7> ), .S(n1849), .Y(n1546) );
  MUX2X1 U1236 ( .B(\mem<10><7> ), .A(\mem<11><7> ), .S(n1849), .Y(n1550) );
  MUX2X1 U1237 ( .B(\mem<8><7> ), .A(\mem<9><7> ), .S(n1849), .Y(n1549) );
  MUX2X1 U1238 ( .B(n1548), .A(n1545), .S(n1820), .Y(n1559) );
  MUX2X1 U1239 ( .B(\mem<6><7> ), .A(\mem<7><7> ), .S(n1848), .Y(n1553) );
  MUX2X1 U1240 ( .B(\mem<4><7> ), .A(\mem<5><7> ), .S(n1841), .Y(n1552) );
  MUX2X1 U1241 ( .B(\mem<2><7> ), .A(\mem<3><7> ), .S(n1848), .Y(n1556) );
  MUX2X1 U1242 ( .B(\mem<0><7> ), .A(\mem<1><7> ), .S(n1849), .Y(n1555) );
  MUX2X1 U1243 ( .B(n1554), .A(n1551), .S(n1820), .Y(n1558) );
  MUX2X1 U1244 ( .B(n1557), .A(n1542), .S(n1816), .Y(n1807) );
  MUX2X1 U1245 ( .B(\mem<30><8> ), .A(\mem<31><8> ), .S(n1841), .Y(n1562) );
  MUX2X1 U1246 ( .B(\mem<28><8> ), .A(\mem<29><8> ), .S(n1841), .Y(n1561) );
  MUX2X1 U1247 ( .B(\mem<26><8> ), .A(\mem<27><8> ), .S(n1847), .Y(n1565) );
  MUX2X1 U1248 ( .B(\mem<24><8> ), .A(\mem<25><8> ), .S(n1849), .Y(n1564) );
  MUX2X1 U1249 ( .B(n1563), .A(n1560), .S(n1820), .Y(n1574) );
  MUX2X1 U1250 ( .B(\mem<22><8> ), .A(\mem<23><8> ), .S(n1848), .Y(n1568) );
  MUX2X1 U1251 ( .B(\mem<20><8> ), .A(\mem<21><8> ), .S(n1847), .Y(n1567) );
  MUX2X1 U1252 ( .B(\mem<18><8> ), .A(\mem<19><8> ), .S(n1851), .Y(n1571) );
  MUX2X1 U1253 ( .B(\mem<16><8> ), .A(\mem<17><8> ), .S(n1856), .Y(n1570) );
  MUX2X1 U1254 ( .B(n1569), .A(n1566), .S(n1820), .Y(n1573) );
  MUX2X1 U1255 ( .B(\mem<14><8> ), .A(\mem<15><8> ), .S(n1849), .Y(n1577) );
  MUX2X1 U1256 ( .B(\mem<12><8> ), .A(\mem<13><8> ), .S(n1846), .Y(n1576) );
  MUX2X1 U1257 ( .B(\mem<10><8> ), .A(\mem<11><8> ), .S(n1847), .Y(n1580) );
  MUX2X1 U1258 ( .B(\mem<8><8> ), .A(\mem<9><8> ), .S(n1848), .Y(n1579) );
  MUX2X1 U1259 ( .B(n1578), .A(n1575), .S(n1820), .Y(n1589) );
  MUX2X1 U1260 ( .B(\mem<6><8> ), .A(\mem<7><8> ), .S(n1845), .Y(n1583) );
  MUX2X1 U1261 ( .B(\mem<4><8> ), .A(\mem<5><8> ), .S(n1851), .Y(n1582) );
  MUX2X1 U1262 ( .B(\mem<2><8> ), .A(\mem<3><8> ), .S(n1849), .Y(n1586) );
  MUX2X1 U1263 ( .B(\mem<0><8> ), .A(\mem<1><8> ), .S(n1846), .Y(n1585) );
  MUX2X1 U1264 ( .B(n1584), .A(n1581), .S(n1820), .Y(n1588) );
  MUX2X1 U1265 ( .B(n1587), .A(n1572), .S(n1816), .Y(n1808) );
  MUX2X1 U1266 ( .B(\mem<30><9> ), .A(\mem<31><9> ), .S(n1845), .Y(n1592) );
  MUX2X1 U1267 ( .B(\mem<28><9> ), .A(\mem<29><9> ), .S(n1848), .Y(n1591) );
  MUX2X1 U1268 ( .B(\mem<26><9> ), .A(\mem<27><9> ), .S(n1848), .Y(n1595) );
  MUX2X1 U1269 ( .B(\mem<24><9> ), .A(\mem<25><9> ), .S(n1848), .Y(n1594) );
  MUX2X1 U1270 ( .B(n1593), .A(n1590), .S(n1819), .Y(n1604) );
  MUX2X1 U1271 ( .B(\mem<22><9> ), .A(\mem<23><9> ), .S(n1850), .Y(n1598) );
  MUX2X1 U1272 ( .B(\mem<20><9> ), .A(\mem<21><9> ), .S(n1850), .Y(n1597) );
  MUX2X1 U1273 ( .B(\mem<18><9> ), .A(\mem<19><9> ), .S(n1850), .Y(n1601) );
  MUX2X1 U1274 ( .B(\mem<16><9> ), .A(\mem<17><9> ), .S(n1850), .Y(n1600) );
  MUX2X1 U1275 ( .B(n1599), .A(n1596), .S(n1819), .Y(n1603) );
  MUX2X1 U1276 ( .B(\mem<14><9> ), .A(\mem<15><9> ), .S(n1850), .Y(n1607) );
  MUX2X1 U1277 ( .B(\mem<12><9> ), .A(\mem<13><9> ), .S(n1850), .Y(n1606) );
  MUX2X1 U1278 ( .B(\mem<10><9> ), .A(\mem<11><9> ), .S(n1850), .Y(n1610) );
  MUX2X1 U1279 ( .B(\mem<8><9> ), .A(\mem<9><9> ), .S(n1850), .Y(n1609) );
  MUX2X1 U1280 ( .B(n1608), .A(n1605), .S(n1819), .Y(n1619) );
  MUX2X1 U1281 ( .B(\mem<6><9> ), .A(\mem<7><9> ), .S(n1850), .Y(n1613) );
  MUX2X1 U1282 ( .B(\mem<4><9> ), .A(\mem<5><9> ), .S(n1850), .Y(n1612) );
  MUX2X1 U1283 ( .B(\mem<2><9> ), .A(\mem<3><9> ), .S(n1850), .Y(n1616) );
  MUX2X1 U1284 ( .B(\mem<0><9> ), .A(\mem<1><9> ), .S(n1850), .Y(n1615) );
  MUX2X1 U1285 ( .B(n1614), .A(n1611), .S(n1819), .Y(n1618) );
  MUX2X1 U1286 ( .B(n1617), .A(n1602), .S(n1816), .Y(n1809) );
  MUX2X1 U1287 ( .B(\mem<30><10> ), .A(\mem<31><10> ), .S(n1851), .Y(n1622) );
  MUX2X1 U1288 ( .B(\mem<28><10> ), .A(\mem<29><10> ), .S(n1846), .Y(n1621) );
  MUX2X1 U1289 ( .B(\mem<26><10> ), .A(\mem<27><10> ), .S(n1845), .Y(n1625) );
  MUX2X1 U1290 ( .B(\mem<24><10> ), .A(\mem<25><10> ), .S(n1849), .Y(n1624) );
  MUX2X1 U1291 ( .B(n1623), .A(n1620), .S(n1819), .Y(n1634) );
  MUX2X1 U1292 ( .B(\mem<22><10> ), .A(\mem<23><10> ), .S(n1845), .Y(n1628) );
  MUX2X1 U1293 ( .B(\mem<20><10> ), .A(\mem<21><10> ), .S(n1849), .Y(n1627) );
  MUX2X1 U1294 ( .B(\mem<18><10> ), .A(\mem<19><10> ), .S(n1850), .Y(n1631) );
  MUX2X1 U1295 ( .B(\mem<16><10> ), .A(\mem<17><10> ), .S(n1847), .Y(n1630) );
  MUX2X1 U1296 ( .B(n1629), .A(n1626), .S(n1819), .Y(n1633) );
  MUX2X1 U1297 ( .B(\mem<14><10> ), .A(\mem<15><10> ), .S(n1846), .Y(n1637) );
  MUX2X1 U1298 ( .B(\mem<12><10> ), .A(\mem<13><10> ), .S(n1848), .Y(n1636) );
  MUX2X1 U1299 ( .B(\mem<10><10> ), .A(\mem<11><10> ), .S(n1846), .Y(n1640) );
  MUX2X1 U1300 ( .B(\mem<8><10> ), .A(\mem<9><10> ), .S(n1845), .Y(n1639) );
  MUX2X1 U1301 ( .B(n1638), .A(n1635), .S(n1819), .Y(n1649) );
  MUX2X1 U1302 ( .B(\mem<6><10> ), .A(\mem<7><10> ), .S(n1851), .Y(n1643) );
  MUX2X1 U1303 ( .B(\mem<4><10> ), .A(\mem<5><10> ), .S(n1851), .Y(n1642) );
  MUX2X1 U1304 ( .B(\mem<2><10> ), .A(\mem<3><10> ), .S(n1851), .Y(n1646) );
  MUX2X1 U1305 ( .B(\mem<0><10> ), .A(\mem<1><10> ), .S(n1851), .Y(n1645) );
  MUX2X1 U1306 ( .B(n1644), .A(n1641), .S(n1819), .Y(n1648) );
  MUX2X1 U1307 ( .B(n1647), .A(n1632), .S(n1816), .Y(n1810) );
  MUX2X1 U1308 ( .B(\mem<30><11> ), .A(\mem<31><11> ), .S(n1851), .Y(n1652) );
  MUX2X1 U1309 ( .B(\mem<28><11> ), .A(\mem<29><11> ), .S(n1851), .Y(n1651) );
  MUX2X1 U1310 ( .B(\mem<26><11> ), .A(\mem<27><11> ), .S(n1851), .Y(n1655) );
  MUX2X1 U1311 ( .B(\mem<24><11> ), .A(\mem<25><11> ), .S(n1851), .Y(n1654) );
  MUX2X1 U1312 ( .B(n1653), .A(n1650), .S(n1819), .Y(n1664) );
  MUX2X1 U1313 ( .B(\mem<22><11> ), .A(\mem<23><11> ), .S(n1851), .Y(n1658) );
  MUX2X1 U1314 ( .B(\mem<20><11> ), .A(\mem<21><11> ), .S(n1851), .Y(n1657) );
  MUX2X1 U1315 ( .B(\mem<18><11> ), .A(\mem<19><11> ), .S(n1851), .Y(n1661) );
  MUX2X1 U1316 ( .B(\mem<16><11> ), .A(\mem<17><11> ), .S(n1851), .Y(n1660) );
  MUX2X1 U1317 ( .B(n1659), .A(n1656), .S(n1819), .Y(n1663) );
  MUX2X1 U1318 ( .B(\mem<14><11> ), .A(\mem<15><11> ), .S(n1852), .Y(n1667) );
  MUX2X1 U1319 ( .B(\mem<12><11> ), .A(\mem<13><11> ), .S(n1852), .Y(n1666) );
  MUX2X1 U1320 ( .B(\mem<10><11> ), .A(\mem<11><11> ), .S(n1852), .Y(n1670) );
  MUX2X1 U1321 ( .B(\mem<8><11> ), .A(\mem<9><11> ), .S(n1852), .Y(n1669) );
  MUX2X1 U1322 ( .B(n1668), .A(n1665), .S(n1819), .Y(n1679) );
  MUX2X1 U1323 ( .B(\mem<6><11> ), .A(\mem<7><11> ), .S(n1852), .Y(n1673) );
  MUX2X1 U1324 ( .B(\mem<4><11> ), .A(\mem<5><11> ), .S(n1852), .Y(n1672) );
  MUX2X1 U1325 ( .B(\mem<2><11> ), .A(\mem<3><11> ), .S(n1852), .Y(n1676) );
  MUX2X1 U1326 ( .B(\mem<0><11> ), .A(\mem<1><11> ), .S(n1852), .Y(n1675) );
  MUX2X1 U1327 ( .B(n1674), .A(n1671), .S(n1819), .Y(n1678) );
  MUX2X1 U1328 ( .B(n1677), .A(n1662), .S(n1816), .Y(n1811) );
  MUX2X1 U1329 ( .B(\mem<30><12> ), .A(\mem<31><12> ), .S(n1852), .Y(n1682) );
  MUX2X1 U1330 ( .B(\mem<28><12> ), .A(\mem<29><12> ), .S(n1852), .Y(n1681) );
  MUX2X1 U1331 ( .B(\mem<26><12> ), .A(\mem<27><12> ), .S(n1852), .Y(n1685) );
  MUX2X1 U1332 ( .B(\mem<24><12> ), .A(\mem<25><12> ), .S(n1852), .Y(n1684) );
  MUX2X1 U1333 ( .B(n1683), .A(n1680), .S(n1822), .Y(n1694) );
  MUX2X1 U1334 ( .B(\mem<22><12> ), .A(\mem<23><12> ), .S(n1842), .Y(n1688) );
  MUX2X1 U1335 ( .B(\mem<20><12> ), .A(\mem<21><12> ), .S(n1850), .Y(n1687) );
  MUX2X1 U1336 ( .B(\mem<18><12> ), .A(\mem<19><12> ), .S(n1856), .Y(n1691) );
  MUX2X1 U1337 ( .B(\mem<16><12> ), .A(\mem<17><12> ), .S(n1856), .Y(n1690) );
  MUX2X1 U1338 ( .B(n1689), .A(n1686), .S(n1822), .Y(n1693) );
  MUX2X1 U1339 ( .B(\mem<14><12> ), .A(\mem<15><12> ), .S(n1845), .Y(n1697) );
  MUX2X1 U1340 ( .B(\mem<12><12> ), .A(\mem<13><12> ), .S(n1844), .Y(n1696) );
  MUX2X1 U1341 ( .B(\mem<10><12> ), .A(\mem<11><12> ), .S(n1851), .Y(n1700) );
  MUX2X1 U1342 ( .B(\mem<8><12> ), .A(\mem<9><12> ), .S(n1851), .Y(n1699) );
  MUX2X1 U1343 ( .B(n1698), .A(n1695), .S(n1822), .Y(n1709) );
  MUX2X1 U1344 ( .B(\mem<6><12> ), .A(\mem<7><12> ), .S(n1841), .Y(n1703) );
  MUX2X1 U1345 ( .B(\mem<4><12> ), .A(\mem<5><12> ), .S(n1843), .Y(n1702) );
  MUX2X1 U1346 ( .B(\mem<2><12> ), .A(\mem<3><12> ), .S(n1854), .Y(n1706) );
  MUX2X1 U1347 ( .B(\mem<0><12> ), .A(\mem<1><12> ), .S(n1849), .Y(n1705) );
  MUX2X1 U1348 ( .B(n1704), .A(n1701), .S(n1822), .Y(n1708) );
  MUX2X1 U1349 ( .B(n1707), .A(n1692), .S(n1816), .Y(n1812) );
  MUX2X1 U1350 ( .B(\mem<30><13> ), .A(\mem<31><13> ), .S(n1848), .Y(n1712) );
  MUX2X1 U1351 ( .B(\mem<28><13> ), .A(\mem<29><13> ), .S(n1843), .Y(n1711) );
  MUX2X1 U1352 ( .B(\mem<26><13> ), .A(\mem<27><13> ), .S(n1851), .Y(n1715) );
  MUX2X1 U1353 ( .B(\mem<24><13> ), .A(\mem<25><13> ), .S(n1844), .Y(n1714) );
  MUX2X1 U1354 ( .B(n1713), .A(n1710), .S(n1822), .Y(n1724) );
  MUX2X1 U1355 ( .B(\mem<22><13> ), .A(\mem<23><13> ), .S(n1849), .Y(n1718) );
  MUX2X1 U1356 ( .B(\mem<20><13> ), .A(\mem<21><13> ), .S(n1849), .Y(n1717) );
  MUX2X1 U1357 ( .B(\mem<18><13> ), .A(\mem<19><13> ), .S(n1851), .Y(n1721) );
  MUX2X1 U1358 ( .B(\mem<16><13> ), .A(\mem<17><13> ), .S(n1841), .Y(n1720) );
  MUX2X1 U1359 ( .B(n1719), .A(n1716), .S(n1822), .Y(n1723) );
  MUX2X1 U1360 ( .B(\mem<14><13> ), .A(\mem<15><13> ), .S(n1842), .Y(n1727) );
  MUX2X1 U1361 ( .B(\mem<12><13> ), .A(\mem<13><13> ), .S(n1851), .Y(n1726) );
  MUX2X1 U1362 ( .B(\mem<10><13> ), .A(\mem<11><13> ), .S(n1842), .Y(n1730) );
  MUX2X1 U1363 ( .B(\mem<8><13> ), .A(\mem<9><13> ), .S(n1846), .Y(n1729) );
  MUX2X1 U1364 ( .B(n1728), .A(n1725), .S(n1822), .Y(n1739) );
  MUX2X1 U1365 ( .B(\mem<6><13> ), .A(\mem<7><13> ), .S(n1853), .Y(n1733) );
  MUX2X1 U1366 ( .B(\mem<4><13> ), .A(\mem<5><13> ), .S(n1853), .Y(n1732) );
  MUX2X1 U1367 ( .B(\mem<2><13> ), .A(\mem<3><13> ), .S(n1853), .Y(n1736) );
  MUX2X1 U1368 ( .B(\mem<0><13> ), .A(\mem<1><13> ), .S(n1853), .Y(n1735) );
  MUX2X1 U1369 ( .B(n1734), .A(n1731), .S(n1822), .Y(n1738) );
  MUX2X1 U1370 ( .B(n1737), .A(n1722), .S(n1816), .Y(n1813) );
  MUX2X1 U1371 ( .B(\mem<30><14> ), .A(\mem<31><14> ), .S(n1853), .Y(n1742) );
  MUX2X1 U1372 ( .B(\mem<28><14> ), .A(\mem<29><14> ), .S(n1853), .Y(n1741) );
  MUX2X1 U1373 ( .B(\mem<26><14> ), .A(\mem<27><14> ), .S(n1853), .Y(n1745) );
  MUX2X1 U1374 ( .B(\mem<24><14> ), .A(\mem<25><14> ), .S(n1853), .Y(n1744) );
  MUX2X1 U1375 ( .B(n1743), .A(n1740), .S(n1822), .Y(n1754) );
  MUX2X1 U1376 ( .B(\mem<22><14> ), .A(\mem<23><14> ), .S(n1853), .Y(n1748) );
  MUX2X1 U1377 ( .B(\mem<20><14> ), .A(\mem<21><14> ), .S(n1853), .Y(n1747) );
  MUX2X1 U1378 ( .B(\mem<18><14> ), .A(\mem<19><14> ), .S(n1853), .Y(n1751) );
  MUX2X1 U1379 ( .B(\mem<16><14> ), .A(\mem<17><14> ), .S(n1853), .Y(n1750) );
  MUX2X1 U1380 ( .B(n1749), .A(n1746), .S(n1822), .Y(n1753) );
  MUX2X1 U1381 ( .B(\mem<14><14> ), .A(\mem<15><14> ), .S(n1854), .Y(n1757) );
  MUX2X1 U1382 ( .B(\mem<12><14> ), .A(\mem<13><14> ), .S(n1854), .Y(n1756) );
  MUX2X1 U1383 ( .B(\mem<10><14> ), .A(\mem<11><14> ), .S(n1854), .Y(n1760) );
  MUX2X1 U1384 ( .B(\mem<8><14> ), .A(\mem<9><14> ), .S(n1854), .Y(n1759) );
  MUX2X1 U1385 ( .B(n1758), .A(n1755), .S(n1822), .Y(n1769) );
  MUX2X1 U1386 ( .B(\mem<6><14> ), .A(\mem<7><14> ), .S(n1854), .Y(n1763) );
  MUX2X1 U1387 ( .B(\mem<4><14> ), .A(\mem<5><14> ), .S(n1854), .Y(n1762) );
  MUX2X1 U1388 ( .B(\mem<2><14> ), .A(\mem<3><14> ), .S(n1854), .Y(n1766) );
  MUX2X1 U1389 ( .B(\mem<0><14> ), .A(\mem<1><14> ), .S(n1854), .Y(n1765) );
  MUX2X1 U1390 ( .B(n1764), .A(n1761), .S(n1822), .Y(n1768) );
  MUX2X1 U1391 ( .B(n1767), .A(n1752), .S(n1816), .Y(n1814) );
  MUX2X1 U1392 ( .B(\mem<30><15> ), .A(\mem<31><15> ), .S(n1854), .Y(n1772) );
  MUX2X1 U1393 ( .B(\mem<28><15> ), .A(\mem<29><15> ), .S(n1854), .Y(n1771) );
  MUX2X1 U1394 ( .B(\mem<26><15> ), .A(\mem<27><15> ), .S(n1854), .Y(n1775) );
  MUX2X1 U1395 ( .B(\mem<24><15> ), .A(\mem<25><15> ), .S(n1854), .Y(n1774) );
  MUX2X1 U1396 ( .B(n1773), .A(n1770), .S(n1819), .Y(n1784) );
  MUX2X1 U1397 ( .B(\mem<22><15> ), .A(\mem<23><15> ), .S(n1842), .Y(n1778) );
  MUX2X1 U1398 ( .B(\mem<20><15> ), .A(\mem<21><15> ), .S(n1851), .Y(n1777) );
  MUX2X1 U1399 ( .B(\mem<18><15> ), .A(\mem<19><15> ), .S(n1847), .Y(n1781) );
  MUX2X1 U1400 ( .B(\mem<16><15> ), .A(\mem<17><15> ), .S(n1845), .Y(n1780) );
  MUX2X1 U1401 ( .B(n1779), .A(n1776), .S(n1821), .Y(n1783) );
  MUX2X1 U1402 ( .B(\mem<14><15> ), .A(\mem<15><15> ), .S(n1846), .Y(n1787) );
  MUX2X1 U1403 ( .B(\mem<12><15> ), .A(\mem<13><15> ), .S(n1847), .Y(n1786) );
  MUX2X1 U1404 ( .B(\mem<10><15> ), .A(\mem<11><15> ), .S(n1856), .Y(n1790) );
  MUX2X1 U1405 ( .B(\mem<8><15> ), .A(\mem<9><15> ), .S(n1856), .Y(n1789) );
  MUX2X1 U1406 ( .B(n1788), .A(n1785), .S(n1822), .Y(n1799) );
  MUX2X1 U1407 ( .B(\mem<6><15> ), .A(\mem<7><15> ), .S(n1843), .Y(n1793) );
  MUX2X1 U1408 ( .B(\mem<4><15> ), .A(\mem<5><15> ), .S(n1843), .Y(n1792) );
  MUX2X1 U1409 ( .B(\mem<2><15> ), .A(\mem<3><15> ), .S(n1856), .Y(n1796) );
  MUX2X1 U1410 ( .B(\mem<0><15> ), .A(\mem<1><15> ), .S(n1845), .Y(n1795) );
  MUX2X1 U1411 ( .B(n1794), .A(n1791), .S(n1820), .Y(n1798) );
  MUX2X1 U1412 ( .B(n1797), .A(n1782), .S(n1816), .Y(n1815) );
  INVX8 U1413 ( .A(n1840), .Y(n1841) );
  INVX8 U1414 ( .A(n1840), .Y(n1842) );
  INVX8 U1415 ( .A(n1840), .Y(n1843) );
  INVX8 U1416 ( .A(n1840), .Y(n1844) );
  INVX8 U1417 ( .A(n1840), .Y(n1850) );
  INVX8 U1418 ( .A(n1938), .Y(n1856) );
  INVX1 U1419 ( .A(N12), .Y(n1942) );
  INVX1 U1420 ( .A(N11), .Y(n1940) );
  INVX1 U1421 ( .A(N10), .Y(n1938) );
  INVX8 U1422 ( .A(n1904), .Y(n1901) );
  INVX8 U1423 ( .A(n1904), .Y(n1902) );
  INVX8 U1424 ( .A(n1904), .Y(n1903) );
  INVX8 U1425 ( .A(n4), .Y(n1905) );
  INVX8 U1426 ( .A(n4), .Y(n1906) );
  INVX8 U1427 ( .A(n6), .Y(n1907) );
  INVX8 U1428 ( .A(n6), .Y(n1908) );
  INVX8 U1429 ( .A(n7), .Y(n1909) );
  INVX8 U1430 ( .A(n7), .Y(n1910) );
  INVX8 U1431 ( .A(n8), .Y(n1911) );
  INVX8 U1432 ( .A(n8), .Y(n1912) );
  INVX8 U1433 ( .A(n9), .Y(n1913) );
  INVX8 U1434 ( .A(n9), .Y(n1914) );
  INVX8 U1435 ( .A(n10), .Y(n1915) );
  INVX8 U1436 ( .A(n10), .Y(n1916) );
  INVX8 U1437 ( .A(n11), .Y(n1917) );
  INVX8 U1438 ( .A(n11), .Y(n1918) );
  INVX8 U1439 ( .A(n12), .Y(n1919) );
  INVX8 U1440 ( .A(n12), .Y(n1920) );
  INVX8 U1441 ( .A(n13), .Y(n1921) );
  INVX8 U1442 ( .A(n13), .Y(n1922) );
  INVX8 U1443 ( .A(n14), .Y(n1923) );
  INVX8 U1444 ( .A(n14), .Y(n1924) );
  INVX8 U1445 ( .A(n15), .Y(n1925) );
  INVX8 U1446 ( .A(n15), .Y(n1926) );
  INVX8 U1447 ( .A(n16), .Y(n1927) );
  INVX8 U1448 ( .A(n16), .Y(n1928) );
  INVX8 U1449 ( .A(n17), .Y(n1929) );
  INVX8 U1450 ( .A(n17), .Y(n1930) );
  INVX8 U1451 ( .A(n18), .Y(n1931) );
  INVX8 U1452 ( .A(n18), .Y(n1932) );
  INVX8 U1453 ( .A(n19), .Y(n1933) );
  INVX8 U1454 ( .A(n19), .Y(n1934) );
  INVX8 U1455 ( .A(n20), .Y(n1935) );
  INVX8 U1456 ( .A(n20), .Y(n1936) );
  AND2X2 U1457 ( .A(N32), .B(n2), .Y(\data_out<0> ) );
  AND2X2 U1458 ( .A(N31), .B(n2), .Y(\data_out<1> ) );
  AND2X2 U1459 ( .A(N30), .B(n2), .Y(\data_out<2> ) );
  AND2X2 U1460 ( .A(N29), .B(n2), .Y(\data_out<3> ) );
  AND2X2 U1461 ( .A(N28), .B(n2), .Y(\data_out<4> ) );
  AND2X2 U1462 ( .A(N27), .B(n2), .Y(\data_out<5> ) );
  AND2X2 U1463 ( .A(N26), .B(n2), .Y(\data_out<6> ) );
  AND2X2 U1464 ( .A(N25), .B(n2), .Y(\data_out<7> ) );
  AND2X2 U1465 ( .A(N24), .B(n2), .Y(\data_out<8> ) );
  AND2X2 U1466 ( .A(n2), .B(N23), .Y(\data_out<9> ) );
  AND2X2 U1467 ( .A(N22), .B(n2), .Y(\data_out<10> ) );
  AND2X2 U1468 ( .A(N21), .B(n2), .Y(\data_out<11> ) );
  AND2X2 U1469 ( .A(N20), .B(n2), .Y(\data_out<12> ) );
  AND2X2 U1470 ( .A(N19), .B(n2), .Y(\data_out<13> ) );
  AND2X2 U1471 ( .A(n2), .B(N18), .Y(\data_out<14> ) );
  AND2X2 U1472 ( .A(N17), .B(n2), .Y(\data_out<15> ) );
  NAND2X1 U1473 ( .A(\mem<31><0> ), .B(n1244), .Y(n1945) );
  OAI21X1 U1474 ( .A(n1243), .B(n1905), .C(n1945), .Y(n2663) );
  NAND2X1 U1475 ( .A(\mem<31><1> ), .B(n1244), .Y(n1946) );
  OAI21X1 U1476 ( .A(n1908), .B(n1243), .C(n1946), .Y(n2662) );
  NAND2X1 U1477 ( .A(\mem<31><2> ), .B(n1244), .Y(n1947) );
  OAI21X1 U1478 ( .A(n1910), .B(n1243), .C(n1947), .Y(n2661) );
  NAND2X1 U1479 ( .A(\mem<31><3> ), .B(n1244), .Y(n1948) );
  OAI21X1 U1480 ( .A(n1912), .B(n1243), .C(n1948), .Y(n2660) );
  NAND2X1 U1481 ( .A(\mem<31><4> ), .B(n1244), .Y(n1949) );
  OAI21X1 U1482 ( .A(n1914), .B(n1243), .C(n1949), .Y(n2659) );
  NAND2X1 U1483 ( .A(\mem<31><5> ), .B(n1244), .Y(n1950) );
  OAI21X1 U1484 ( .A(n1916), .B(n1243), .C(n1950), .Y(n2658) );
  NAND2X1 U1485 ( .A(\mem<31><6> ), .B(n1244), .Y(n1951) );
  OAI21X1 U1486 ( .A(n1918), .B(n1243), .C(n1951), .Y(n2657) );
  NAND2X1 U1487 ( .A(\mem<31><7> ), .B(n1244), .Y(n1952) );
  OAI21X1 U1488 ( .A(n1920), .B(n1243), .C(n1952), .Y(n2656) );
  NAND2X1 U1489 ( .A(\mem<31><8> ), .B(n1244), .Y(n1953) );
  OAI21X1 U1490 ( .A(n1922), .B(n1243), .C(n1953), .Y(n2655) );
  NAND2X1 U1491 ( .A(\mem<31><9> ), .B(n1244), .Y(n1954) );
  OAI21X1 U1492 ( .A(n1924), .B(n1243), .C(n1954), .Y(n2654) );
  NAND2X1 U1493 ( .A(\mem<31><10> ), .B(n1244), .Y(n1955) );
  OAI21X1 U1494 ( .A(n1926), .B(n1243), .C(n1955), .Y(n2653) );
  NAND2X1 U1495 ( .A(\mem<31><11> ), .B(n1244), .Y(n1956) );
  OAI21X1 U1496 ( .A(n1928), .B(n1243), .C(n1956), .Y(n2652) );
  NAND2X1 U1497 ( .A(\mem<31><12> ), .B(n1244), .Y(n1957) );
  OAI21X1 U1498 ( .A(n1930), .B(n1243), .C(n1957), .Y(n2651) );
  NAND2X1 U1499 ( .A(\mem<31><13> ), .B(n1244), .Y(n1958) );
  OAI21X1 U1500 ( .A(n1932), .B(n1243), .C(n1958), .Y(n2650) );
  NAND2X1 U1501 ( .A(\mem<31><14> ), .B(n1244), .Y(n1959) );
  OAI21X1 U1502 ( .A(n1934), .B(n1243), .C(n1959), .Y(n2649) );
  NAND2X1 U1503 ( .A(\mem<31><15> ), .B(n1244), .Y(n1960) );
  OAI21X1 U1504 ( .A(n1936), .B(n1243), .C(n1960), .Y(n2648) );
  NAND2X1 U1505 ( .A(\mem<30><0> ), .B(n1247), .Y(n1961) );
  OAI21X1 U1506 ( .A(n1246), .B(n1905), .C(n1961), .Y(n2647) );
  NAND2X1 U1507 ( .A(\mem<30><1> ), .B(n1247), .Y(n1962) );
  OAI21X1 U1508 ( .A(n1246), .B(n1908), .C(n1962), .Y(n2646) );
  NAND2X1 U1509 ( .A(\mem<30><2> ), .B(n1247), .Y(n1963) );
  OAI21X1 U1510 ( .A(n1246), .B(n1910), .C(n1963), .Y(n2645) );
  NAND2X1 U1511 ( .A(\mem<30><3> ), .B(n1247), .Y(n1964) );
  OAI21X1 U1512 ( .A(n1246), .B(n1912), .C(n1964), .Y(n2644) );
  NAND2X1 U1513 ( .A(\mem<30><4> ), .B(n1247), .Y(n1965) );
  OAI21X1 U1514 ( .A(n1246), .B(n1914), .C(n1965), .Y(n2643) );
  NAND2X1 U1515 ( .A(\mem<30><5> ), .B(n1247), .Y(n1966) );
  OAI21X1 U1516 ( .A(n1246), .B(n1916), .C(n1966), .Y(n2642) );
  NAND2X1 U1517 ( .A(\mem<30><6> ), .B(n1247), .Y(n1967) );
  OAI21X1 U1518 ( .A(n1246), .B(n1918), .C(n1967), .Y(n2641) );
  NAND2X1 U1519 ( .A(\mem<30><7> ), .B(n1247), .Y(n1968) );
  OAI21X1 U1520 ( .A(n1246), .B(n1920), .C(n1968), .Y(n2640) );
  NAND2X1 U1521 ( .A(\mem<30><8> ), .B(n1247), .Y(n1969) );
  OAI21X1 U1522 ( .A(n1246), .B(n1921), .C(n1969), .Y(n2639) );
  NAND2X1 U1523 ( .A(\mem<30><9> ), .B(n1247), .Y(n1970) );
  OAI21X1 U1524 ( .A(n1246), .B(n1923), .C(n1970), .Y(n2638) );
  NAND2X1 U1525 ( .A(\mem<30><10> ), .B(n1247), .Y(n1971) );
  OAI21X1 U1526 ( .A(n1246), .B(n1925), .C(n1971), .Y(n2637) );
  NAND2X1 U1527 ( .A(\mem<30><11> ), .B(n1247), .Y(n1972) );
  OAI21X1 U1528 ( .A(n1246), .B(n1927), .C(n1972), .Y(n2636) );
  NAND2X1 U1529 ( .A(\mem<30><12> ), .B(n1247), .Y(n1973) );
  OAI21X1 U1530 ( .A(n1246), .B(n1929), .C(n1973), .Y(n2635) );
  NAND2X1 U1531 ( .A(\mem<30><13> ), .B(n1247), .Y(n1974) );
  OAI21X1 U1532 ( .A(n1246), .B(n1931), .C(n1974), .Y(n2634) );
  NAND2X1 U1533 ( .A(\mem<30><14> ), .B(n1247), .Y(n1975) );
  OAI21X1 U1534 ( .A(n1246), .B(n1933), .C(n1975), .Y(n2633) );
  NAND2X1 U1535 ( .A(\mem<30><15> ), .B(n1247), .Y(n1976) );
  OAI21X1 U1536 ( .A(n1246), .B(n1935), .C(n1976), .Y(n2632) );
  NAND3X1 U1537 ( .A(n1853), .B(n1941), .C(n1940), .Y(n1977) );
  NAND2X1 U1538 ( .A(\mem<29><0> ), .B(n1251), .Y(n1978) );
  OAI21X1 U1539 ( .A(n1249), .B(n1905), .C(n1978), .Y(n2631) );
  NAND2X1 U1540 ( .A(\mem<29><1> ), .B(n1251), .Y(n1979) );
  OAI21X1 U1541 ( .A(n1249), .B(n1907), .C(n1979), .Y(n2630) );
  NAND2X1 U1542 ( .A(\mem<29><2> ), .B(n1251), .Y(n1980) );
  OAI21X1 U1543 ( .A(n1249), .B(n1909), .C(n1980), .Y(n2629) );
  NAND2X1 U1544 ( .A(\mem<29><3> ), .B(n1251), .Y(n1981) );
  OAI21X1 U1545 ( .A(n1249), .B(n1911), .C(n1981), .Y(n2628) );
  NAND2X1 U1546 ( .A(\mem<29><4> ), .B(n1251), .Y(n1982) );
  OAI21X1 U1547 ( .A(n1249), .B(n1913), .C(n1982), .Y(n2627) );
  NAND2X1 U1548 ( .A(\mem<29><5> ), .B(n1251), .Y(n1983) );
  OAI21X1 U1549 ( .A(n1249), .B(n1915), .C(n1983), .Y(n2626) );
  NAND2X1 U1550 ( .A(\mem<29><6> ), .B(n1251), .Y(n1984) );
  OAI21X1 U1551 ( .A(n1249), .B(n1917), .C(n1984), .Y(n2625) );
  NAND2X1 U1552 ( .A(\mem<29><7> ), .B(n1251), .Y(n1985) );
  OAI21X1 U1553 ( .A(n1249), .B(n1919), .C(n1985), .Y(n2624) );
  NAND2X1 U1554 ( .A(\mem<29><8> ), .B(n1250), .Y(n1986) );
  OAI21X1 U1555 ( .A(n1249), .B(n1922), .C(n1986), .Y(n2623) );
  NAND2X1 U1556 ( .A(\mem<29><9> ), .B(n1250), .Y(n1987) );
  OAI21X1 U1557 ( .A(n1249), .B(n1924), .C(n1987), .Y(n2622) );
  NAND2X1 U1558 ( .A(\mem<29><10> ), .B(n1250), .Y(n1988) );
  OAI21X1 U1559 ( .A(n1249), .B(n1926), .C(n1988), .Y(n2621) );
  NAND2X1 U1560 ( .A(\mem<29><11> ), .B(n1250), .Y(n1989) );
  OAI21X1 U1561 ( .A(n1249), .B(n1928), .C(n1989), .Y(n2620) );
  NAND2X1 U1562 ( .A(\mem<29><12> ), .B(n1250), .Y(n1990) );
  OAI21X1 U1563 ( .A(n1249), .B(n1930), .C(n1990), .Y(n2619) );
  NAND2X1 U1564 ( .A(\mem<29><13> ), .B(n1250), .Y(n1991) );
  OAI21X1 U1565 ( .A(n1249), .B(n1932), .C(n1991), .Y(n2618) );
  NAND2X1 U1566 ( .A(\mem<29><14> ), .B(n1250), .Y(n1992) );
  OAI21X1 U1567 ( .A(n1249), .B(n1934), .C(n1992), .Y(n2617) );
  NAND2X1 U1568 ( .A(\mem<29><15> ), .B(n1250), .Y(n1993) );
  OAI21X1 U1569 ( .A(n1249), .B(n1936), .C(n1993), .Y(n2616) );
  NAND3X1 U1570 ( .A(n1941), .B(n1940), .C(n1938), .Y(n1994) );
  NAND2X1 U1571 ( .A(\mem<28><0> ), .B(n1255), .Y(n1995) );
  OAI21X1 U1572 ( .A(n1253), .B(n1905), .C(n1995), .Y(n2615) );
  NAND2X1 U1573 ( .A(\mem<28><1> ), .B(n1255), .Y(n1996) );
  OAI21X1 U1574 ( .A(n1253), .B(n1908), .C(n1996), .Y(n2614) );
  NAND2X1 U1575 ( .A(\mem<28><2> ), .B(n1255), .Y(n1997) );
  OAI21X1 U1576 ( .A(n1253), .B(n1910), .C(n1997), .Y(n2613) );
  NAND2X1 U1577 ( .A(\mem<28><3> ), .B(n1255), .Y(n1998) );
  OAI21X1 U1578 ( .A(n1253), .B(n1912), .C(n1998), .Y(n2612) );
  NAND2X1 U1579 ( .A(\mem<28><4> ), .B(n1255), .Y(n1999) );
  OAI21X1 U1580 ( .A(n1253), .B(n1914), .C(n1999), .Y(n2611) );
  NAND2X1 U1581 ( .A(\mem<28><5> ), .B(n1255), .Y(n2000) );
  OAI21X1 U1582 ( .A(n1253), .B(n1916), .C(n2000), .Y(n2610) );
  NAND2X1 U1583 ( .A(\mem<28><6> ), .B(n1255), .Y(n2001) );
  OAI21X1 U1584 ( .A(n1253), .B(n1918), .C(n2001), .Y(n2609) );
  NAND2X1 U1585 ( .A(\mem<28><7> ), .B(n1255), .Y(n2002) );
  OAI21X1 U1586 ( .A(n1253), .B(n1920), .C(n2002), .Y(n2608) );
  NAND2X1 U1587 ( .A(\mem<28><8> ), .B(n1254), .Y(n2003) );
  OAI21X1 U1588 ( .A(n1253), .B(n1921), .C(n2003), .Y(n2607) );
  NAND2X1 U1589 ( .A(\mem<28><9> ), .B(n1254), .Y(n2004) );
  OAI21X1 U1590 ( .A(n1253), .B(n1923), .C(n2004), .Y(n2606) );
  NAND2X1 U1591 ( .A(\mem<28><10> ), .B(n1254), .Y(n2005) );
  OAI21X1 U1592 ( .A(n1253), .B(n1925), .C(n2005), .Y(n2605) );
  NAND2X1 U1593 ( .A(\mem<28><11> ), .B(n1254), .Y(n2006) );
  OAI21X1 U1594 ( .A(n1253), .B(n1927), .C(n2006), .Y(n2604) );
  NAND2X1 U1595 ( .A(\mem<28><12> ), .B(n1254), .Y(n2007) );
  OAI21X1 U1596 ( .A(n1253), .B(n1929), .C(n2007), .Y(n2603) );
  NAND2X1 U1597 ( .A(\mem<28><13> ), .B(n1254), .Y(n2008) );
  OAI21X1 U1598 ( .A(n1253), .B(n1931), .C(n2008), .Y(n2602) );
  NAND2X1 U1599 ( .A(\mem<28><14> ), .B(n1254), .Y(n2009) );
  OAI21X1 U1600 ( .A(n1253), .B(n1933), .C(n2009), .Y(n2601) );
  NAND2X1 U1601 ( .A(\mem<28><15> ), .B(n1254), .Y(n2010) );
  OAI21X1 U1602 ( .A(n1253), .B(n1935), .C(n2010), .Y(n2600) );
  NAND3X1 U1603 ( .A(n1853), .B(n1939), .C(n1942), .Y(n2011) );
  NAND2X1 U1604 ( .A(\mem<27><0> ), .B(n1259), .Y(n2012) );
  OAI21X1 U1605 ( .A(n1257), .B(n1905), .C(n2012), .Y(n2599) );
  NAND2X1 U1606 ( .A(\mem<27><1> ), .B(n1259), .Y(n2013) );
  OAI21X1 U1607 ( .A(n1257), .B(n1907), .C(n2013), .Y(n2598) );
  NAND2X1 U1608 ( .A(\mem<27><2> ), .B(n1259), .Y(n2014) );
  OAI21X1 U1609 ( .A(n1257), .B(n1909), .C(n2014), .Y(n2597) );
  NAND2X1 U1610 ( .A(\mem<27><3> ), .B(n1259), .Y(n2015) );
  OAI21X1 U1611 ( .A(n1257), .B(n1911), .C(n2015), .Y(n2596) );
  NAND2X1 U1612 ( .A(\mem<27><4> ), .B(n1259), .Y(n2016) );
  OAI21X1 U1613 ( .A(n1257), .B(n1913), .C(n2016), .Y(n2595) );
  NAND2X1 U1614 ( .A(\mem<27><5> ), .B(n1259), .Y(n2017) );
  OAI21X1 U1615 ( .A(n1257), .B(n1915), .C(n2017), .Y(n2594) );
  NAND2X1 U1616 ( .A(\mem<27><6> ), .B(n1259), .Y(n2018) );
  OAI21X1 U1617 ( .A(n1257), .B(n1917), .C(n2018), .Y(n2593) );
  NAND2X1 U1618 ( .A(\mem<27><7> ), .B(n1259), .Y(n2019) );
  OAI21X1 U1619 ( .A(n1257), .B(n1919), .C(n2019), .Y(n2592) );
  NAND2X1 U1620 ( .A(\mem<27><8> ), .B(n1258), .Y(n2020) );
  OAI21X1 U1621 ( .A(n1257), .B(n1922), .C(n2020), .Y(n2591) );
  NAND2X1 U1622 ( .A(\mem<27><9> ), .B(n1258), .Y(n2021) );
  OAI21X1 U1623 ( .A(n1257), .B(n1924), .C(n2021), .Y(n2590) );
  NAND2X1 U1624 ( .A(\mem<27><10> ), .B(n1258), .Y(n2022) );
  OAI21X1 U1625 ( .A(n1257), .B(n1926), .C(n2022), .Y(n2589) );
  NAND2X1 U1626 ( .A(\mem<27><11> ), .B(n1258), .Y(n2023) );
  OAI21X1 U1627 ( .A(n1257), .B(n1928), .C(n2023), .Y(n2588) );
  NAND2X1 U1628 ( .A(\mem<27><12> ), .B(n1258), .Y(n2024) );
  OAI21X1 U1629 ( .A(n1257), .B(n1930), .C(n2024), .Y(n2587) );
  NAND2X1 U1630 ( .A(\mem<27><13> ), .B(n1258), .Y(n2025) );
  OAI21X1 U1631 ( .A(n1257), .B(n1932), .C(n2025), .Y(n2586) );
  NAND2X1 U1632 ( .A(\mem<27><14> ), .B(n1258), .Y(n2026) );
  OAI21X1 U1633 ( .A(n1257), .B(n1934), .C(n2026), .Y(n2585) );
  NAND2X1 U1634 ( .A(\mem<27><15> ), .B(n1258), .Y(n2027) );
  OAI21X1 U1635 ( .A(n1257), .B(n1936), .C(n2027), .Y(n2584) );
  NAND3X1 U1636 ( .A(n1942), .B(n1939), .C(n1938), .Y(n2028) );
  NAND2X1 U1637 ( .A(\mem<26><0> ), .B(n1263), .Y(n2029) );
  OAI21X1 U1638 ( .A(n1261), .B(n1905), .C(n2029), .Y(n2583) );
  NAND2X1 U1639 ( .A(\mem<26><1> ), .B(n1263), .Y(n2030) );
  OAI21X1 U1640 ( .A(n1261), .B(n1908), .C(n2030), .Y(n2582) );
  NAND2X1 U1641 ( .A(\mem<26><2> ), .B(n1263), .Y(n2031) );
  OAI21X1 U1642 ( .A(n1261), .B(n1910), .C(n2031), .Y(n2581) );
  NAND2X1 U1643 ( .A(\mem<26><3> ), .B(n1263), .Y(n2032) );
  OAI21X1 U1644 ( .A(n1261), .B(n1912), .C(n2032), .Y(n2580) );
  NAND2X1 U1645 ( .A(\mem<26><4> ), .B(n1263), .Y(n2033) );
  OAI21X1 U1646 ( .A(n1261), .B(n1914), .C(n2033), .Y(n2579) );
  NAND2X1 U1647 ( .A(\mem<26><5> ), .B(n1263), .Y(n2034) );
  OAI21X1 U1648 ( .A(n1261), .B(n1916), .C(n2034), .Y(n2578) );
  NAND2X1 U1649 ( .A(\mem<26><6> ), .B(n1263), .Y(n2035) );
  OAI21X1 U1650 ( .A(n1261), .B(n1918), .C(n2035), .Y(n2577) );
  NAND2X1 U1651 ( .A(\mem<26><7> ), .B(n1263), .Y(n2036) );
  OAI21X1 U1652 ( .A(n1261), .B(n1920), .C(n2036), .Y(n2576) );
  NAND2X1 U1653 ( .A(\mem<26><8> ), .B(n1262), .Y(n2037) );
  OAI21X1 U1654 ( .A(n1261), .B(n1921), .C(n2037), .Y(n2575) );
  NAND2X1 U1655 ( .A(\mem<26><9> ), .B(n1262), .Y(n2038) );
  OAI21X1 U1656 ( .A(n1261), .B(n1923), .C(n2038), .Y(n2574) );
  NAND2X1 U1657 ( .A(\mem<26><10> ), .B(n1262), .Y(n2039) );
  OAI21X1 U1658 ( .A(n1261), .B(n1925), .C(n2039), .Y(n2573) );
  NAND2X1 U1659 ( .A(\mem<26><11> ), .B(n1262), .Y(n2040) );
  OAI21X1 U1660 ( .A(n1261), .B(n1927), .C(n2040), .Y(n2572) );
  NAND2X1 U1661 ( .A(\mem<26><12> ), .B(n1262), .Y(n2041) );
  OAI21X1 U1662 ( .A(n1261), .B(n1929), .C(n2041), .Y(n2571) );
  NAND2X1 U1663 ( .A(\mem<26><13> ), .B(n1262), .Y(n2042) );
  OAI21X1 U1664 ( .A(n1261), .B(n1931), .C(n2042), .Y(n2570) );
  NAND2X1 U1665 ( .A(\mem<26><14> ), .B(n1262), .Y(n2043) );
  OAI21X1 U1666 ( .A(n1261), .B(n1933), .C(n2043), .Y(n2569) );
  NAND2X1 U1667 ( .A(\mem<26><15> ), .B(n1262), .Y(n2044) );
  OAI21X1 U1668 ( .A(n1261), .B(n1935), .C(n2044), .Y(n2568) );
  NAND3X1 U1669 ( .A(n1854), .B(n1942), .C(n1940), .Y(n2045) );
  NAND2X1 U1670 ( .A(\mem<25><0> ), .B(n1267), .Y(n2046) );
  OAI21X1 U1671 ( .A(n1265), .B(n1905), .C(n2046), .Y(n2567) );
  NAND2X1 U1672 ( .A(\mem<25><1> ), .B(n1267), .Y(n2047) );
  OAI21X1 U1673 ( .A(n1265), .B(n1907), .C(n2047), .Y(n2566) );
  NAND2X1 U1674 ( .A(\mem<25><2> ), .B(n1267), .Y(n2048) );
  OAI21X1 U1675 ( .A(n1265), .B(n1909), .C(n2048), .Y(n2565) );
  NAND2X1 U1676 ( .A(\mem<25><3> ), .B(n1267), .Y(n2049) );
  OAI21X1 U1677 ( .A(n1265), .B(n1911), .C(n2049), .Y(n2564) );
  NAND2X1 U1678 ( .A(\mem<25><4> ), .B(n1267), .Y(n2050) );
  OAI21X1 U1679 ( .A(n1265), .B(n1913), .C(n2050), .Y(n2563) );
  NAND2X1 U1680 ( .A(\mem<25><5> ), .B(n1267), .Y(n2051) );
  OAI21X1 U1681 ( .A(n1265), .B(n1915), .C(n2051), .Y(n2562) );
  NAND2X1 U1682 ( .A(\mem<25><6> ), .B(n1267), .Y(n2052) );
  OAI21X1 U1683 ( .A(n1265), .B(n1917), .C(n2052), .Y(n2561) );
  NAND2X1 U1684 ( .A(\mem<25><7> ), .B(n1267), .Y(n2053) );
  OAI21X1 U1685 ( .A(n1265), .B(n1919), .C(n2053), .Y(n2560) );
  NAND2X1 U1686 ( .A(\mem<25><8> ), .B(n1266), .Y(n2054) );
  OAI21X1 U1687 ( .A(n1265), .B(n1922), .C(n2054), .Y(n2559) );
  NAND2X1 U1688 ( .A(\mem<25><9> ), .B(n1266), .Y(n2055) );
  OAI21X1 U1689 ( .A(n1265), .B(n1924), .C(n2055), .Y(n2558) );
  NAND2X1 U1690 ( .A(\mem<25><10> ), .B(n1266), .Y(n2056) );
  OAI21X1 U1691 ( .A(n1265), .B(n1926), .C(n2056), .Y(n2557) );
  NAND2X1 U1692 ( .A(\mem<25><11> ), .B(n1266), .Y(n2057) );
  OAI21X1 U1693 ( .A(n1265), .B(n1928), .C(n2057), .Y(n2556) );
  NAND2X1 U1694 ( .A(\mem<25><12> ), .B(n1266), .Y(n2058) );
  OAI21X1 U1695 ( .A(n1265), .B(n1930), .C(n2058), .Y(n2555) );
  NAND2X1 U1696 ( .A(\mem<25><13> ), .B(n1266), .Y(n2059) );
  OAI21X1 U1697 ( .A(n1265), .B(n1932), .C(n2059), .Y(n2554) );
  NAND2X1 U1698 ( .A(\mem<25><14> ), .B(n1266), .Y(n2060) );
  OAI21X1 U1699 ( .A(n1265), .B(n1934), .C(n2060), .Y(n2553) );
  NAND2X1 U1700 ( .A(\mem<25><15> ), .B(n1266), .Y(n2061) );
  OAI21X1 U1701 ( .A(n1265), .B(n1936), .C(n2061), .Y(n2552) );
  NOR3X1 U1702 ( .A(n1851), .B(n1939), .C(n1941), .Y(n2151) );
  NAND2X1 U1703 ( .A(\mem<24><0> ), .B(n1269), .Y(n2062) );
  OAI21X1 U1704 ( .A(n1857), .B(n1905), .C(n2062), .Y(n2551) );
  NAND2X1 U1705 ( .A(\mem<24><1> ), .B(n1269), .Y(n2063) );
  OAI21X1 U1706 ( .A(n1857), .B(n1907), .C(n2063), .Y(n2550) );
  NAND2X1 U1707 ( .A(\mem<24><2> ), .B(n1269), .Y(n2064) );
  OAI21X1 U1708 ( .A(n1857), .B(n1909), .C(n2064), .Y(n2549) );
  NAND2X1 U1709 ( .A(\mem<24><3> ), .B(n1269), .Y(n2065) );
  OAI21X1 U1710 ( .A(n1857), .B(n1911), .C(n2065), .Y(n2548) );
  NAND2X1 U1711 ( .A(\mem<24><4> ), .B(n1269), .Y(n2066) );
  OAI21X1 U1712 ( .A(n1857), .B(n1913), .C(n2066), .Y(n2547) );
  NAND2X1 U1713 ( .A(\mem<24><5> ), .B(n1269), .Y(n2067) );
  OAI21X1 U1714 ( .A(n1857), .B(n1915), .C(n2067), .Y(n2546) );
  NAND2X1 U1715 ( .A(\mem<24><6> ), .B(n1269), .Y(n2068) );
  OAI21X1 U1716 ( .A(n1857), .B(n1917), .C(n2068), .Y(n2545) );
  NAND2X1 U1717 ( .A(\mem<24><7> ), .B(n1269), .Y(n2069) );
  OAI21X1 U1718 ( .A(n1857), .B(n1919), .C(n2069), .Y(n2544) );
  NAND2X1 U1719 ( .A(\mem<24><8> ), .B(n1268), .Y(n2070) );
  OAI21X1 U1720 ( .A(n1857), .B(n1921), .C(n2070), .Y(n2543) );
  NAND2X1 U1721 ( .A(\mem<24><9> ), .B(n1268), .Y(n2071) );
  OAI21X1 U1722 ( .A(n1857), .B(n1923), .C(n2071), .Y(n2542) );
  NAND2X1 U1723 ( .A(\mem<24><10> ), .B(n1268), .Y(n2072) );
  OAI21X1 U1724 ( .A(n1857), .B(n1925), .C(n2072), .Y(n2541) );
  NAND2X1 U1725 ( .A(\mem<24><11> ), .B(n1268), .Y(n2073) );
  OAI21X1 U1726 ( .A(n1857), .B(n1927), .C(n2073), .Y(n2540) );
  NAND2X1 U1727 ( .A(\mem<24><12> ), .B(n1268), .Y(n2074) );
  OAI21X1 U1728 ( .A(n1857), .B(n1929), .C(n2074), .Y(n2539) );
  NAND2X1 U1729 ( .A(\mem<24><13> ), .B(n1268), .Y(n2075) );
  OAI21X1 U1730 ( .A(n1857), .B(n1931), .C(n2075), .Y(n2538) );
  NAND2X1 U1731 ( .A(\mem<24><14> ), .B(n1268), .Y(n2076) );
  OAI21X1 U1732 ( .A(n1857), .B(n1933), .C(n2076), .Y(n2537) );
  NAND2X1 U1733 ( .A(\mem<24><15> ), .B(n1268), .Y(n2077) );
  OAI21X1 U1734 ( .A(n1857), .B(n1935), .C(n2077), .Y(n2536) );
  NAND2X1 U1735 ( .A(\mem<23><0> ), .B(n1273), .Y(n2078) );
  OAI21X1 U1736 ( .A(n1271), .B(n1905), .C(n2078), .Y(n2535) );
  NAND2X1 U1737 ( .A(\mem<23><1> ), .B(n1273), .Y(n2079) );
  OAI21X1 U1738 ( .A(n1271), .B(n1908), .C(n2079), .Y(n2534) );
  NAND2X1 U1739 ( .A(\mem<23><2> ), .B(n1273), .Y(n2080) );
  OAI21X1 U1740 ( .A(n1271), .B(n1910), .C(n2080), .Y(n2533) );
  NAND2X1 U1741 ( .A(\mem<23><3> ), .B(n1273), .Y(n2081) );
  OAI21X1 U1742 ( .A(n1271), .B(n1912), .C(n2081), .Y(n2532) );
  NAND2X1 U1743 ( .A(\mem<23><4> ), .B(n1273), .Y(n2082) );
  OAI21X1 U1744 ( .A(n1271), .B(n1914), .C(n2082), .Y(n2531) );
  NAND2X1 U1745 ( .A(\mem<23><5> ), .B(n1273), .Y(n2083) );
  OAI21X1 U1746 ( .A(n1271), .B(n1916), .C(n2083), .Y(n2530) );
  NAND2X1 U1747 ( .A(\mem<23><6> ), .B(n1273), .Y(n2084) );
  OAI21X1 U1748 ( .A(n1271), .B(n1918), .C(n2084), .Y(n2529) );
  NAND2X1 U1749 ( .A(\mem<23><7> ), .B(n1273), .Y(n2085) );
  OAI21X1 U1750 ( .A(n1271), .B(n1920), .C(n2085), .Y(n2528) );
  NAND2X1 U1751 ( .A(\mem<23><8> ), .B(n1272), .Y(n2086) );
  OAI21X1 U1752 ( .A(n1271), .B(n1922), .C(n2086), .Y(n2527) );
  NAND2X1 U1753 ( .A(\mem<23><9> ), .B(n1272), .Y(n2087) );
  OAI21X1 U1754 ( .A(n1271), .B(n1924), .C(n2087), .Y(n2526) );
  NAND2X1 U1755 ( .A(\mem<23><10> ), .B(n1272), .Y(n2088) );
  OAI21X1 U1756 ( .A(n1271), .B(n1926), .C(n2088), .Y(n2525) );
  NAND2X1 U1757 ( .A(\mem<23><11> ), .B(n1272), .Y(n2089) );
  OAI21X1 U1758 ( .A(n1271), .B(n1928), .C(n2089), .Y(n2524) );
  NAND2X1 U1759 ( .A(\mem<23><12> ), .B(n1272), .Y(n2090) );
  OAI21X1 U1760 ( .A(n1271), .B(n1930), .C(n2090), .Y(n2523) );
  NAND2X1 U1761 ( .A(\mem<23><13> ), .B(n1272), .Y(n2091) );
  OAI21X1 U1762 ( .A(n1271), .B(n1932), .C(n2091), .Y(n2522) );
  NAND2X1 U1763 ( .A(\mem<23><14> ), .B(n1272), .Y(n2092) );
  OAI21X1 U1764 ( .A(n1271), .B(n1934), .C(n2092), .Y(n2521) );
  NAND2X1 U1765 ( .A(\mem<23><15> ), .B(n1272), .Y(n2093) );
  OAI21X1 U1766 ( .A(n1271), .B(n1936), .C(n2093), .Y(n2520) );
  NAND2X1 U1767 ( .A(\mem<22><0> ), .B(n1277), .Y(n2094) );
  OAI21X1 U1768 ( .A(n1275), .B(n1905), .C(n2094), .Y(n2519) );
  NAND2X1 U1769 ( .A(\mem<22><1> ), .B(n1277), .Y(n2095) );
  OAI21X1 U1770 ( .A(n1275), .B(n1908), .C(n2095), .Y(n2518) );
  NAND2X1 U1771 ( .A(\mem<22><2> ), .B(n1277), .Y(n2096) );
  OAI21X1 U1772 ( .A(n1275), .B(n1910), .C(n2096), .Y(n2517) );
  NAND2X1 U1773 ( .A(\mem<22><3> ), .B(n1277), .Y(n2097) );
  OAI21X1 U1774 ( .A(n1275), .B(n1912), .C(n2097), .Y(n2516) );
  NAND2X1 U1775 ( .A(\mem<22><4> ), .B(n1277), .Y(n2098) );
  OAI21X1 U1776 ( .A(n1275), .B(n1914), .C(n2098), .Y(n2515) );
  NAND2X1 U1777 ( .A(\mem<22><5> ), .B(n1277), .Y(n2099) );
  OAI21X1 U1778 ( .A(n1275), .B(n1916), .C(n2099), .Y(n2514) );
  NAND2X1 U1779 ( .A(\mem<22><6> ), .B(n1277), .Y(n2100) );
  OAI21X1 U1780 ( .A(n1275), .B(n1918), .C(n2100), .Y(n2513) );
  NAND2X1 U1781 ( .A(\mem<22><7> ), .B(n1277), .Y(n2101) );
  OAI21X1 U1782 ( .A(n1275), .B(n1920), .C(n2101), .Y(n2512) );
  NAND2X1 U1783 ( .A(\mem<22><8> ), .B(n1276), .Y(n2102) );
  OAI21X1 U1784 ( .A(n1275), .B(n1922), .C(n2102), .Y(n2511) );
  NAND2X1 U1785 ( .A(\mem<22><9> ), .B(n1276), .Y(n2103) );
  OAI21X1 U1786 ( .A(n1275), .B(n1924), .C(n2103), .Y(n2510) );
  NAND2X1 U1787 ( .A(\mem<22><10> ), .B(n1276), .Y(n2104) );
  OAI21X1 U1788 ( .A(n1275), .B(n1926), .C(n2104), .Y(n2509) );
  NAND2X1 U1789 ( .A(\mem<22><11> ), .B(n1276), .Y(n2105) );
  OAI21X1 U1790 ( .A(n1275), .B(n1928), .C(n2105), .Y(n2508) );
  NAND2X1 U1791 ( .A(\mem<22><12> ), .B(n1276), .Y(n2106) );
  OAI21X1 U1792 ( .A(n1275), .B(n1930), .C(n2106), .Y(n2507) );
  NAND2X1 U1793 ( .A(\mem<22><13> ), .B(n1276), .Y(n2107) );
  OAI21X1 U1794 ( .A(n1275), .B(n1932), .C(n2107), .Y(n2506) );
  NAND2X1 U1795 ( .A(\mem<22><14> ), .B(n1276), .Y(n2108) );
  OAI21X1 U1796 ( .A(n1275), .B(n1934), .C(n2108), .Y(n2505) );
  NAND2X1 U1797 ( .A(\mem<22><15> ), .B(n1276), .Y(n2109) );
  OAI21X1 U1798 ( .A(n1275), .B(n1936), .C(n2109), .Y(n2504) );
  NAND2X1 U1799 ( .A(\mem<21><0> ), .B(n1281), .Y(n2110) );
  OAI21X1 U1800 ( .A(n1279), .B(n1905), .C(n2110), .Y(n2503) );
  NAND2X1 U1801 ( .A(\mem<21><1> ), .B(n1281), .Y(n2111) );
  OAI21X1 U1802 ( .A(n1279), .B(n1908), .C(n2111), .Y(n2502) );
  NAND2X1 U1803 ( .A(\mem<21><2> ), .B(n1281), .Y(n2112) );
  OAI21X1 U1804 ( .A(n1279), .B(n1910), .C(n2112), .Y(n2501) );
  NAND2X1 U1805 ( .A(\mem<21><3> ), .B(n1281), .Y(n2113) );
  OAI21X1 U1806 ( .A(n1279), .B(n1912), .C(n2113), .Y(n2500) );
  NAND2X1 U1807 ( .A(\mem<21><4> ), .B(n1281), .Y(n2114) );
  OAI21X1 U1808 ( .A(n1279), .B(n1914), .C(n2114), .Y(n2499) );
  NAND2X1 U1809 ( .A(\mem<21><5> ), .B(n1281), .Y(n2115) );
  OAI21X1 U1810 ( .A(n1279), .B(n1916), .C(n2115), .Y(n2498) );
  NAND2X1 U1811 ( .A(\mem<21><6> ), .B(n1281), .Y(n2116) );
  OAI21X1 U1812 ( .A(n1279), .B(n1918), .C(n2116), .Y(n2497) );
  NAND2X1 U1813 ( .A(\mem<21><7> ), .B(n1281), .Y(n2117) );
  OAI21X1 U1814 ( .A(n1279), .B(n1920), .C(n2117), .Y(n2496) );
  NAND2X1 U1815 ( .A(\mem<21><8> ), .B(n1280), .Y(n2118) );
  OAI21X1 U1816 ( .A(n1279), .B(n1922), .C(n2118), .Y(n2495) );
  NAND2X1 U1817 ( .A(\mem<21><9> ), .B(n1280), .Y(n2119) );
  OAI21X1 U1818 ( .A(n1279), .B(n1924), .C(n2119), .Y(n2494) );
  NAND2X1 U1819 ( .A(\mem<21><10> ), .B(n1280), .Y(n2120) );
  OAI21X1 U1820 ( .A(n1279), .B(n1926), .C(n2120), .Y(n2493) );
  NAND2X1 U1821 ( .A(\mem<21><11> ), .B(n1280), .Y(n2121) );
  OAI21X1 U1822 ( .A(n1279), .B(n1928), .C(n2121), .Y(n2492) );
  NAND2X1 U1823 ( .A(\mem<21><12> ), .B(n1280), .Y(n2122) );
  OAI21X1 U1824 ( .A(n1279), .B(n1930), .C(n2122), .Y(n2491) );
  NAND2X1 U1825 ( .A(\mem<21><13> ), .B(n1280), .Y(n2123) );
  OAI21X1 U1826 ( .A(n1279), .B(n1932), .C(n2123), .Y(n2490) );
  NAND2X1 U1827 ( .A(\mem<21><14> ), .B(n1280), .Y(n2124) );
  OAI21X1 U1828 ( .A(n1279), .B(n1934), .C(n2124), .Y(n2489) );
  NAND2X1 U1829 ( .A(\mem<21><15> ), .B(n1280), .Y(n2125) );
  OAI21X1 U1830 ( .A(n1279), .B(n1936), .C(n2125), .Y(n2488) );
  NAND2X1 U1831 ( .A(\mem<20><0> ), .B(n1285), .Y(n2126) );
  OAI21X1 U1832 ( .A(n1283), .B(n1905), .C(n2126), .Y(n2487) );
  NAND2X1 U1833 ( .A(\mem<20><1> ), .B(n1285), .Y(n2127) );
  OAI21X1 U1834 ( .A(n1283), .B(n1908), .C(n2127), .Y(n2486) );
  NAND2X1 U1835 ( .A(\mem<20><2> ), .B(n1285), .Y(n2128) );
  OAI21X1 U1836 ( .A(n1283), .B(n1910), .C(n2128), .Y(n2485) );
  NAND2X1 U1837 ( .A(\mem<20><3> ), .B(n1285), .Y(n2129) );
  OAI21X1 U1838 ( .A(n1283), .B(n1912), .C(n2129), .Y(n2484) );
  NAND2X1 U1839 ( .A(\mem<20><4> ), .B(n1285), .Y(n2130) );
  OAI21X1 U1840 ( .A(n1283), .B(n1914), .C(n2130), .Y(n2483) );
  NAND2X1 U1841 ( .A(\mem<20><5> ), .B(n1285), .Y(n2131) );
  OAI21X1 U1842 ( .A(n1283), .B(n1916), .C(n2131), .Y(n2482) );
  NAND2X1 U1843 ( .A(\mem<20><6> ), .B(n1285), .Y(n2132) );
  OAI21X1 U1844 ( .A(n1283), .B(n1918), .C(n2132), .Y(n2481) );
  NAND2X1 U1845 ( .A(\mem<20><7> ), .B(n1285), .Y(n2133) );
  OAI21X1 U1846 ( .A(n1283), .B(n1920), .C(n2133), .Y(n2480) );
  NAND2X1 U1847 ( .A(\mem<20><8> ), .B(n1284), .Y(n2134) );
  OAI21X1 U1848 ( .A(n1283), .B(n1922), .C(n2134), .Y(n2479) );
  NAND2X1 U1849 ( .A(\mem<20><9> ), .B(n1284), .Y(n2135) );
  OAI21X1 U1850 ( .A(n1283), .B(n1924), .C(n2135), .Y(n2478) );
  NAND2X1 U1851 ( .A(\mem<20><10> ), .B(n1284), .Y(n2136) );
  OAI21X1 U1852 ( .A(n1283), .B(n1926), .C(n2136), .Y(n2477) );
  NAND2X1 U1853 ( .A(\mem<20><11> ), .B(n1284), .Y(n2137) );
  OAI21X1 U1854 ( .A(n1283), .B(n1928), .C(n2137), .Y(n2476) );
  NAND2X1 U1855 ( .A(\mem<20><12> ), .B(n1284), .Y(n2138) );
  OAI21X1 U1856 ( .A(n1283), .B(n1930), .C(n2138), .Y(n2475) );
  NAND2X1 U1857 ( .A(\mem<20><13> ), .B(n1284), .Y(n2139) );
  OAI21X1 U1858 ( .A(n1283), .B(n1932), .C(n2139), .Y(n2474) );
  NAND2X1 U1859 ( .A(\mem<20><14> ), .B(n1284), .Y(n2140) );
  OAI21X1 U1860 ( .A(n1283), .B(n1934), .C(n2140), .Y(n2473) );
  NAND2X1 U1861 ( .A(\mem<20><15> ), .B(n1284), .Y(n2141) );
  OAI21X1 U1862 ( .A(n1283), .B(n1936), .C(n2141), .Y(n2472) );
  OAI21X1 U1863 ( .A(n1287), .B(n1906), .C(n73), .Y(n2471) );
  OAI21X1 U1864 ( .A(n1287), .B(n1908), .C(n75), .Y(n2470) );
  OAI21X1 U1865 ( .A(n1287), .B(n1910), .C(n77), .Y(n2469) );
  OAI21X1 U1866 ( .A(n1287), .B(n1912), .C(n79), .Y(n2468) );
  OAI21X1 U1867 ( .A(n1287), .B(n1914), .C(n81), .Y(n2467) );
  OAI21X1 U1868 ( .A(n1287), .B(n1916), .C(n83), .Y(n2466) );
  OAI21X1 U1869 ( .A(n1287), .B(n1918), .C(n85), .Y(n2465) );
  OAI21X1 U1870 ( .A(n1287), .B(n1920), .C(n87), .Y(n2464) );
  OAI21X1 U1871 ( .A(n1287), .B(n1922), .C(n89), .Y(n2463) );
  OAI21X1 U1872 ( .A(n1287), .B(n1924), .C(n91), .Y(n2462) );
  OAI21X1 U1873 ( .A(n1287), .B(n1926), .C(n93), .Y(n2461) );
  OAI21X1 U1874 ( .A(n1287), .B(n1928), .C(n95), .Y(n2460) );
  OAI21X1 U1875 ( .A(n1287), .B(n1930), .C(n97), .Y(n2459) );
  OAI21X1 U1876 ( .A(n1287), .B(n1932), .C(n99), .Y(n2458) );
  OAI21X1 U1877 ( .A(n1287), .B(n1934), .C(n101), .Y(n2457) );
  OAI21X1 U1878 ( .A(n1287), .B(n1936), .C(n103), .Y(n2456) );
  OAI21X1 U1879 ( .A(n1289), .B(n1906), .C(n105), .Y(n2455) );
  OAI21X1 U1880 ( .A(n1289), .B(n1908), .C(n107), .Y(n2454) );
  OAI21X1 U1881 ( .A(n1289), .B(n1910), .C(n109), .Y(n2453) );
  OAI21X1 U1882 ( .A(n1289), .B(n1912), .C(n111), .Y(n2452) );
  OAI21X1 U1883 ( .A(n1289), .B(n1914), .C(n113), .Y(n2451) );
  OAI21X1 U1884 ( .A(n1289), .B(n1916), .C(n115), .Y(n2450) );
  OAI21X1 U1885 ( .A(n1289), .B(n1918), .C(n117), .Y(n2449) );
  OAI21X1 U1886 ( .A(n1289), .B(n1920), .C(n119), .Y(n2448) );
  OAI21X1 U1887 ( .A(n1289), .B(n1922), .C(n121), .Y(n2447) );
  OAI21X1 U1888 ( .A(n1289), .B(n1924), .C(n123), .Y(n2446) );
  OAI21X1 U1889 ( .A(n1289), .B(n1926), .C(n125), .Y(n2445) );
  OAI21X1 U1890 ( .A(n1289), .B(n1928), .C(n127), .Y(n2444) );
  OAI21X1 U1891 ( .A(n1289), .B(n1930), .C(n129), .Y(n2443) );
  OAI21X1 U1892 ( .A(n1289), .B(n1932), .C(n131), .Y(n2442) );
  OAI21X1 U1893 ( .A(n1289), .B(n1934), .C(n133), .Y(n2441) );
  OAI21X1 U1894 ( .A(n1289), .B(n1936), .C(n135), .Y(n2440) );
  OAI21X1 U1895 ( .A(n1291), .B(n1906), .C(n137), .Y(n2439) );
  OAI21X1 U1896 ( .A(n1291), .B(n1908), .C(n139), .Y(n2438) );
  OAI21X1 U1897 ( .A(n1291), .B(n1910), .C(n141), .Y(n2437) );
  OAI21X1 U1898 ( .A(n1291), .B(n1912), .C(n143), .Y(n2436) );
  OAI21X1 U1899 ( .A(n1291), .B(n1914), .C(n145), .Y(n2435) );
  OAI21X1 U1900 ( .A(n1291), .B(n1916), .C(n147), .Y(n2434) );
  OAI21X1 U1901 ( .A(n1291), .B(n1918), .C(n149), .Y(n2433) );
  OAI21X1 U1902 ( .A(n1291), .B(n1920), .C(n151), .Y(n2432) );
  OAI21X1 U1903 ( .A(n1291), .B(n1922), .C(n153), .Y(n2431) );
  OAI21X1 U1904 ( .A(n1291), .B(n1924), .C(n155), .Y(n2430) );
  OAI21X1 U1905 ( .A(n1291), .B(n1926), .C(n157), .Y(n2429) );
  OAI21X1 U1906 ( .A(n1291), .B(n1928), .C(n159), .Y(n2428) );
  OAI21X1 U1907 ( .A(n1291), .B(n1930), .C(n161), .Y(n2427) );
  OAI21X1 U1908 ( .A(n1291), .B(n1932), .C(n163), .Y(n2426) );
  OAI21X1 U1909 ( .A(n1291), .B(n1934), .C(n165), .Y(n2425) );
  OAI21X1 U1910 ( .A(n1291), .B(n1936), .C(n167), .Y(n2424) );
  OAI21X1 U1911 ( .A(n1864), .B(n1906), .C(n169), .Y(n2423) );
  OAI21X1 U1912 ( .A(n1864), .B(n1908), .C(n171), .Y(n2422) );
  OAI21X1 U1913 ( .A(n1864), .B(n1910), .C(n173), .Y(n2421) );
  OAI21X1 U1914 ( .A(n1864), .B(n1912), .C(n175), .Y(n2420) );
  OAI21X1 U1915 ( .A(n1864), .B(n1914), .C(n177), .Y(n2419) );
  OAI21X1 U1916 ( .A(n1864), .B(n1916), .C(n179), .Y(n2418) );
  OAI21X1 U1917 ( .A(n1864), .B(n1918), .C(n181), .Y(n2417) );
  OAI21X1 U1918 ( .A(n1864), .B(n1920), .C(n183), .Y(n2416) );
  OAI21X1 U1919 ( .A(n1864), .B(n1922), .C(n185), .Y(n2415) );
  OAI21X1 U1920 ( .A(n1864), .B(n1924), .C(n187), .Y(n2414) );
  OAI21X1 U1921 ( .A(n1864), .B(n1926), .C(n189), .Y(n2413) );
  OAI21X1 U1922 ( .A(n1864), .B(n1928), .C(n191), .Y(n2412) );
  OAI21X1 U1923 ( .A(n1864), .B(n1930), .C(n193), .Y(n2411) );
  OAI21X1 U1924 ( .A(n1864), .B(n1932), .C(n195), .Y(n2410) );
  OAI21X1 U1925 ( .A(n1864), .B(n1934), .C(n197), .Y(n2409) );
  OAI21X1 U1926 ( .A(n1864), .B(n1936), .C(n199), .Y(n2408) );
  NAND3X1 U1927 ( .A(n1817), .B(n2664), .C(n1944), .Y(n2142) );
  OAI21X1 U1928 ( .A(n1293), .B(n1906), .C(n201), .Y(n2407) );
  OAI21X1 U1929 ( .A(n1293), .B(n1908), .C(n203), .Y(n2406) );
  OAI21X1 U1930 ( .A(n1293), .B(n1910), .C(n205), .Y(n2405) );
  OAI21X1 U1931 ( .A(n1293), .B(n1912), .C(n207), .Y(n2404) );
  OAI21X1 U1932 ( .A(n1293), .B(n1914), .C(n209), .Y(n2403) );
  OAI21X1 U1933 ( .A(n1293), .B(n1916), .C(n211), .Y(n2402) );
  OAI21X1 U1934 ( .A(n1293), .B(n1918), .C(n213), .Y(n2401) );
  OAI21X1 U1935 ( .A(n1293), .B(n1920), .C(n216), .Y(n2400) );
  OAI21X1 U1936 ( .A(n1293), .B(n1922), .C(n218), .Y(n2399) );
  OAI21X1 U1937 ( .A(n1293), .B(n1924), .C(n220), .Y(n2398) );
  OAI21X1 U1938 ( .A(n1293), .B(n1926), .C(n222), .Y(n2397) );
  OAI21X1 U1939 ( .A(n1293), .B(n1928), .C(n224), .Y(n2396) );
  OAI21X1 U1940 ( .A(n1293), .B(n1930), .C(n226), .Y(n2395) );
  OAI21X1 U1941 ( .A(n1293), .B(n1932), .C(n228), .Y(n2394) );
  OAI21X1 U1942 ( .A(n1293), .B(n1934), .C(n230), .Y(n2393) );
  OAI21X1 U1943 ( .A(n1293), .B(n1936), .C(n232), .Y(n2392) );
  OAI21X1 U1944 ( .A(n1295), .B(n1906), .C(n234), .Y(n2391) );
  OAI21X1 U1945 ( .A(n1295), .B(n1908), .C(n236), .Y(n2390) );
  OAI21X1 U1946 ( .A(n1295), .B(n1910), .C(n238), .Y(n2389) );
  OAI21X1 U1947 ( .A(n1295), .B(n1912), .C(n240), .Y(n2388) );
  OAI21X1 U1948 ( .A(n1295), .B(n1914), .C(n242), .Y(n2387) );
  OAI21X1 U1949 ( .A(n1295), .B(n1916), .C(n244), .Y(n2386) );
  OAI21X1 U1950 ( .A(n1295), .B(n1918), .C(n246), .Y(n2385) );
  OAI21X1 U1951 ( .A(n1295), .B(n1920), .C(n248), .Y(n2384) );
  OAI21X1 U1952 ( .A(n1295), .B(n1922), .C(n250), .Y(n2383) );
  OAI21X1 U1953 ( .A(n1295), .B(n1924), .C(n252), .Y(n2382) );
  OAI21X1 U1954 ( .A(n1295), .B(n1926), .C(n254), .Y(n2381) );
  OAI21X1 U1955 ( .A(n1295), .B(n1928), .C(n256), .Y(n2380) );
  OAI21X1 U1956 ( .A(n1295), .B(n1930), .C(n258), .Y(n2379) );
  OAI21X1 U1957 ( .A(n1295), .B(n1932), .C(n260), .Y(n2378) );
  OAI21X1 U1958 ( .A(n1295), .B(n1934), .C(n262), .Y(n2377) );
  OAI21X1 U1959 ( .A(n1295), .B(n1936), .C(n264), .Y(n2376) );
  OAI21X1 U1960 ( .A(n1297), .B(n1906), .C(n266), .Y(n2375) );
  OAI21X1 U1961 ( .A(n1297), .B(n1908), .C(n268), .Y(n2374) );
  OAI21X1 U1962 ( .A(n1297), .B(n1910), .C(n270), .Y(n2373) );
  OAI21X1 U1963 ( .A(n1297), .B(n1912), .C(n272), .Y(n2372) );
  OAI21X1 U1964 ( .A(n1297), .B(n1914), .C(n274), .Y(n2371) );
  OAI21X1 U1965 ( .A(n1297), .B(n1916), .C(n276), .Y(n2370) );
  OAI21X1 U1966 ( .A(n1297), .B(n1918), .C(n278), .Y(n2369) );
  OAI21X1 U1967 ( .A(n1297), .B(n1920), .C(n280), .Y(n2368) );
  OAI21X1 U1968 ( .A(n1297), .B(n1922), .C(n282), .Y(n2367) );
  OAI21X1 U1969 ( .A(n1297), .B(n1924), .C(n284), .Y(n2366) );
  OAI21X1 U1970 ( .A(n1297), .B(n1926), .C(n286), .Y(n2365) );
  OAI21X1 U1971 ( .A(n1297), .B(n1928), .C(n288), .Y(n2364) );
  OAI21X1 U1972 ( .A(n1297), .B(n1930), .C(n290), .Y(n2363) );
  OAI21X1 U1973 ( .A(n1297), .B(n1932), .C(n292), .Y(n2362) );
  OAI21X1 U1974 ( .A(n1297), .B(n1934), .C(n294), .Y(n2361) );
  OAI21X1 U1975 ( .A(n1297), .B(n1936), .C(n296), .Y(n2360) );
  OAI21X1 U1976 ( .A(n1299), .B(n1906), .C(n298), .Y(n2359) );
  OAI21X1 U1977 ( .A(n1299), .B(n1908), .C(n300), .Y(n2358) );
  OAI21X1 U1978 ( .A(n1299), .B(n1910), .C(n302), .Y(n2357) );
  OAI21X1 U1979 ( .A(n1299), .B(n1912), .C(n304), .Y(n2356) );
  OAI21X1 U1980 ( .A(n1299), .B(n1914), .C(n306), .Y(n2355) );
  OAI21X1 U1981 ( .A(n1299), .B(n1916), .C(n308), .Y(n2354) );
  OAI21X1 U1982 ( .A(n1299), .B(n1918), .C(n310), .Y(n2353) );
  OAI21X1 U1983 ( .A(n1299), .B(n1920), .C(n312), .Y(n2352) );
  OAI21X1 U1984 ( .A(n1299), .B(n1922), .C(n314), .Y(n2351) );
  OAI21X1 U1985 ( .A(n1299), .B(n1924), .C(n316), .Y(n2350) );
  OAI21X1 U1986 ( .A(n1299), .B(n1926), .C(n318), .Y(n2349) );
  OAI21X1 U1987 ( .A(n1299), .B(n1928), .C(n320), .Y(n2348) );
  OAI21X1 U1988 ( .A(n1299), .B(n1930), .C(n322), .Y(n2347) );
  OAI21X1 U1989 ( .A(n1299), .B(n1932), .C(n324), .Y(n2346) );
  OAI21X1 U1990 ( .A(n1299), .B(n1934), .C(n326), .Y(n2345) );
  OAI21X1 U1991 ( .A(n1299), .B(n1936), .C(n328), .Y(n2344) );
  OAI21X1 U1992 ( .A(n1301), .B(n1906), .C(n330), .Y(n2343) );
  OAI21X1 U1993 ( .A(n1301), .B(n1907), .C(n332), .Y(n2342) );
  OAI21X1 U1994 ( .A(n1301), .B(n1909), .C(n334), .Y(n2341) );
  OAI21X1 U1995 ( .A(n1301), .B(n1911), .C(n336), .Y(n2340) );
  OAI21X1 U1996 ( .A(n1301), .B(n1913), .C(n338), .Y(n2339) );
  OAI21X1 U1997 ( .A(n1301), .B(n1915), .C(n340), .Y(n2338) );
  OAI21X1 U1998 ( .A(n1301), .B(n1917), .C(n342), .Y(n2337) );
  OAI21X1 U1999 ( .A(n1301), .B(n1919), .C(n344), .Y(n2336) );
  OAI21X1 U2000 ( .A(n1301), .B(n1921), .C(n346), .Y(n2335) );
  OAI21X1 U2001 ( .A(n1301), .B(n1923), .C(n348), .Y(n2334) );
  OAI21X1 U2002 ( .A(n1301), .B(n1925), .C(n350), .Y(n2333) );
  OAI21X1 U2003 ( .A(n1301), .B(n1927), .C(n352), .Y(n2332) );
  OAI21X1 U2004 ( .A(n1301), .B(n1929), .C(n354), .Y(n2331) );
  OAI21X1 U2005 ( .A(n1301), .B(n1931), .C(n356), .Y(n2330) );
  OAI21X1 U2006 ( .A(n1301), .B(n1933), .C(n358), .Y(n2329) );
  OAI21X1 U2007 ( .A(n1301), .B(n1935), .C(n360), .Y(n2328) );
  OAI21X1 U2008 ( .A(n1303), .B(n1906), .C(n362), .Y(n2327) );
  OAI21X1 U2009 ( .A(n1303), .B(n1907), .C(n364), .Y(n2326) );
  OAI21X1 U2010 ( .A(n1303), .B(n1909), .C(n366), .Y(n2325) );
  OAI21X1 U2011 ( .A(n1303), .B(n1911), .C(n368), .Y(n2324) );
  OAI21X1 U2012 ( .A(n1303), .B(n1913), .C(n370), .Y(n2323) );
  OAI21X1 U2013 ( .A(n1303), .B(n1915), .C(n372), .Y(n2322) );
  OAI21X1 U2014 ( .A(n1303), .B(n1917), .C(n374), .Y(n2321) );
  OAI21X1 U2015 ( .A(n1303), .B(n1919), .C(n376), .Y(n2320) );
  OAI21X1 U2016 ( .A(n1303), .B(n1921), .C(n378), .Y(n2319) );
  OAI21X1 U2017 ( .A(n1303), .B(n1923), .C(n380), .Y(n2318) );
  OAI21X1 U2018 ( .A(n1303), .B(n1925), .C(n382), .Y(n2317) );
  OAI21X1 U2019 ( .A(n1303), .B(n1927), .C(n384), .Y(n2316) );
  OAI21X1 U2020 ( .A(n1303), .B(n1929), .C(n386), .Y(n2315) );
  OAI21X1 U2021 ( .A(n1303), .B(n1931), .C(n388), .Y(n2314) );
  OAI21X1 U2022 ( .A(n1303), .B(n1933), .C(n390), .Y(n2313) );
  OAI21X1 U2023 ( .A(n1303), .B(n1935), .C(n392), .Y(n2312) );
  OAI21X1 U2024 ( .A(n1305), .B(n1906), .C(n394), .Y(n2311) );
  OAI21X1 U2025 ( .A(n1305), .B(n1907), .C(n396), .Y(n2310) );
  OAI21X1 U2026 ( .A(n1305), .B(n1909), .C(n398), .Y(n2309) );
  OAI21X1 U2027 ( .A(n1305), .B(n1911), .C(n400), .Y(n2308) );
  OAI21X1 U2028 ( .A(n1305), .B(n1913), .C(n402), .Y(n2307) );
  OAI21X1 U2029 ( .A(n1305), .B(n1915), .C(n404), .Y(n2306) );
  OAI21X1 U2030 ( .A(n1305), .B(n1917), .C(n406), .Y(n2305) );
  OAI21X1 U2031 ( .A(n1305), .B(n1919), .C(n408), .Y(n2304) );
  OAI21X1 U2032 ( .A(n1305), .B(n1921), .C(n410), .Y(n2303) );
  OAI21X1 U2033 ( .A(n1305), .B(n1923), .C(n412), .Y(n2302) );
  OAI21X1 U2034 ( .A(n1305), .B(n1925), .C(n414), .Y(n2301) );
  OAI21X1 U2035 ( .A(n1305), .B(n1927), .C(n416), .Y(n2300) );
  OAI21X1 U2036 ( .A(n1305), .B(n1929), .C(n418), .Y(n2299) );
  OAI21X1 U2037 ( .A(n1305), .B(n1931), .C(n420), .Y(n2298) );
  OAI21X1 U2038 ( .A(n1305), .B(n1933), .C(n422), .Y(n2297) );
  OAI21X1 U2039 ( .A(n1305), .B(n1935), .C(n424), .Y(n2296) );
  OAI21X1 U2040 ( .A(n1881), .B(n1906), .C(n426), .Y(n2295) );
  OAI21X1 U2041 ( .A(n1881), .B(n1907), .C(n428), .Y(n2294) );
  OAI21X1 U2042 ( .A(n1881), .B(n1909), .C(n430), .Y(n2293) );
  OAI21X1 U2043 ( .A(n1881), .B(n1911), .C(n432), .Y(n2292) );
  OAI21X1 U2044 ( .A(n1881), .B(n1913), .C(n434), .Y(n2291) );
  OAI21X1 U2045 ( .A(n1881), .B(n1915), .C(n436), .Y(n2290) );
  OAI21X1 U2046 ( .A(n1881), .B(n1917), .C(n438), .Y(n2289) );
  OAI21X1 U2047 ( .A(n1881), .B(n1919), .C(n440), .Y(n2288) );
  OAI21X1 U2048 ( .A(n1881), .B(n1921), .C(n442), .Y(n2287) );
  OAI21X1 U2049 ( .A(n1881), .B(n1923), .C(n444), .Y(n2286) );
  OAI21X1 U2050 ( .A(n1881), .B(n1925), .C(n446), .Y(n2285) );
  OAI21X1 U2051 ( .A(n1881), .B(n1927), .C(n448), .Y(n2284) );
  OAI21X1 U2052 ( .A(n1881), .B(n1929), .C(n450), .Y(n2283) );
  OAI21X1 U2053 ( .A(n1881), .B(n1931), .C(n452), .Y(n2282) );
  OAI21X1 U2054 ( .A(n1881), .B(n1933), .C(n454), .Y(n2281) );
  OAI21X1 U2055 ( .A(n1881), .B(n1935), .C(n456), .Y(n2280) );
  NAND3X1 U2056 ( .A(n1943), .B(n2664), .C(n1944), .Y(n2144) );
  OAI21X1 U2057 ( .A(n1307), .B(n1905), .C(n458), .Y(n2279) );
  OAI21X1 U2058 ( .A(n1307), .B(n1907), .C(n460), .Y(n2278) );
  OAI21X1 U2059 ( .A(n1307), .B(n1909), .C(n462), .Y(n2277) );
  OAI21X1 U2060 ( .A(n1307), .B(n1911), .C(n464), .Y(n2276) );
  OAI21X1 U2061 ( .A(n1307), .B(n1913), .C(n466), .Y(n2275) );
  OAI21X1 U2062 ( .A(n1307), .B(n1915), .C(n468), .Y(n2274) );
  OAI21X1 U2063 ( .A(n1307), .B(n1917), .C(n470), .Y(n2273) );
  OAI21X1 U2064 ( .A(n1307), .B(n1919), .C(n472), .Y(n2272) );
  OAI21X1 U2065 ( .A(n1307), .B(n1921), .C(n474), .Y(n2271) );
  OAI21X1 U2066 ( .A(n1307), .B(n1923), .C(n476), .Y(n2270) );
  OAI21X1 U2067 ( .A(n1307), .B(n1925), .C(n478), .Y(n2269) );
  OAI21X1 U2068 ( .A(n1307), .B(n1927), .C(n480), .Y(n2268) );
  OAI21X1 U2069 ( .A(n1307), .B(n1929), .C(n482), .Y(n2267) );
  OAI21X1 U2070 ( .A(n1307), .B(n1931), .C(n484), .Y(n2266) );
  OAI21X1 U2071 ( .A(n1307), .B(n1933), .C(n486), .Y(n2265) );
  OAI21X1 U2072 ( .A(n1307), .B(n1935), .C(n488), .Y(n2264) );
  OAI21X1 U2073 ( .A(n1309), .B(n1906), .C(n490), .Y(n2263) );
  OAI21X1 U2074 ( .A(n1309), .B(n1907), .C(n492), .Y(n2262) );
  OAI21X1 U2075 ( .A(n1309), .B(n1909), .C(n494), .Y(n2261) );
  OAI21X1 U2076 ( .A(n1309), .B(n1911), .C(n496), .Y(n2260) );
  OAI21X1 U2077 ( .A(n1309), .B(n1913), .C(n498), .Y(n2259) );
  OAI21X1 U2078 ( .A(n1309), .B(n1915), .C(n500), .Y(n2258) );
  OAI21X1 U2079 ( .A(n1309), .B(n1917), .C(n502), .Y(n2257) );
  OAI21X1 U2080 ( .A(n1309), .B(n1919), .C(n504), .Y(n2256) );
  OAI21X1 U2081 ( .A(n1309), .B(n1921), .C(n506), .Y(n2255) );
  OAI21X1 U2082 ( .A(n1309), .B(n1923), .C(n508), .Y(n2254) );
  OAI21X1 U2083 ( .A(n1309), .B(n1925), .C(n510), .Y(n2253) );
  OAI21X1 U2084 ( .A(n1309), .B(n1927), .C(n512), .Y(n2252) );
  OAI21X1 U2085 ( .A(n1309), .B(n1929), .C(n514), .Y(n2251) );
  OAI21X1 U2086 ( .A(n1309), .B(n1931), .C(n516), .Y(n2250) );
  OAI21X1 U2087 ( .A(n1309), .B(n1933), .C(n518), .Y(n2249) );
  OAI21X1 U2088 ( .A(n1309), .B(n1935), .C(n520), .Y(n2248) );
  OAI21X1 U2089 ( .A(n1311), .B(n1905), .C(n522), .Y(n2247) );
  OAI21X1 U2090 ( .A(n1311), .B(n1907), .C(n524), .Y(n2246) );
  OAI21X1 U2091 ( .A(n1311), .B(n1909), .C(n526), .Y(n2245) );
  OAI21X1 U2092 ( .A(n1311), .B(n1911), .C(n528), .Y(n2244) );
  OAI21X1 U2093 ( .A(n1311), .B(n1913), .C(n530), .Y(n2243) );
  OAI21X1 U2094 ( .A(n1311), .B(n1915), .C(n532), .Y(n2242) );
  OAI21X1 U2095 ( .A(n1311), .B(n1917), .C(n534), .Y(n2241) );
  OAI21X1 U2096 ( .A(n1311), .B(n1919), .C(n536), .Y(n2240) );
  OAI21X1 U2097 ( .A(n1311), .B(n1921), .C(n538), .Y(n2239) );
  OAI21X1 U2098 ( .A(n1311), .B(n1923), .C(n540), .Y(n2238) );
  OAI21X1 U2099 ( .A(n1311), .B(n1925), .C(n542), .Y(n2237) );
  OAI21X1 U2100 ( .A(n1311), .B(n1927), .C(n544), .Y(n2236) );
  OAI21X1 U2101 ( .A(n1311), .B(n1929), .C(n546), .Y(n2235) );
  OAI21X1 U2102 ( .A(n1311), .B(n1931), .C(n548), .Y(n2234) );
  OAI21X1 U2103 ( .A(n1311), .B(n1933), .C(n550), .Y(n2233) );
  OAI21X1 U2104 ( .A(n1311), .B(n1935), .C(n552), .Y(n2232) );
  OAI21X1 U2105 ( .A(n1313), .B(n1906), .C(n554), .Y(n2231) );
  OAI21X1 U2106 ( .A(n1313), .B(n1907), .C(n556), .Y(n2230) );
  OAI21X1 U2107 ( .A(n1313), .B(n1909), .C(n558), .Y(n2229) );
  OAI21X1 U2108 ( .A(n1313), .B(n1911), .C(n560), .Y(n2228) );
  OAI21X1 U2109 ( .A(n1313), .B(n1913), .C(n562), .Y(n2227) );
  OAI21X1 U2110 ( .A(n1313), .B(n1915), .C(n564), .Y(n2226) );
  OAI21X1 U2111 ( .A(n1313), .B(n1917), .C(n566), .Y(n2225) );
  OAI21X1 U2112 ( .A(n1313), .B(n1919), .C(n568), .Y(n2224) );
  OAI21X1 U2113 ( .A(n1313), .B(n1921), .C(n570), .Y(n2223) );
  OAI21X1 U2114 ( .A(n1313), .B(n1923), .C(n572), .Y(n2222) );
  OAI21X1 U2115 ( .A(n1313), .B(n1925), .C(n574), .Y(n2221) );
  OAI21X1 U2116 ( .A(n1313), .B(n1927), .C(n576), .Y(n2220) );
  OAI21X1 U2117 ( .A(n1313), .B(n1929), .C(n578), .Y(n2219) );
  OAI21X1 U2118 ( .A(n1313), .B(n1931), .C(n580), .Y(n2218) );
  OAI21X1 U2119 ( .A(n1313), .B(n1933), .C(n582), .Y(n2217) );
  OAI21X1 U2120 ( .A(n1313), .B(n1935), .C(n584), .Y(n2216) );
  OAI21X1 U2121 ( .A(n1315), .B(n1905), .C(n586), .Y(n2215) );
  OAI21X1 U2122 ( .A(n1315), .B(n1907), .C(n588), .Y(n2214) );
  OAI21X1 U2123 ( .A(n1315), .B(n1909), .C(n590), .Y(n2213) );
  OAI21X1 U2124 ( .A(n1315), .B(n1911), .C(n592), .Y(n2212) );
  OAI21X1 U2125 ( .A(n1315), .B(n1913), .C(n594), .Y(n2211) );
  OAI21X1 U2126 ( .A(n1315), .B(n1915), .C(n596), .Y(n2210) );
  OAI21X1 U2127 ( .A(n1315), .B(n1917), .C(n598), .Y(n2209) );
  OAI21X1 U2128 ( .A(n1315), .B(n1919), .C(n600), .Y(n2208) );
  OAI21X1 U2129 ( .A(n1315), .B(n1921), .C(n602), .Y(n2207) );
  OAI21X1 U2130 ( .A(n1315), .B(n1923), .C(n604), .Y(n2206) );
  OAI21X1 U2131 ( .A(n1315), .B(n1925), .C(n606), .Y(n2205) );
  OAI21X1 U2132 ( .A(n1315), .B(n1927), .C(n608), .Y(n2204) );
  OAI21X1 U2133 ( .A(n1315), .B(n1929), .C(n610), .Y(n2203) );
  OAI21X1 U2134 ( .A(n1315), .B(n1931), .C(n612), .Y(n2202) );
  OAI21X1 U2135 ( .A(n1315), .B(n1933), .C(n614), .Y(n2201) );
  OAI21X1 U2136 ( .A(n1315), .B(n1935), .C(n616), .Y(n2200) );
  OAI21X1 U2137 ( .A(n1317), .B(n1906), .C(n618), .Y(n2199) );
  OAI21X1 U2138 ( .A(n1317), .B(n1907), .C(n620), .Y(n2198) );
  OAI21X1 U2139 ( .A(n1317), .B(n1909), .C(n622), .Y(n2197) );
  OAI21X1 U2140 ( .A(n1317), .B(n1911), .C(n624), .Y(n2196) );
  OAI21X1 U2141 ( .A(n1317), .B(n1913), .C(n626), .Y(n2195) );
  OAI21X1 U2142 ( .A(n1317), .B(n1915), .C(n628), .Y(n2194) );
  OAI21X1 U2143 ( .A(n1317), .B(n1917), .C(n630), .Y(n2193) );
  OAI21X1 U2144 ( .A(n1317), .B(n1919), .C(n632), .Y(n2192) );
  OAI21X1 U2145 ( .A(n1317), .B(n1921), .C(n634), .Y(n2191) );
  OAI21X1 U2146 ( .A(n1317), .B(n1923), .C(n636), .Y(n2190) );
  OAI21X1 U2147 ( .A(n1317), .B(n1925), .C(n638), .Y(n2189) );
  OAI21X1 U2148 ( .A(n1317), .B(n1927), .C(n640), .Y(n2188) );
  OAI21X1 U2149 ( .A(n1317), .B(n1929), .C(n642), .Y(n2187) );
  OAI21X1 U2150 ( .A(n1317), .B(n1931), .C(n644), .Y(n2186) );
  OAI21X1 U2151 ( .A(n1317), .B(n1933), .C(n646), .Y(n2185) );
  OAI21X1 U2152 ( .A(n1317), .B(n1935), .C(n648), .Y(n2184) );
  OAI21X1 U2153 ( .A(n1319), .B(n1905), .C(n650), .Y(n2183) );
  OAI21X1 U2154 ( .A(n1319), .B(n1907), .C(n1164), .Y(n2182) );
  OAI21X1 U2155 ( .A(n1319), .B(n1909), .C(n1166), .Y(n2181) );
  OAI21X1 U2156 ( .A(n1319), .B(n1911), .C(n1168), .Y(n2180) );
  OAI21X1 U2157 ( .A(n1319), .B(n1913), .C(n1170), .Y(n2179) );
  OAI21X1 U2158 ( .A(n1319), .B(n1915), .C(n1172), .Y(n2178) );
  OAI21X1 U2159 ( .A(n1319), .B(n1917), .C(n1174), .Y(n2177) );
  OAI21X1 U2160 ( .A(n1319), .B(n1919), .C(n1176), .Y(n2176) );
  OAI21X1 U2161 ( .A(n1319), .B(n1921), .C(n1178), .Y(n2175) );
  OAI21X1 U2162 ( .A(n1319), .B(n1923), .C(n1180), .Y(n2174) );
  OAI21X1 U2163 ( .A(n1319), .B(n1925), .C(n1182), .Y(n2173) );
  OAI21X1 U2164 ( .A(n1319), .B(n1927), .C(n1184), .Y(n2172) );
  OAI21X1 U2165 ( .A(n1319), .B(n1929), .C(n1186), .Y(n2171) );
  OAI21X1 U2166 ( .A(n1319), .B(n1931), .C(n1188), .Y(n2170) );
  OAI21X1 U2167 ( .A(n1319), .B(n1933), .C(n1190), .Y(n2169) );
  OAI21X1 U2168 ( .A(n1319), .B(n1935), .C(n1192), .Y(n2168) );
  OAI21X1 U2169 ( .A(n1898), .B(n1906), .C(n1194), .Y(n2167) );
  OAI21X1 U2170 ( .A(n1898), .B(n1907), .C(n1196), .Y(n2166) );
  OAI21X1 U2171 ( .A(n1898), .B(n1909), .C(n1198), .Y(n2165) );
  OAI21X1 U2172 ( .A(n1898), .B(n1911), .C(n1200), .Y(n2164) );
  OAI21X1 U2173 ( .A(n1898), .B(n1913), .C(n1202), .Y(n2163) );
  OAI21X1 U2174 ( .A(n1898), .B(n1915), .C(n1204), .Y(n2162) );
  OAI21X1 U2175 ( .A(n1898), .B(n1917), .C(n1206), .Y(n2161) );
  OAI21X1 U2176 ( .A(n1898), .B(n1919), .C(n1208), .Y(n2160) );
  OAI21X1 U2177 ( .A(n1898), .B(n1921), .C(n1210), .Y(n2159) );
  OAI21X1 U2178 ( .A(n1898), .B(n1923), .C(n1212), .Y(n2158) );
  OAI21X1 U2179 ( .A(n1898), .B(n1925), .C(n1214), .Y(n2157) );
  OAI21X1 U2180 ( .A(n1898), .B(n1927), .C(n1216), .Y(n2156) );
  OAI21X1 U2181 ( .A(n1898), .B(n1929), .C(n1218), .Y(n2155) );
  OAI21X1 U2182 ( .A(n1898), .B(n1931), .C(n1220), .Y(n2154) );
  OAI21X1 U2183 ( .A(n1898), .B(n1933), .C(n1222), .Y(n2153) );
  OAI21X1 U2184 ( .A(n1898), .B(n1935), .C(n1224), .Y(n2152) );
endmodule


module memc_Size5 ( .data_out({\data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), .addr({\addr<7> , \addr<6> , \addr<5> , 
        \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), .data_in({
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        write, clk, rst, createdump, .file_id({\file_id<4> , \file_id<3> , 
        \file_id<2> , \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<4> , \data_in<3> , \data_in<2> ,
         \data_in<1> , \data_in<0> , write, clk, rst, createdump, \file_id<4> ,
         \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> ,
         \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><4> , \mem<0><3> , \mem<0><2> ,
         \mem<0><1> , \mem<0><0> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><4> , \mem<2><3> , \mem<2><2> ,
         \mem<2><1> , \mem<2><0> , \mem<3><4> , \mem<3><3> , \mem<3><2> ,
         \mem<3><1> , \mem<3><0> , \mem<4><4> , \mem<4><3> , \mem<4><2> ,
         \mem<4><1> , \mem<4><0> , \mem<5><4> , \mem<5><3> , \mem<5><2> ,
         \mem<5><1> , \mem<5><0> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><4> , \mem<7><3> , \mem<7><2> ,
         \mem<7><1> , \mem<7><0> , \mem<8><4> , \mem<8><3> , \mem<8><2> ,
         \mem<8><1> , \mem<8><0> , \mem<9><4> , \mem<9><3> , \mem<9><2> ,
         \mem<9><1> , \mem<9><0> , \mem<10><4> , \mem<10><3> , \mem<10><2> ,
         \mem<10><1> , \mem<10><0> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><4> , \mem<12><3> , \mem<12><2> ,
         \mem<12><1> , \mem<12><0> , \mem<13><4> , \mem<13><3> , \mem<13><2> ,
         \mem<13><1> , \mem<13><0> , \mem<14><4> , \mem<14><3> , \mem<14><2> ,
         \mem<14><1> , \mem<14><0> , \mem<15><4> , \mem<15><3> , \mem<15><2> ,
         \mem<15><1> , \mem<15><0> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><4> , \mem<17><3> , \mem<17><2> ,
         \mem<17><1> , \mem<17><0> , \mem<18><4> , \mem<18><3> , \mem<18><2> ,
         \mem<18><1> , \mem<18><0> , \mem<19><4> , \mem<19><3> , \mem<19><2> ,
         \mem<19><1> , \mem<19><0> , \mem<20><4> , \mem<20><3> , \mem<20><2> ,
         \mem<20><1> , \mem<20><0> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><4> , \mem<22><3> , \mem<22><2> ,
         \mem<22><1> , \mem<22><0> , \mem<23><4> , \mem<23><3> , \mem<23><2> ,
         \mem<23><1> , \mem<23><0> , \mem<24><4> , \mem<24><3> , \mem<24><2> ,
         \mem<24><1> , \mem<24><0> , \mem<25><4> , \mem<25><3> , \mem<25><2> ,
         \mem<25><1> , \mem<25><0> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><4> , \mem<27><3> , \mem<27><2> ,
         \mem<27><1> , \mem<27><0> , \mem<28><4> , \mem<28><3> , \mem<28><2> ,
         \mem<28><1> , \mem<28><0> , \mem<29><4> , \mem<29><3> , \mem<29><2> ,
         \mem<29><1> , \mem<29><0> , \mem<30><4> , \mem<30><3> , \mem<30><2> ,
         \mem<30><1> , \mem<30><0> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , N17, N18, N19, N20, N21, n46, n49, n51,
         n53, n55, n56, n57, n59, n61, n62, n63, n64, n65, n67, n69, n70, n71,
         n72, n73, n75, n77, n78, n79, n80, n81, n83, n85, n86, n87, n88, n89,
         n91, n93, n94, n95, n96, n97, n99, n101, n102, n103, n104, n105, n107,
         n109, n110, n111, n112, n113, n114, n115, n117, n119, n120, n121,
         n122, n124, n126, n127, n128, n129, n131, n133, n134, n135, n136,
         n138, n140, n141, n142, n143, n145, n147, n148, n149, n150, n152,
         n154, n155, n156, n157, n159, n161, n162, n163, n164, n166, n168,
         n169, n170, n171, n172, n174, n176, n177, n178, n179, n181, n183,
         n184, n185, n186, n188, n190, n191, n192, n193, n195, n197, n198,
         n199, n200, n202, n204, n205, n206, n207, n209, n211, n212, n213,
         n214, n216, n218, n219, n220, n221, n223, n225, n226, n227, n228,
         n229, n231, n233, n234, n235, n236, n238, n240, n241, n242, n243,
         n245, n247, n248, n249, n250, n252, n254, n255, n256, n257, n259,
         n261, n262, n263, n264, n266, n268, n269, n270, n271, n273, n275,
         n276, n277, n278, n280, n282, n283, n284, n285, n286, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n47, n48, n50, n52, n54, n58, n60, n66,
         n68, n74, n76, n82, n84, n90, n92, n98, n100, n106, n108, n116, n118,
         n123, n125, n130, n132, n137, n139, n144, n146, n151, n153, n158,
         n160, n165, n167, n173, n175, n180, n182, n187, n189, n194, n196,
         n201, n203, n208, n210, n215, n217, n222, n224, n230, n232, n237,
         n239, n244, n246, n251, n253, n258, n260, n265, n267, n272, n274,
         n279, n281, n287, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><4>  ( .D(n447), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n446), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n445), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n444), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n443), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n442), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n441), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n440), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n439), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n438), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n437), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n436), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n435), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n434), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n433), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n432), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n431), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n430), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n429), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n428), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n427), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n426), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n425), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n424), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n423), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n422), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n421), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n420), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n419), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n418), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n417), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n416), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n415), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n414), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n413), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n412), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n411), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n410), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n409), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n408), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n407), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n406), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n405), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n404), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n403), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n402), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n401), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n400), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n399), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n398), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n397), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n396), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n395), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n394), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n393), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n392), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n391), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n390), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n389), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n388), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n387), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n386), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n385), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n384), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n383), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n382), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n381), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n380), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n379), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n378), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n377), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n376), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n375), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n374), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n373), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n372), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n371), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n370), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n369), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n368), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n367), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n366), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n365), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n364), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n363), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n362), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n361), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n360), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n359), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n358), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n357), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n356), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n355), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n354), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n353), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n352), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n351), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n350), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n349), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n348), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n347), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n346), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n345), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n344), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n343), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n342), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n341), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n340), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n339), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n338), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n337), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n336), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n335), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n334), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n333), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n332), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n331), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n330), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n329), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n328), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n327), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n326), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n325), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n324), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n323), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n322), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n321), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n320), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n319), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n318), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n317), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n316), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n315), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n314), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n313), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n312), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n311), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n310), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n309), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n308), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n307), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n306), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n305), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n304), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n303), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n302), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n301), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n300), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n299), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n298), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n297), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n296), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n295), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n294), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n293), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n292), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n291), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n290), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n289), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n288), .CLK(clk), .Q(\mem<31><0> ) );
  OAI21X1 U50 ( .A(n173), .B(n663), .C(n46), .Y(n288) );
  NAND2X1 U51 ( .A(\mem<31><0> ), .B(n167), .Y(n46) );
  OAI21X1 U52 ( .A(n173), .B(n661), .C(n49), .Y(n289) );
  NAND2X1 U53 ( .A(\mem<31><1> ), .B(n167), .Y(n49) );
  OAI21X1 U54 ( .A(n173), .B(n659), .C(n51), .Y(n290) );
  NAND2X1 U55 ( .A(\mem<31><2> ), .B(n167), .Y(n51) );
  OAI21X1 U56 ( .A(n173), .B(n657), .C(n53), .Y(n291) );
  NAND2X1 U57 ( .A(\mem<31><3> ), .B(n167), .Y(n53) );
  OAI21X1 U58 ( .A(n173), .B(n655), .C(n55), .Y(n292) );
  NAND2X1 U59 ( .A(\mem<31><4> ), .B(n167), .Y(n55) );
  OAI21X1 U62 ( .A(n663), .B(n477), .C(n59), .Y(n293) );
  NAND2X1 U63 ( .A(\mem<30><0> ), .B(n160), .Y(n59) );
  OAI21X1 U64 ( .A(n661), .B(n477), .C(n61), .Y(n294) );
  NAND2X1 U65 ( .A(\mem<30><1> ), .B(n160), .Y(n61) );
  OAI21X1 U66 ( .A(n659), .B(n477), .C(n62), .Y(n295) );
  NAND2X1 U67 ( .A(\mem<30><2> ), .B(n160), .Y(n62) );
  OAI21X1 U68 ( .A(n657), .B(n477), .C(n63), .Y(n296) );
  NAND2X1 U69 ( .A(\mem<30><3> ), .B(n160), .Y(n63) );
  OAI21X1 U70 ( .A(n655), .B(n477), .C(n64), .Y(n297) );
  NAND2X1 U71 ( .A(\mem<30><4> ), .B(n160), .Y(n64) );
  OAI21X1 U74 ( .A(n663), .B(n475), .C(n67), .Y(n298) );
  NAND2X1 U75 ( .A(\mem<29><0> ), .B(n153), .Y(n67) );
  OAI21X1 U76 ( .A(n661), .B(n475), .C(n69), .Y(n299) );
  NAND2X1 U77 ( .A(\mem<29><1> ), .B(n153), .Y(n69) );
  OAI21X1 U78 ( .A(n659), .B(n475), .C(n70), .Y(n300) );
  NAND2X1 U79 ( .A(\mem<29><2> ), .B(n153), .Y(n70) );
  OAI21X1 U80 ( .A(n657), .B(n475), .C(n71), .Y(n301) );
  NAND2X1 U81 ( .A(\mem<29><3> ), .B(n153), .Y(n71) );
  OAI21X1 U82 ( .A(n655), .B(n475), .C(n72), .Y(n302) );
  NAND2X1 U83 ( .A(\mem<29><4> ), .B(n153), .Y(n72) );
  OAI21X1 U86 ( .A(n663), .B(n473), .C(n75), .Y(n303) );
  NAND2X1 U87 ( .A(\mem<28><0> ), .B(n146), .Y(n75) );
  OAI21X1 U88 ( .A(n661), .B(n473), .C(n77), .Y(n304) );
  NAND2X1 U89 ( .A(\mem<28><1> ), .B(n146), .Y(n77) );
  OAI21X1 U90 ( .A(n659), .B(n473), .C(n78), .Y(n305) );
  NAND2X1 U91 ( .A(\mem<28><2> ), .B(n146), .Y(n78) );
  OAI21X1 U92 ( .A(n657), .B(n473), .C(n79), .Y(n306) );
  NAND2X1 U93 ( .A(\mem<28><3> ), .B(n146), .Y(n79) );
  OAI21X1 U94 ( .A(n655), .B(n473), .C(n80), .Y(n307) );
  NAND2X1 U95 ( .A(\mem<28><4> ), .B(n146), .Y(n80) );
  OAI21X1 U98 ( .A(n663), .B(n471), .C(n83), .Y(n308) );
  NAND2X1 U99 ( .A(\mem<27><0> ), .B(n139), .Y(n83) );
  OAI21X1 U100 ( .A(n661), .B(n471), .C(n85), .Y(n309) );
  NAND2X1 U101 ( .A(\mem<27><1> ), .B(n139), .Y(n85) );
  OAI21X1 U102 ( .A(n659), .B(n471), .C(n86), .Y(n310) );
  NAND2X1 U103 ( .A(\mem<27><2> ), .B(n139), .Y(n86) );
  OAI21X1 U104 ( .A(n657), .B(n471), .C(n87), .Y(n311) );
  NAND2X1 U105 ( .A(\mem<27><3> ), .B(n139), .Y(n87) );
  OAI21X1 U106 ( .A(n655), .B(n471), .C(n88), .Y(n312) );
  NAND2X1 U107 ( .A(\mem<27><4> ), .B(n139), .Y(n88) );
  OAI21X1 U110 ( .A(n663), .B(n469), .C(n91), .Y(n313) );
  NAND2X1 U111 ( .A(\mem<26><0> ), .B(n132), .Y(n91) );
  OAI21X1 U112 ( .A(n661), .B(n469), .C(n93), .Y(n314) );
  NAND2X1 U113 ( .A(\mem<26><1> ), .B(n132), .Y(n93) );
  OAI21X1 U114 ( .A(n659), .B(n469), .C(n94), .Y(n315) );
  NAND2X1 U115 ( .A(\mem<26><2> ), .B(n132), .Y(n94) );
  OAI21X1 U116 ( .A(n657), .B(n469), .C(n95), .Y(n316) );
  NAND2X1 U117 ( .A(\mem<26><3> ), .B(n132), .Y(n95) );
  OAI21X1 U118 ( .A(n655), .B(n469), .C(n96), .Y(n317) );
  NAND2X1 U119 ( .A(\mem<26><4> ), .B(n132), .Y(n96) );
  OAI21X1 U122 ( .A(n663), .B(n467), .C(n99), .Y(n318) );
  NAND2X1 U123 ( .A(\mem<25><0> ), .B(n125), .Y(n99) );
  OAI21X1 U124 ( .A(n661), .B(n467), .C(n101), .Y(n319) );
  NAND2X1 U125 ( .A(\mem<25><1> ), .B(n125), .Y(n101) );
  OAI21X1 U126 ( .A(n659), .B(n467), .C(n102), .Y(n320) );
  NAND2X1 U127 ( .A(\mem<25><2> ), .B(n125), .Y(n102) );
  OAI21X1 U128 ( .A(n657), .B(n467), .C(n103), .Y(n321) );
  NAND2X1 U129 ( .A(\mem<25><3> ), .B(n125), .Y(n103) );
  OAI21X1 U130 ( .A(n655), .B(n467), .C(n104), .Y(n322) );
  NAND2X1 U131 ( .A(\mem<25><4> ), .B(n125), .Y(n104) );
  OAI21X1 U134 ( .A(n663), .B(n465), .C(n107), .Y(n323) );
  NAND2X1 U135 ( .A(\mem<24><0> ), .B(n118), .Y(n107) );
  OAI21X1 U136 ( .A(n661), .B(n465), .C(n109), .Y(n324) );
  NAND2X1 U137 ( .A(\mem<24><1> ), .B(n118), .Y(n109) );
  OAI21X1 U138 ( .A(n659), .B(n465), .C(n110), .Y(n325) );
  NAND2X1 U139 ( .A(\mem<24><2> ), .B(n118), .Y(n110) );
  OAI21X1 U140 ( .A(n657), .B(n465), .C(n111), .Y(n326) );
  NAND2X1 U141 ( .A(\mem<24><3> ), .B(n118), .Y(n111) );
  OAI21X1 U142 ( .A(n655), .B(n465), .C(n112), .Y(n327) );
  NAND2X1 U143 ( .A(\mem<24><4> ), .B(n118), .Y(n112) );
  NAND3X1 U146 ( .A(N13), .B(n115), .C(N14), .Y(n114) );
  OAI21X1 U147 ( .A(n663), .B(n464), .C(n117), .Y(n328) );
  NAND2X1 U148 ( .A(\mem<23><0> ), .B(n108), .Y(n117) );
  OAI21X1 U149 ( .A(n661), .B(n464), .C(n119), .Y(n329) );
  NAND2X1 U150 ( .A(\mem<23><1> ), .B(n108), .Y(n119) );
  OAI21X1 U151 ( .A(n659), .B(n464), .C(n120), .Y(n330) );
  NAND2X1 U152 ( .A(\mem<23><2> ), .B(n108), .Y(n120) );
  OAI21X1 U153 ( .A(n657), .B(n464), .C(n121), .Y(n331) );
  NAND2X1 U154 ( .A(\mem<23><3> ), .B(n108), .Y(n121) );
  OAI21X1 U155 ( .A(n655), .B(n464), .C(n122), .Y(n332) );
  NAND2X1 U156 ( .A(\mem<23><4> ), .B(n108), .Y(n122) );
  OAI21X1 U159 ( .A(n663), .B(n462), .C(n124), .Y(n333) );
  NAND2X1 U160 ( .A(\mem<22><0> ), .B(n100), .Y(n124) );
  OAI21X1 U161 ( .A(n661), .B(n462), .C(n126), .Y(n334) );
  NAND2X1 U162 ( .A(\mem<22><1> ), .B(n100), .Y(n126) );
  OAI21X1 U163 ( .A(n659), .B(n462), .C(n127), .Y(n335) );
  NAND2X1 U164 ( .A(\mem<22><2> ), .B(n100), .Y(n127) );
  OAI21X1 U165 ( .A(n657), .B(n462), .C(n128), .Y(n336) );
  NAND2X1 U166 ( .A(\mem<22><3> ), .B(n100), .Y(n128) );
  OAI21X1 U167 ( .A(n655), .B(n462), .C(n129), .Y(n337) );
  NAND2X1 U168 ( .A(\mem<22><4> ), .B(n100), .Y(n129) );
  OAI21X1 U171 ( .A(n663), .B(n460), .C(n131), .Y(n338) );
  NAND2X1 U172 ( .A(\mem<21><0> ), .B(n92), .Y(n131) );
  OAI21X1 U173 ( .A(n661), .B(n460), .C(n133), .Y(n339) );
  NAND2X1 U174 ( .A(\mem<21><1> ), .B(n92), .Y(n133) );
  OAI21X1 U175 ( .A(n659), .B(n460), .C(n134), .Y(n340) );
  NAND2X1 U176 ( .A(\mem<21><2> ), .B(n92), .Y(n134) );
  OAI21X1 U177 ( .A(n657), .B(n460), .C(n135), .Y(n341) );
  NAND2X1 U178 ( .A(\mem<21><3> ), .B(n92), .Y(n135) );
  OAI21X1 U179 ( .A(n655), .B(n460), .C(n136), .Y(n342) );
  NAND2X1 U180 ( .A(\mem<21><4> ), .B(n92), .Y(n136) );
  OAI21X1 U183 ( .A(n663), .B(n458), .C(n138), .Y(n343) );
  NAND2X1 U184 ( .A(\mem<20><0> ), .B(n84), .Y(n138) );
  OAI21X1 U185 ( .A(n661), .B(n458), .C(n140), .Y(n344) );
  NAND2X1 U186 ( .A(\mem<20><1> ), .B(n84), .Y(n140) );
  OAI21X1 U187 ( .A(n659), .B(n458), .C(n141), .Y(n345) );
  NAND2X1 U188 ( .A(\mem<20><2> ), .B(n84), .Y(n141) );
  OAI21X1 U189 ( .A(n657), .B(n458), .C(n142), .Y(n346) );
  NAND2X1 U190 ( .A(\mem<20><3> ), .B(n84), .Y(n142) );
  OAI21X1 U191 ( .A(n655), .B(n458), .C(n143), .Y(n347) );
  NAND2X1 U192 ( .A(\mem<20><4> ), .B(n84), .Y(n143) );
  OAI21X1 U195 ( .A(n663), .B(n456), .C(n145), .Y(n348) );
  NAND2X1 U196 ( .A(\mem<19><0> ), .B(n76), .Y(n145) );
  OAI21X1 U197 ( .A(n661), .B(n456), .C(n147), .Y(n349) );
  NAND2X1 U198 ( .A(\mem<19><1> ), .B(n76), .Y(n147) );
  OAI21X1 U199 ( .A(n659), .B(n456), .C(n148), .Y(n350) );
  NAND2X1 U200 ( .A(\mem<19><2> ), .B(n76), .Y(n148) );
  OAI21X1 U201 ( .A(n657), .B(n456), .C(n149), .Y(n351) );
  NAND2X1 U202 ( .A(\mem<19><3> ), .B(n76), .Y(n149) );
  OAI21X1 U203 ( .A(n655), .B(n456), .C(n150), .Y(n352) );
  NAND2X1 U204 ( .A(\mem<19><4> ), .B(n76), .Y(n150) );
  OAI21X1 U207 ( .A(n664), .B(n454), .C(n152), .Y(n353) );
  NAND2X1 U208 ( .A(\mem<18><0> ), .B(n68), .Y(n152) );
  OAI21X1 U209 ( .A(n662), .B(n454), .C(n154), .Y(n354) );
  NAND2X1 U210 ( .A(\mem<18><1> ), .B(n68), .Y(n154) );
  OAI21X1 U211 ( .A(n660), .B(n454), .C(n155), .Y(n355) );
  NAND2X1 U212 ( .A(\mem<18><2> ), .B(n68), .Y(n155) );
  OAI21X1 U213 ( .A(n658), .B(n454), .C(n156), .Y(n356) );
  NAND2X1 U214 ( .A(\mem<18><3> ), .B(n68), .Y(n156) );
  OAI21X1 U215 ( .A(n656), .B(n454), .C(n157), .Y(n357) );
  NAND2X1 U216 ( .A(\mem<18><4> ), .B(n68), .Y(n157) );
  OAI21X1 U219 ( .A(n664), .B(n452), .C(n159), .Y(n358) );
  NAND2X1 U220 ( .A(\mem<17><0> ), .B(n60), .Y(n159) );
  OAI21X1 U221 ( .A(n662), .B(n452), .C(n161), .Y(n359) );
  NAND2X1 U222 ( .A(\mem<17><1> ), .B(n60), .Y(n161) );
  OAI21X1 U223 ( .A(n660), .B(n452), .C(n162), .Y(n360) );
  NAND2X1 U224 ( .A(\mem<17><2> ), .B(n60), .Y(n162) );
  OAI21X1 U225 ( .A(n658), .B(n452), .C(n163), .Y(n361) );
  NAND2X1 U226 ( .A(\mem<17><3> ), .B(n60), .Y(n163) );
  OAI21X1 U227 ( .A(n656), .B(n452), .C(n164), .Y(n362) );
  NAND2X1 U228 ( .A(\mem<17><4> ), .B(n60), .Y(n164) );
  OAI21X1 U231 ( .A(n664), .B(n450), .C(n166), .Y(n363) );
  NAND2X1 U232 ( .A(\mem<16><0> ), .B(n54), .Y(n166) );
  OAI21X1 U233 ( .A(n662), .B(n450), .C(n168), .Y(n364) );
  NAND2X1 U234 ( .A(\mem<16><1> ), .B(n54), .Y(n168) );
  OAI21X1 U235 ( .A(n660), .B(n450), .C(n169), .Y(n365) );
  NAND2X1 U236 ( .A(\mem<16><2> ), .B(n54), .Y(n169) );
  OAI21X1 U237 ( .A(n658), .B(n450), .C(n170), .Y(n366) );
  NAND2X1 U238 ( .A(\mem<16><3> ), .B(n54), .Y(n170) );
  OAI21X1 U239 ( .A(n656), .B(n450), .C(n171), .Y(n367) );
  NAND2X1 U240 ( .A(\mem<16><4> ), .B(n54), .Y(n171) );
  NAND3X1 U243 ( .A(n115), .B(n669), .C(N14), .Y(n172) );
  OAI21X1 U244 ( .A(n664), .B(n448), .C(n174), .Y(n368) );
  NAND2X1 U245 ( .A(\mem<15><0> ), .B(n50), .Y(n174) );
  OAI21X1 U246 ( .A(n662), .B(n448), .C(n176), .Y(n369) );
  NAND2X1 U247 ( .A(\mem<15><1> ), .B(n50), .Y(n176) );
  OAI21X1 U248 ( .A(n660), .B(n448), .C(n177), .Y(n370) );
  NAND2X1 U249 ( .A(\mem<15><2> ), .B(n50), .Y(n177) );
  OAI21X1 U250 ( .A(n658), .B(n448), .C(n178), .Y(n371) );
  NAND2X1 U251 ( .A(\mem<15><3> ), .B(n50), .Y(n178) );
  OAI21X1 U252 ( .A(n656), .B(n448), .C(n179), .Y(n372) );
  NAND2X1 U253 ( .A(\mem<15><4> ), .B(n50), .Y(n179) );
  OAI21X1 U256 ( .A(n664), .B(n281), .C(n181), .Y(n373) );
  NAND2X1 U257 ( .A(\mem<14><0> ), .B(n47), .Y(n181) );
  OAI21X1 U258 ( .A(n662), .B(n281), .C(n183), .Y(n374) );
  NAND2X1 U259 ( .A(\mem<14><1> ), .B(n47), .Y(n183) );
  OAI21X1 U260 ( .A(n660), .B(n281), .C(n184), .Y(n375) );
  NAND2X1 U261 ( .A(\mem<14><2> ), .B(n47), .Y(n184) );
  OAI21X1 U262 ( .A(n658), .B(n281), .C(n185), .Y(n376) );
  NAND2X1 U263 ( .A(\mem<14><3> ), .B(n47), .Y(n185) );
  OAI21X1 U264 ( .A(n656), .B(n281), .C(n186), .Y(n377) );
  NAND2X1 U265 ( .A(\mem<14><4> ), .B(n47), .Y(n186) );
  OAI21X1 U268 ( .A(n664), .B(n274), .C(n188), .Y(n378) );
  NAND2X1 U269 ( .A(\mem<13><0> ), .B(n44), .Y(n188) );
  OAI21X1 U270 ( .A(n662), .B(n274), .C(n190), .Y(n379) );
  NAND2X1 U271 ( .A(\mem<13><1> ), .B(n44), .Y(n190) );
  OAI21X1 U272 ( .A(n660), .B(n274), .C(n191), .Y(n380) );
  NAND2X1 U273 ( .A(\mem<13><2> ), .B(n44), .Y(n191) );
  OAI21X1 U274 ( .A(n658), .B(n274), .C(n192), .Y(n381) );
  NAND2X1 U275 ( .A(\mem<13><3> ), .B(n44), .Y(n192) );
  OAI21X1 U276 ( .A(n656), .B(n274), .C(n193), .Y(n382) );
  NAND2X1 U277 ( .A(\mem<13><4> ), .B(n44), .Y(n193) );
  OAI21X1 U280 ( .A(n664), .B(n267), .C(n195), .Y(n383) );
  NAND2X1 U281 ( .A(\mem<12><0> ), .B(n42), .Y(n195) );
  OAI21X1 U282 ( .A(n662), .B(n267), .C(n197), .Y(n384) );
  NAND2X1 U283 ( .A(\mem<12><1> ), .B(n42), .Y(n197) );
  OAI21X1 U284 ( .A(n660), .B(n267), .C(n198), .Y(n385) );
  NAND2X1 U285 ( .A(\mem<12><2> ), .B(n42), .Y(n198) );
  OAI21X1 U286 ( .A(n658), .B(n267), .C(n199), .Y(n386) );
  NAND2X1 U287 ( .A(\mem<12><3> ), .B(n42), .Y(n199) );
  OAI21X1 U288 ( .A(n656), .B(n267), .C(n200), .Y(n387) );
  NAND2X1 U289 ( .A(\mem<12><4> ), .B(n42), .Y(n200) );
  OAI21X1 U292 ( .A(n664), .B(n260), .C(n202), .Y(n388) );
  NAND2X1 U293 ( .A(\mem<11><0> ), .B(n40), .Y(n202) );
  OAI21X1 U294 ( .A(n662), .B(n260), .C(n204), .Y(n389) );
  NAND2X1 U295 ( .A(\mem<11><1> ), .B(n40), .Y(n204) );
  OAI21X1 U296 ( .A(n660), .B(n260), .C(n205), .Y(n390) );
  NAND2X1 U297 ( .A(\mem<11><2> ), .B(n40), .Y(n205) );
  OAI21X1 U298 ( .A(n658), .B(n260), .C(n206), .Y(n391) );
  NAND2X1 U299 ( .A(\mem<11><3> ), .B(n40), .Y(n206) );
  OAI21X1 U300 ( .A(n656), .B(n260), .C(n207), .Y(n392) );
  NAND2X1 U301 ( .A(\mem<11><4> ), .B(n40), .Y(n207) );
  OAI21X1 U304 ( .A(n664), .B(n253), .C(n209), .Y(n393) );
  NAND2X1 U305 ( .A(\mem<10><0> ), .B(n38), .Y(n209) );
  OAI21X1 U306 ( .A(n662), .B(n253), .C(n211), .Y(n394) );
  NAND2X1 U307 ( .A(\mem<10><1> ), .B(n38), .Y(n211) );
  OAI21X1 U308 ( .A(n660), .B(n253), .C(n212), .Y(n395) );
  NAND2X1 U309 ( .A(\mem<10><2> ), .B(n38), .Y(n212) );
  OAI21X1 U310 ( .A(n658), .B(n253), .C(n213), .Y(n396) );
  NAND2X1 U311 ( .A(\mem<10><3> ), .B(n38), .Y(n213) );
  OAI21X1 U312 ( .A(n656), .B(n253), .C(n214), .Y(n397) );
  NAND2X1 U313 ( .A(\mem<10><4> ), .B(n38), .Y(n214) );
  OAI21X1 U316 ( .A(n664), .B(n246), .C(n216), .Y(n398) );
  NAND2X1 U317 ( .A(\mem<9><0> ), .B(n36), .Y(n216) );
  OAI21X1 U318 ( .A(n662), .B(n246), .C(n218), .Y(n399) );
  NAND2X1 U319 ( .A(\mem<9><1> ), .B(n36), .Y(n218) );
  OAI21X1 U320 ( .A(n660), .B(n246), .C(n219), .Y(n400) );
  NAND2X1 U321 ( .A(\mem<9><2> ), .B(n36), .Y(n219) );
  OAI21X1 U322 ( .A(n658), .B(n246), .C(n220), .Y(n401) );
  NAND2X1 U323 ( .A(\mem<9><3> ), .B(n36), .Y(n220) );
  OAI21X1 U324 ( .A(n656), .B(n246), .C(n221), .Y(n402) );
  NAND2X1 U325 ( .A(\mem<9><4> ), .B(n36), .Y(n221) );
  OAI21X1 U328 ( .A(n664), .B(n239), .C(n223), .Y(n403) );
  NAND2X1 U329 ( .A(\mem<8><0> ), .B(n34), .Y(n223) );
  OAI21X1 U330 ( .A(n662), .B(n239), .C(n225), .Y(n404) );
  NAND2X1 U331 ( .A(\mem<8><1> ), .B(n34), .Y(n225) );
  OAI21X1 U332 ( .A(n660), .B(n239), .C(n226), .Y(n405) );
  NAND2X1 U333 ( .A(\mem<8><2> ), .B(n34), .Y(n226) );
  OAI21X1 U334 ( .A(n658), .B(n239), .C(n227), .Y(n406) );
  NAND2X1 U335 ( .A(\mem<8><3> ), .B(n34), .Y(n227) );
  OAI21X1 U336 ( .A(n656), .B(n239), .C(n228), .Y(n407) );
  NAND2X1 U337 ( .A(\mem<8><4> ), .B(n34), .Y(n228) );
  NAND3X1 U340 ( .A(n115), .B(n670), .C(N13), .Y(n229) );
  OAI21X1 U341 ( .A(n664), .B(n232), .C(n231), .Y(n408) );
  NAND2X1 U342 ( .A(\mem<7><0> ), .B(n32), .Y(n231) );
  OAI21X1 U343 ( .A(n662), .B(n232), .C(n233), .Y(n409) );
  NAND2X1 U344 ( .A(\mem<7><1> ), .B(n32), .Y(n233) );
  OAI21X1 U345 ( .A(n660), .B(n232), .C(n234), .Y(n410) );
  NAND2X1 U346 ( .A(\mem<7><2> ), .B(n32), .Y(n234) );
  OAI21X1 U347 ( .A(n658), .B(n232), .C(n235), .Y(n411) );
  NAND2X1 U348 ( .A(\mem<7><3> ), .B(n32), .Y(n235) );
  OAI21X1 U349 ( .A(n656), .B(n232), .C(n236), .Y(n412) );
  NAND2X1 U350 ( .A(\mem<7><4> ), .B(n32), .Y(n236) );
  NOR3X1 U353 ( .A(n667), .B(n666), .C(n668), .Y(n57) );
  OAI21X1 U354 ( .A(n664), .B(n224), .C(n238), .Y(n413) );
  NAND2X1 U355 ( .A(\mem<6><0> ), .B(n30), .Y(n238) );
  OAI21X1 U356 ( .A(n662), .B(n224), .C(n240), .Y(n414) );
  NAND2X1 U357 ( .A(\mem<6><1> ), .B(n30), .Y(n240) );
  OAI21X1 U358 ( .A(n660), .B(n224), .C(n241), .Y(n415) );
  NAND2X1 U359 ( .A(\mem<6><2> ), .B(n30), .Y(n241) );
  OAI21X1 U360 ( .A(n658), .B(n224), .C(n242), .Y(n416) );
  NAND2X1 U361 ( .A(\mem<6><3> ), .B(n30), .Y(n242) );
  OAI21X1 U362 ( .A(n656), .B(n224), .C(n243), .Y(n417) );
  NAND2X1 U363 ( .A(\mem<6><4> ), .B(n30), .Y(n243) );
  NOR3X1 U366 ( .A(n667), .B(n654), .C(n668), .Y(n65) );
  OAI21X1 U367 ( .A(n663), .B(n217), .C(n245), .Y(n418) );
  NAND2X1 U368 ( .A(\mem<5><0> ), .B(n28), .Y(n245) );
  OAI21X1 U369 ( .A(n661), .B(n217), .C(n247), .Y(n419) );
  NAND2X1 U370 ( .A(\mem<5><1> ), .B(n28), .Y(n247) );
  OAI21X1 U371 ( .A(n659), .B(n217), .C(n248), .Y(n420) );
  NAND2X1 U372 ( .A(\mem<5><2> ), .B(n28), .Y(n248) );
  OAI21X1 U373 ( .A(n657), .B(n217), .C(n249), .Y(n421) );
  NAND2X1 U374 ( .A(\mem<5><3> ), .B(n28), .Y(n249) );
  OAI21X1 U375 ( .A(n655), .B(n217), .C(n250), .Y(n422) );
  NAND2X1 U376 ( .A(\mem<5><4> ), .B(n28), .Y(n250) );
  NOR3X1 U379 ( .A(n666), .B(n5), .C(n668), .Y(n73) );
  OAI21X1 U380 ( .A(n664), .B(n210), .C(n252), .Y(n423) );
  NAND2X1 U381 ( .A(\mem<4><0> ), .B(n26), .Y(n252) );
  OAI21X1 U382 ( .A(n662), .B(n210), .C(n254), .Y(n424) );
  NAND2X1 U383 ( .A(\mem<4><1> ), .B(n26), .Y(n254) );
  OAI21X1 U384 ( .A(n660), .B(n210), .C(n255), .Y(n425) );
  NAND2X1 U385 ( .A(\mem<4><2> ), .B(n26), .Y(n255) );
  OAI21X1 U386 ( .A(n658), .B(n210), .C(n256), .Y(n426) );
  NAND2X1 U387 ( .A(\mem<4><3> ), .B(n26), .Y(n256) );
  OAI21X1 U388 ( .A(n656), .B(n210), .C(n257), .Y(n427) );
  NAND2X1 U389 ( .A(\mem<4><4> ), .B(n26), .Y(n257) );
  NOR3X1 U392 ( .A(n654), .B(n5), .C(n668), .Y(n81) );
  OAI21X1 U393 ( .A(n663), .B(n203), .C(n259), .Y(n428) );
  NAND2X1 U394 ( .A(\mem<3><0> ), .B(n24), .Y(n259) );
  OAI21X1 U395 ( .A(n661), .B(n203), .C(n261), .Y(n429) );
  NAND2X1 U396 ( .A(\mem<3><1> ), .B(n24), .Y(n261) );
  OAI21X1 U397 ( .A(n659), .B(n203), .C(n262), .Y(n430) );
  NAND2X1 U398 ( .A(\mem<3><2> ), .B(n24), .Y(n262) );
  OAI21X1 U399 ( .A(n657), .B(n203), .C(n263), .Y(n431) );
  NAND2X1 U400 ( .A(\mem<3><3> ), .B(n24), .Y(n263) );
  OAI21X1 U401 ( .A(n655), .B(n203), .C(n264), .Y(n432) );
  NAND2X1 U402 ( .A(\mem<3><4> ), .B(n24), .Y(n264) );
  NOR3X1 U405 ( .A(n666), .B(N12), .C(n667), .Y(n89) );
  OAI21X1 U406 ( .A(n664), .B(n196), .C(n266), .Y(n433) );
  NAND2X1 U407 ( .A(\mem<2><0> ), .B(n22), .Y(n266) );
  OAI21X1 U408 ( .A(n662), .B(n196), .C(n268), .Y(n434) );
  NAND2X1 U409 ( .A(\mem<2><1> ), .B(n22), .Y(n268) );
  OAI21X1 U410 ( .A(n660), .B(n196), .C(n269), .Y(n435) );
  NAND2X1 U411 ( .A(\mem<2><2> ), .B(n22), .Y(n269) );
  OAI21X1 U412 ( .A(n658), .B(n196), .C(n270), .Y(n436) );
  NAND2X1 U413 ( .A(\mem<2><3> ), .B(n22), .Y(n270) );
  OAI21X1 U414 ( .A(n656), .B(n196), .C(n271), .Y(n437) );
  NAND2X1 U415 ( .A(\mem<2><4> ), .B(n22), .Y(n271) );
  NOR3X1 U418 ( .A(n654), .B(N12), .C(n667), .Y(n97) );
  OAI21X1 U419 ( .A(n663), .B(n189), .C(n273), .Y(n438) );
  NAND2X1 U420 ( .A(\mem<1><0> ), .B(n20), .Y(n273) );
  OAI21X1 U421 ( .A(n661), .B(n189), .C(n275), .Y(n439) );
  NAND2X1 U422 ( .A(\mem<1><1> ), .B(n20), .Y(n275) );
  OAI21X1 U423 ( .A(n659), .B(n189), .C(n276), .Y(n440) );
  NAND2X1 U424 ( .A(\mem<1><2> ), .B(n20), .Y(n276) );
  OAI21X1 U425 ( .A(n657), .B(n189), .C(n277), .Y(n441) );
  NAND2X1 U426 ( .A(\mem<1><3> ), .B(n20), .Y(n277) );
  OAI21X1 U427 ( .A(n655), .B(n189), .C(n278), .Y(n442) );
  NAND2X1 U428 ( .A(\mem<1><4> ), .B(n20), .Y(n278) );
  NOR3X1 U431 ( .A(n5), .B(N12), .C(n666), .Y(n105) );
  OAI21X1 U432 ( .A(n664), .B(n182), .C(n280), .Y(n443) );
  NAND2X1 U433 ( .A(\mem<0><0> ), .B(n18), .Y(n280) );
  OAI21X1 U435 ( .A(n662), .B(n182), .C(n282), .Y(n444) );
  NAND2X1 U436 ( .A(\mem<0><1> ), .B(n18), .Y(n282) );
  OAI21X1 U438 ( .A(n660), .B(n182), .C(n283), .Y(n445) );
  NAND2X1 U439 ( .A(\mem<0><2> ), .B(n18), .Y(n283) );
  OAI21X1 U441 ( .A(n658), .B(n182), .C(n284), .Y(n446) );
  NAND2X1 U442 ( .A(\mem<0><3> ), .B(n18), .Y(n284) );
  OAI21X1 U444 ( .A(n656), .B(n182), .C(n285), .Y(n447) );
  NAND2X1 U445 ( .A(\mem<0><4> ), .B(n18), .Y(n285) );
  NOR3X1 U448 ( .A(n5), .B(N12), .C(n654), .Y(n113) );
  NAND3X1 U449 ( .A(n669), .B(n670), .C(n115), .Y(n286) );
  NOR3X1 U450 ( .A(\addr<5> ), .B(\addr<7> ), .C(\addr<6> ), .Y(n115) );
  MUX2X1 U2 ( .B(n597), .A(n598), .S(N13), .Y(n596) );
  INVX2 U3 ( .A(n6), .Y(n671) );
  MUX2X1 U4 ( .B(n613), .A(n612), .S(n634), .Y(n611) );
  MUX2X1 U5 ( .B(n622), .A(n621), .S(n639), .Y(n620) );
  MUX2X1 U6 ( .B(n583), .A(n582), .S(n634), .Y(n581) );
  MUX2X1 U7 ( .B(n625), .A(n624), .S(n639), .Y(n623) );
  INVX1 U8 ( .A(n645), .Y(n1) );
  MUX2X1 U9 ( .B(n523), .A(n522), .S(n634), .Y(n521) );
  AND2X1 U10 ( .A(n653), .B(n665), .Y(n56) );
  INVX1 U11 ( .A(n12), .Y(n656) );
  INVX1 U12 ( .A(n12), .Y(n655) );
  INVX1 U13 ( .A(n13), .Y(n658) );
  INVX1 U14 ( .A(n13), .Y(n657) );
  INVX1 U15 ( .A(n14), .Y(n660) );
  INVX1 U16 ( .A(n14), .Y(n659) );
  INVX1 U17 ( .A(n15), .Y(n662) );
  INVX1 U18 ( .A(n15), .Y(n661) );
  INVX1 U19 ( .A(n16), .Y(n664) );
  INVX1 U20 ( .A(n16), .Y(n663) );
  INVX1 U21 ( .A(N14), .Y(n670) );
  INVX1 U22 ( .A(rst), .Y(n665) );
  INVX1 U23 ( .A(N12), .Y(n668) );
  INVX1 U24 ( .A(N13), .Y(n669) );
  MUX2X1 U25 ( .B(n628), .A(n627), .S(n634), .Y(n626) );
  MUX2X1 U26 ( .B(n599), .A(n602), .S(n636), .Y(n613) );
  INVX1 U27 ( .A(n3), .Y(n2) );
  MUX2X1 U28 ( .B(\mem<1><4> ), .A(\mem<0><4> ), .S(n2), .Y(n624) );
  INVX1 U29 ( .A(n645), .Y(n3) );
  INVX1 U30 ( .A(n3), .Y(n4) );
  INVX1 U31 ( .A(n639), .Y(n5) );
  INVX1 U32 ( .A(n5), .Y(n667) );
  INVX4 U33 ( .A(n644), .Y(n650) );
  MUX2X1 U34 ( .B(\mem<11><3> ), .A(\mem<10><3> ), .S(n4), .Y(n589) );
  OR2X2 U35 ( .A(write), .B(rst), .Y(n6) );
  MUX2X1 U36 ( .B(n521), .A(n536), .S(n670), .Y(n630) );
  MUX2X1 U37 ( .B(n499), .A(n498), .S(n639), .Y(n497) );
  INVX8 U38 ( .A(n639), .Y(n640) );
  MUX2X1 U39 ( .B(n568), .A(n567), .S(n634), .Y(n566) );
  INVX1 U40 ( .A(n633), .Y(N17) );
  INVX1 U41 ( .A(n6), .Y(n7) );
  BUFX2 U42 ( .A(n286), .Y(n8) );
  INVX1 U43 ( .A(n8), .Y(n672) );
  BUFX2 U44 ( .A(n229), .Y(n9) );
  INVX1 U45 ( .A(n9), .Y(n673) );
  BUFX2 U46 ( .A(n172), .Y(n10) );
  INVX1 U47 ( .A(n10), .Y(n674) );
  BUFX2 U48 ( .A(n114), .Y(n11) );
  INVX1 U49 ( .A(n11), .Y(n675) );
  AND2X1 U60 ( .A(\data_in<4> ), .B(n56), .Y(n12) );
  AND2X1 U61 ( .A(\data_in<3> ), .B(n56), .Y(n13) );
  AND2X1 U72 ( .A(\data_in<2> ), .B(n56), .Y(n14) );
  AND2X1 U73 ( .A(\data_in<1> ), .B(n56), .Y(n15) );
  AND2X1 U84 ( .A(\data_in<0> ), .B(n56), .Y(n16) );
  AND2X1 U85 ( .A(n180), .B(n56), .Y(n17) );
  INVX1 U96 ( .A(n17), .Y(n18) );
  AND2X1 U97 ( .A(n187), .B(n56), .Y(n19) );
  INVX1 U108 ( .A(n19), .Y(n20) );
  AND2X1 U109 ( .A(n194), .B(n56), .Y(n21) );
  INVX1 U120 ( .A(n21), .Y(n22) );
  AND2X1 U121 ( .A(n201), .B(n56), .Y(n23) );
  INVX1 U132 ( .A(n23), .Y(n24) );
  AND2X1 U133 ( .A(n208), .B(n56), .Y(n25) );
  INVX1 U144 ( .A(n25), .Y(n26) );
  AND2X1 U145 ( .A(n215), .B(n56), .Y(n27) );
  INVX1 U157 ( .A(n27), .Y(n28) );
  AND2X1 U158 ( .A(n222), .B(n56), .Y(n29) );
  INVX1 U169 ( .A(n29), .Y(n30) );
  AND2X1 U170 ( .A(n230), .B(n56), .Y(n31) );
  INVX1 U181 ( .A(n31), .Y(n32) );
  AND2X1 U182 ( .A(n237), .B(n56), .Y(n33) );
  INVX1 U193 ( .A(n33), .Y(n34) );
  AND2X1 U194 ( .A(n244), .B(n56), .Y(n35) );
  INVX1 U205 ( .A(n35), .Y(n36) );
  AND2X1 U206 ( .A(n251), .B(n56), .Y(n37) );
  INVX1 U217 ( .A(n37), .Y(n38) );
  AND2X1 U218 ( .A(n258), .B(n56), .Y(n39) );
  INVX1 U229 ( .A(n39), .Y(n40) );
  AND2X1 U230 ( .A(n265), .B(n56), .Y(n41) );
  INVX1 U241 ( .A(n41), .Y(n42) );
  AND2X1 U242 ( .A(n272), .B(n56), .Y(n43) );
  INVX1 U254 ( .A(n43), .Y(n44) );
  AND2X1 U255 ( .A(n279), .B(n56), .Y(n45) );
  INVX1 U266 ( .A(n45), .Y(n47) );
  AND2X1 U267 ( .A(n287), .B(n56), .Y(n48) );
  INVX1 U278 ( .A(n48), .Y(n50) );
  AND2X1 U279 ( .A(n449), .B(n56), .Y(n52) );
  INVX1 U290 ( .A(n52), .Y(n54) );
  AND2X1 U291 ( .A(n451), .B(n56), .Y(n58) );
  INVX1 U302 ( .A(n58), .Y(n60) );
  AND2X1 U303 ( .A(n453), .B(n56), .Y(n66) );
  INVX1 U314 ( .A(n66), .Y(n68) );
  AND2X1 U315 ( .A(n455), .B(n56), .Y(n74) );
  INVX1 U326 ( .A(n74), .Y(n76) );
  AND2X1 U327 ( .A(n457), .B(n56), .Y(n82) );
  INVX1 U338 ( .A(n82), .Y(n84) );
  AND2X1 U339 ( .A(n459), .B(n56), .Y(n90) );
  INVX1 U351 ( .A(n90), .Y(n92) );
  AND2X1 U352 ( .A(n461), .B(n56), .Y(n98) );
  INVX1 U364 ( .A(n98), .Y(n100) );
  AND2X1 U365 ( .A(n463), .B(n56), .Y(n106) );
  INVX1 U377 ( .A(n106), .Y(n108) );
  AND2X1 U378 ( .A(n466), .B(n56), .Y(n116) );
  INVX1 U390 ( .A(n116), .Y(n118) );
  AND2X1 U391 ( .A(n468), .B(n56), .Y(n123) );
  INVX1 U403 ( .A(n123), .Y(n125) );
  AND2X1 U404 ( .A(n470), .B(n56), .Y(n130) );
  INVX1 U416 ( .A(n130), .Y(n132) );
  AND2X1 U417 ( .A(n472), .B(n56), .Y(n137) );
  INVX1 U429 ( .A(n137), .Y(n139) );
  AND2X1 U430 ( .A(n474), .B(n56), .Y(n144) );
  INVX1 U434 ( .A(n144), .Y(n146) );
  AND2X1 U437 ( .A(n476), .B(n56), .Y(n151) );
  INVX1 U440 ( .A(n151), .Y(n153) );
  AND2X1 U443 ( .A(n478), .B(n56), .Y(n158) );
  INVX1 U446 ( .A(n158), .Y(n160) );
  AND2X1 U447 ( .A(n175), .B(n56), .Y(n165) );
  INVX1 U451 ( .A(n165), .Y(n167) );
  INVX1 U452 ( .A(n175), .Y(n173) );
  AND2X1 U453 ( .A(n57), .B(n675), .Y(n175) );
  AND2X1 U454 ( .A(n672), .B(n113), .Y(n180) );
  INVX1 U455 ( .A(n180), .Y(n182) );
  AND2X1 U456 ( .A(n672), .B(n105), .Y(n187) );
  INVX1 U457 ( .A(n187), .Y(n189) );
  AND2X1 U458 ( .A(n672), .B(n97), .Y(n194) );
  INVX1 U459 ( .A(n194), .Y(n196) );
  AND2X1 U460 ( .A(n672), .B(n89), .Y(n201) );
  INVX1 U461 ( .A(n201), .Y(n203) );
  AND2X1 U462 ( .A(n672), .B(n81), .Y(n208) );
  INVX1 U463 ( .A(n208), .Y(n210) );
  AND2X1 U464 ( .A(n672), .B(n73), .Y(n215) );
  INVX1 U465 ( .A(n215), .Y(n217) );
  AND2X1 U466 ( .A(n672), .B(n65), .Y(n222) );
  INVX1 U467 ( .A(n222), .Y(n224) );
  AND2X1 U468 ( .A(n672), .B(n57), .Y(n230) );
  INVX1 U469 ( .A(n230), .Y(n232) );
  AND2X1 U470 ( .A(n673), .B(n113), .Y(n237) );
  INVX1 U471 ( .A(n237), .Y(n239) );
  AND2X1 U472 ( .A(n673), .B(n105), .Y(n244) );
  INVX1 U473 ( .A(n244), .Y(n246) );
  AND2X1 U474 ( .A(n673), .B(n97), .Y(n251) );
  INVX1 U475 ( .A(n251), .Y(n253) );
  AND2X1 U476 ( .A(n673), .B(n89), .Y(n258) );
  INVX1 U477 ( .A(n258), .Y(n260) );
  AND2X1 U478 ( .A(n673), .B(n81), .Y(n265) );
  INVX1 U479 ( .A(n265), .Y(n267) );
  AND2X1 U480 ( .A(n673), .B(n73), .Y(n272) );
  INVX1 U481 ( .A(n272), .Y(n274) );
  AND2X1 U482 ( .A(n673), .B(n65), .Y(n279) );
  INVX1 U483 ( .A(n279), .Y(n281) );
  AND2X1 U484 ( .A(n673), .B(n57), .Y(n287) );
  INVX1 U485 ( .A(n287), .Y(n448) );
  AND2X1 U486 ( .A(n674), .B(n113), .Y(n449) );
  INVX1 U487 ( .A(n449), .Y(n450) );
  AND2X1 U488 ( .A(n674), .B(n105), .Y(n451) );
  INVX1 U489 ( .A(n451), .Y(n452) );
  AND2X1 U490 ( .A(n674), .B(n97), .Y(n453) );
  INVX1 U491 ( .A(n453), .Y(n454) );
  AND2X1 U492 ( .A(n674), .B(n89), .Y(n455) );
  INVX1 U493 ( .A(n455), .Y(n456) );
  AND2X1 U494 ( .A(n674), .B(n81), .Y(n457) );
  INVX1 U495 ( .A(n457), .Y(n458) );
  AND2X1 U496 ( .A(n674), .B(n73), .Y(n459) );
  INVX1 U497 ( .A(n459), .Y(n460) );
  AND2X1 U498 ( .A(n674), .B(n65), .Y(n461) );
  INVX1 U499 ( .A(n461), .Y(n462) );
  AND2X1 U500 ( .A(n674), .B(n57), .Y(n463) );
  INVX1 U501 ( .A(n463), .Y(n464) );
  INVX1 U502 ( .A(n466), .Y(n465) );
  AND2X1 U503 ( .A(n113), .B(n675), .Y(n466) );
  INVX1 U504 ( .A(n468), .Y(n467) );
  AND2X1 U505 ( .A(n105), .B(n675), .Y(n468) );
  INVX1 U506 ( .A(n470), .Y(n469) );
  AND2X1 U507 ( .A(n97), .B(n675), .Y(n470) );
  INVX1 U508 ( .A(n472), .Y(n471) );
  AND2X1 U509 ( .A(n89), .B(n675), .Y(n472) );
  INVX1 U510 ( .A(n474), .Y(n473) );
  AND2X1 U511 ( .A(n81), .B(n675), .Y(n474) );
  INVX1 U512 ( .A(n476), .Y(n475) );
  AND2X1 U513 ( .A(n73), .B(n675), .Y(n476) );
  INVX1 U514 ( .A(n478), .Y(n477) );
  AND2X1 U515 ( .A(n65), .B(n675), .Y(n478) );
  MUX2X1 U516 ( .B(n480), .A(n481), .S(n651), .Y(n479) );
  MUX2X1 U517 ( .B(n483), .A(n484), .S(n643), .Y(n482) );
  MUX2X1 U518 ( .B(n486), .A(n487), .S(n651), .Y(n485) );
  MUX2X1 U519 ( .B(n489), .A(n490), .S(n643), .Y(n488) );
  MUX2X1 U520 ( .B(n492), .A(n493), .S(n635), .Y(n491) );
  MUX2X1 U521 ( .B(n495), .A(n496), .S(n643), .Y(n494) );
  MUX2X1 U522 ( .B(n501), .A(n502), .S(n643), .Y(n500) );
  MUX2X1 U523 ( .B(n504), .A(n505), .S(n643), .Y(n503) );
  MUX2X1 U524 ( .B(n507), .A(n508), .S(n635), .Y(n506) );
  MUX2X1 U525 ( .B(n510), .A(n511), .S(n643), .Y(n509) );
  MUX2X1 U526 ( .B(n513), .A(n514), .S(n643), .Y(n512) );
  MUX2X1 U527 ( .B(n516), .A(n517), .S(n651), .Y(n515) );
  MUX2X1 U528 ( .B(n519), .A(n520), .S(n643), .Y(n518) );
  MUX2X1 U529 ( .B(n525), .A(n526), .S(n640), .Y(n524) );
  MUX2X1 U530 ( .B(n528), .A(n529), .S(n640), .Y(n527) );
  MUX2X1 U531 ( .B(n531), .A(n532), .S(n641), .Y(n530) );
  MUX2X1 U532 ( .B(n534), .A(n535), .S(n641), .Y(n533) );
  MUX2X1 U533 ( .B(n537), .A(n538), .S(n635), .Y(n536) );
  MUX2X1 U534 ( .B(n540), .A(n541), .S(n640), .Y(n539) );
  MUX2X1 U535 ( .B(n543), .A(n544), .S(n641), .Y(n542) );
  MUX2X1 U536 ( .B(n546), .A(n547), .S(n640), .Y(n545) );
  MUX2X1 U537 ( .B(n549), .A(n550), .S(n640), .Y(n548) );
  MUX2X1 U538 ( .B(n552), .A(n553), .S(n635), .Y(n551) );
  MUX2X1 U539 ( .B(n555), .A(n556), .S(n641), .Y(n554) );
  MUX2X1 U540 ( .B(n558), .A(n559), .S(n640), .Y(n557) );
  MUX2X1 U541 ( .B(n561), .A(n562), .S(n640), .Y(n560) );
  MUX2X1 U542 ( .B(n564), .A(n565), .S(n642), .Y(n563) );
  MUX2X1 U543 ( .B(n570), .A(n571), .S(n640), .Y(n569) );
  MUX2X1 U544 ( .B(n573), .A(n574), .S(n642), .Y(n572) );
  MUX2X1 U545 ( .B(n576), .A(n577), .S(n641), .Y(n575) );
  MUX2X1 U546 ( .B(n579), .A(n580), .S(n641), .Y(n578) );
  MUX2X1 U547 ( .B(n585), .A(n586), .S(n642), .Y(n584) );
  MUX2X1 U548 ( .B(n588), .A(n589), .S(n642), .Y(n587) );
  MUX2X1 U549 ( .B(n591), .A(n592), .S(n640), .Y(n590) );
  MUX2X1 U550 ( .B(n594), .A(n595), .S(n642), .Y(n593) );
  MUX2X1 U551 ( .B(n600), .A(n601), .S(n641), .Y(n599) );
  MUX2X1 U552 ( .B(n603), .A(n604), .S(n641), .Y(n602) );
  MUX2X1 U553 ( .B(n606), .A(n607), .S(n641), .Y(n605) );
  MUX2X1 U554 ( .B(n609), .A(n610), .S(n640), .Y(n608) );
  MUX2X1 U555 ( .B(n615), .A(n616), .S(n640), .Y(n614) );
  MUX2X1 U556 ( .B(n618), .A(n619), .S(n642), .Y(n617) );
  MUX2X1 U557 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n647), .Y(n481) );
  MUX2X1 U558 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n1), .Y(n480) );
  MUX2X1 U559 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n647), .Y(n484) );
  MUX2X1 U560 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n647), .Y(n483) );
  MUX2X1 U561 ( .B(n482), .A(n479), .S(n638), .Y(n493) );
  MUX2X1 U562 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n1), .Y(n487) );
  MUX2X1 U563 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n1), .Y(n486) );
  MUX2X1 U564 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n647), .Y(n490) );
  MUX2X1 U565 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n647), .Y(n489) );
  MUX2X1 U566 ( .B(n488), .A(n485), .S(n637), .Y(n492) );
  MUX2X1 U567 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n648), .Y(n496) );
  MUX2X1 U568 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n647), .Y(n495) );
  MUX2X1 U569 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n650), .Y(n499) );
  MUX2X1 U570 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n652), .Y(n498) );
  MUX2X1 U571 ( .B(n497), .A(n494), .S(n637), .Y(n508) );
  MUX2X1 U572 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n646), .Y(n502) );
  MUX2X1 U573 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n646), .Y(n501) );
  MUX2X1 U574 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n650), .Y(n505) );
  MUX2X1 U575 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n648), .Y(n504) );
  MUX2X1 U576 ( .B(n503), .A(n500), .S(n637), .Y(n507) );
  MUX2X1 U577 ( .B(n506), .A(n491), .S(N14), .Y(n629) );
  MUX2X1 U578 ( .B(\mem<30><1> ), .A(\mem<31><1> ), .S(n649), .Y(n511) );
  MUX2X1 U579 ( .B(\mem<28><1> ), .A(\mem<29><1> ), .S(n648), .Y(n510) );
  MUX2X1 U580 ( .B(\mem<26><1> ), .A(\mem<27><1> ), .S(n649), .Y(n514) );
  MUX2X1 U581 ( .B(\mem<24><1> ), .A(\mem<25><1> ), .S(n649), .Y(n513) );
  MUX2X1 U582 ( .B(n512), .A(n509), .S(n638), .Y(n523) );
  MUX2X1 U583 ( .B(\mem<22><1> ), .A(\mem<23><1> ), .S(n649), .Y(n517) );
  MUX2X1 U584 ( .B(\mem<20><1> ), .A(\mem<21><1> ), .S(n649), .Y(n516) );
  MUX2X1 U585 ( .B(\mem<18><1> ), .A(\mem<19><1> ), .S(n646), .Y(n520) );
  MUX2X1 U586 ( .B(\mem<16><1> ), .A(\mem<17><1> ), .S(n646), .Y(n519) );
  MUX2X1 U587 ( .B(n518), .A(n515), .S(n638), .Y(n522) );
  MUX2X1 U588 ( .B(\mem<14><1> ), .A(\mem<15><1> ), .S(n649), .Y(n526) );
  MUX2X1 U589 ( .B(\mem<12><1> ), .A(\mem<13><1> ), .S(n649), .Y(n525) );
  MUX2X1 U590 ( .B(\mem<10><1> ), .A(\mem<11><1> ), .S(n646), .Y(n529) );
  MUX2X1 U591 ( .B(\mem<8><1> ), .A(\mem<9><1> ), .S(n646), .Y(n528) );
  MUX2X1 U592 ( .B(n527), .A(n524), .S(n638), .Y(n538) );
  MUX2X1 U593 ( .B(\mem<6><1> ), .A(\mem<7><1> ), .S(n646), .Y(n532) );
  MUX2X1 U594 ( .B(\mem<4><1> ), .A(\mem<5><1> ), .S(n648), .Y(n531) );
  MUX2X1 U595 ( .B(\mem<2><1> ), .A(\mem<3><1> ), .S(n648), .Y(n535) );
  MUX2X1 U596 ( .B(\mem<0><1> ), .A(\mem<1><1> ), .S(n646), .Y(n534) );
  MUX2X1 U597 ( .B(n533), .A(n530), .S(n638), .Y(n537) );
  MUX2X1 U598 ( .B(\mem<30><2> ), .A(\mem<31><2> ), .S(n646), .Y(n541) );
  MUX2X1 U599 ( .B(\mem<28><2> ), .A(\mem<29><2> ), .S(n646), .Y(n540) );
  MUX2X1 U600 ( .B(\mem<26><2> ), .A(\mem<27><2> ), .S(n646), .Y(n544) );
  MUX2X1 U601 ( .B(\mem<24><2> ), .A(\mem<25><2> ), .S(n649), .Y(n543) );
  MUX2X1 U602 ( .B(n542), .A(n539), .S(n638), .Y(n553) );
  MUX2X1 U603 ( .B(\mem<22><2> ), .A(\mem<23><2> ), .S(n648), .Y(n547) );
  MUX2X1 U604 ( .B(\mem<20><2> ), .A(\mem<21><2> ), .S(n649), .Y(n546) );
  MUX2X1 U605 ( .B(\mem<18><2> ), .A(\mem<19><2> ), .S(n646), .Y(n550) );
  MUX2X1 U606 ( .B(\mem<16><2> ), .A(\mem<17><2> ), .S(n649), .Y(n549) );
  MUX2X1 U607 ( .B(n548), .A(n545), .S(n637), .Y(n552) );
  MUX2X1 U608 ( .B(\mem<14><2> ), .A(\mem<15><2> ), .S(n649), .Y(n556) );
  MUX2X1 U609 ( .B(\mem<12><2> ), .A(\mem<13><2> ), .S(n646), .Y(n555) );
  MUX2X1 U610 ( .B(\mem<10><2> ), .A(\mem<11><2> ), .S(n648), .Y(n559) );
  MUX2X1 U611 ( .B(\mem<8><2> ), .A(\mem<9><2> ), .S(n649), .Y(n558) );
  MUX2X1 U612 ( .B(n557), .A(n554), .S(n637), .Y(n568) );
  MUX2X1 U613 ( .B(\mem<6><2> ), .A(\mem<7><2> ), .S(n649), .Y(n562) );
  MUX2X1 U614 ( .B(\mem<4><2> ), .A(\mem<5><2> ), .S(n646), .Y(n561) );
  MUX2X1 U615 ( .B(\mem<2><2> ), .A(\mem<3><2> ), .S(n648), .Y(n565) );
  MUX2X1 U616 ( .B(\mem<0><2> ), .A(\mem<1><2> ), .S(n648), .Y(n564) );
  MUX2X1 U617 ( .B(n563), .A(n560), .S(n638), .Y(n567) );
  MUX2X1 U618 ( .B(n566), .A(n551), .S(N14), .Y(n631) );
  MUX2X1 U619 ( .B(\mem<30><3> ), .A(\mem<31><3> ), .S(n647), .Y(n571) );
  MUX2X1 U620 ( .B(\mem<28><3> ), .A(\mem<29><3> ), .S(n647), .Y(n570) );
  MUX2X1 U621 ( .B(\mem<26><3> ), .A(\mem<27><3> ), .S(n648), .Y(n574) );
  MUX2X1 U622 ( .B(\mem<24><3> ), .A(\mem<25><3> ), .S(n646), .Y(n573) );
  MUX2X1 U623 ( .B(n572), .A(n569), .S(n637), .Y(n583) );
  MUX2X1 U624 ( .B(\mem<22><3> ), .A(\mem<23><3> ), .S(n649), .Y(n577) );
  MUX2X1 U625 ( .B(\mem<20><3> ), .A(\mem<21><3> ), .S(n647), .Y(n576) );
  MUX2X1 U626 ( .B(\mem<18><3> ), .A(\mem<19><3> ), .S(n648), .Y(n580) );
  MUX2X1 U627 ( .B(\mem<16><3> ), .A(\mem<17><3> ), .S(n647), .Y(n579) );
  MUX2X1 U628 ( .B(n578), .A(n575), .S(n638), .Y(n582) );
  MUX2X1 U629 ( .B(\mem<14><3> ), .A(\mem<15><3> ), .S(n648), .Y(n586) );
  MUX2X1 U630 ( .B(\mem<12><3> ), .A(\mem<13><3> ), .S(n647), .Y(n585) );
  MUX2X1 U631 ( .B(\mem<8><3> ), .A(\mem<9><3> ), .S(n652), .Y(n588) );
  MUX2X1 U632 ( .B(n587), .A(n584), .S(n638), .Y(n598) );
  MUX2X1 U633 ( .B(\mem<6><3> ), .A(\mem<7><3> ), .S(n650), .Y(n592) );
  MUX2X1 U634 ( .B(\mem<4><3> ), .A(\mem<5><3> ), .S(n648), .Y(n591) );
  MUX2X1 U635 ( .B(\mem<2><3> ), .A(\mem<3><3> ), .S(n652), .Y(n595) );
  MUX2X1 U636 ( .B(\mem<0><3> ), .A(\mem<1><3> ), .S(n652), .Y(n594) );
  MUX2X1 U637 ( .B(n593), .A(n590), .S(n638), .Y(n597) );
  MUX2X1 U638 ( .B(n596), .A(n581), .S(N14), .Y(n632) );
  MUX2X1 U639 ( .B(\mem<30><4> ), .A(\mem<31><4> ), .S(n649), .Y(n601) );
  MUX2X1 U640 ( .B(\mem<28><4> ), .A(\mem<29><4> ), .S(n647), .Y(n600) );
  MUX2X1 U641 ( .B(\mem<26><4> ), .A(\mem<27><4> ), .S(n647), .Y(n604) );
  MUX2X1 U642 ( .B(\mem<24><4> ), .A(\mem<25><4> ), .S(n647), .Y(n603) );
  MUX2X1 U643 ( .B(\mem<22><4> ), .A(\mem<23><4> ), .S(n646), .Y(n607) );
  MUX2X1 U644 ( .B(\mem<20><4> ), .A(\mem<21><4> ), .S(n649), .Y(n606) );
  MUX2X1 U645 ( .B(\mem<18><4> ), .A(\mem<19><4> ), .S(n647), .Y(n610) );
  MUX2X1 U646 ( .B(\mem<16><4> ), .A(\mem<17><4> ), .S(n648), .Y(n609) );
  MUX2X1 U647 ( .B(n608), .A(n605), .S(n637), .Y(n612) );
  MUX2X1 U648 ( .B(\mem<14><4> ), .A(\mem<15><4> ), .S(n649), .Y(n616) );
  MUX2X1 U649 ( .B(\mem<12><4> ), .A(\mem<13><4> ), .S(n646), .Y(n615) );
  MUX2X1 U650 ( .B(\mem<10><4> ), .A(\mem<11><4> ), .S(n650), .Y(n619) );
  MUX2X1 U651 ( .B(\mem<8><4> ), .A(\mem<9><4> ), .S(n650), .Y(n618) );
  MUX2X1 U652 ( .B(n617), .A(n614), .S(n637), .Y(n628) );
  MUX2X1 U653 ( .B(\mem<6><4> ), .A(\mem<7><4> ), .S(n649), .Y(n622) );
  MUX2X1 U654 ( .B(\mem<4><4> ), .A(\mem<5><4> ), .S(n647), .Y(n621) );
  MUX2X1 U655 ( .B(\mem<2><4> ), .A(\mem<3><4> ), .S(n650), .Y(n625) );
  MUX2X1 U656 ( .B(n623), .A(n620), .S(n637), .Y(n627) );
  MUX2X1 U657 ( .B(n626), .A(n611), .S(N14), .Y(n633) );
  INVX8 U658 ( .A(N13), .Y(n634) );
  INVX8 U659 ( .A(n634), .Y(n635) );
  INVX8 U660 ( .A(N12), .Y(n636) );
  INVX8 U661 ( .A(n636), .Y(n637) );
  INVX8 U662 ( .A(n636), .Y(n638) );
  INVX8 U663 ( .A(N11), .Y(n639) );
  INVX8 U664 ( .A(n639), .Y(n641) );
  INVX8 U665 ( .A(n639), .Y(n642) );
  INVX8 U666 ( .A(n639), .Y(n643) );
  INVX8 U667 ( .A(N10), .Y(n645) );
  INVX8 U668 ( .A(n644), .Y(n646) );
  INVX8 U669 ( .A(n645), .Y(n647) );
  INVX8 U670 ( .A(n645), .Y(n648) );
  INVX8 U671 ( .A(n645), .Y(n649) );
  INVX1 U672 ( .A(n631), .Y(N19) );
  INVX1 U673 ( .A(n629), .Y(N21) );
  INVX1 U674 ( .A(n630), .Y(N20) );
  INVX4 U675 ( .A(N10), .Y(n644) );
  INVX1 U676 ( .A(n632), .Y(N18) );
  INVX2 U677 ( .A(n639), .Y(n651) );
  BUFX2 U678 ( .A(N10), .Y(n652) );
  BUFX2 U679 ( .A(write), .Y(n653) );
  INVX1 U680 ( .A(n666), .Y(n654) );
  INVX1 U681 ( .A(n648), .Y(n666) );
  AND2X2 U682 ( .A(N21), .B(n7), .Y(\data_out<0> ) );
  AND2X2 U683 ( .A(N20), .B(n671), .Y(\data_out<1> ) );
  AND2X2 U684 ( .A(N19), .B(n671), .Y(\data_out<2> ) );
  AND2X2 U685 ( .A(N18), .B(n671), .Y(\data_out<3> ) );
  AND2X2 U686 ( .A(N17), .B(n7), .Y(\data_out<4> ) );
endmodule


module memc_Size1 ( .data_out(\data_out<0> ), .addr({\addr<7> , \addr<6> , 
        \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> }), 
    .data_in(\data_in<0> ), write, clk, rst, createdump, .file_id({
        \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> })
 );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , \data_in<0> , write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output \data_out<0> ;
  wire   N10, N11, N12, N13, N14, \mem<0><0> , \mem<1><0> , \mem<2><0> ,
         \mem<3><0> , \mem<4><0> , \mem<5><0> , \mem<6><0> , \mem<7><0> ,
         \mem<8><0> , \mem<9><0> , \mem<10><0> , \mem<11><0> , \mem<12><0> ,
         \mem<13><0> , \mem<14><0> , \mem<15><0> , \mem<16><0> , \mem<17><0> ,
         \mem<18><0> , \mem<19><0> , \mem<20><0> , \mem<21><0> , \mem<22><0> ,
         \mem<23><0> , \mem<24><0> , \mem<25><0> , \mem<26><0> , \mem<27><0> ,
         \mem<28><0> , \mem<29><0> , \mem<30><0> , \mem<31><0> , N17, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206;
  assign N10 = \addr<0> ;
  assign N11 = \addr<1> ;
  assign N12 = \addr<2> ;
  assign N13 = \addr<3> ;
  assign N14 = \addr<4> ;

  DFFPOSX1 \mem_reg<0><0>  ( .D(n92), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n91), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n90), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n89), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n88), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n87), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n86), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n85), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n84), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n83), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n82), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n81), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n80), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n79), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n78), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n77), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n76), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n75), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n74), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n73), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n72), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n71), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n70), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n69), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n68), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n67), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n66), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n65), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n64), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n63), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n62), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n61), .CLK(clk), .Q(\mem<31><0> ) );
  AND2X2 U2 ( .A(n2), .B(n57), .Y(\data_out<0> ) );
  INVX1 U3 ( .A(rst), .Y(n150) );
  INVX1 U4 ( .A(n154), .Y(n141) );
  INVX1 U5 ( .A(n140), .Y(N17) );
  INVX1 U6 ( .A(n97), .Y(n190) );
  INVX1 U7 ( .A(n98), .Y(n193) );
  INVX1 U8 ( .A(n99), .Y(n196) );
  INVX1 U9 ( .A(n100), .Y(n199) );
  INVX1 U10 ( .A(n101), .Y(n202) );
  BUFX2 U11 ( .A(write), .Y(n1) );
  INVX4 U12 ( .A(n109), .Y(n108) );
  AND2X2 U13 ( .A(\data_in<0> ), .B(n143), .Y(n94) );
  INVX2 U14 ( .A(n143), .Y(n205) );
  AND2X2 U15 ( .A(n103), .B(n94), .Y(n43) );
  AND2X2 U16 ( .A(n196), .B(n94), .Y(n49) );
  AND2X2 U17 ( .A(n105), .B(n94), .Y(n55) );
  AND2X2 U18 ( .A(\data_in<0> ), .B(n145), .Y(n93) );
  INVX2 U19 ( .A(n145), .Y(n186) );
  INVX1 U20 ( .A(write), .Y(n2) );
  OR2X2 U21 ( .A(\addr<5> ), .B(n59), .Y(n4) );
  INVX1 U22 ( .A(n4), .Y(n5) );
  AND2X2 U23 ( .A(n106), .B(n38), .Y(n6) );
  INVX1 U24 ( .A(n6), .Y(n7) );
  AND2X2 U25 ( .A(n103), .B(n38), .Y(n8) );
  INVX1 U26 ( .A(n8), .Y(n9) );
  AND2X2 U27 ( .A(n190), .B(n38), .Y(n10) );
  INVX1 U28 ( .A(n10), .Y(n11) );
  AND2X2 U29 ( .A(n193), .B(n38), .Y(n12) );
  INVX1 U30 ( .A(n12), .Y(n13) );
  AND2X2 U31 ( .A(n196), .B(n38), .Y(n14) );
  INVX1 U32 ( .A(n14), .Y(n15) );
  AND2X2 U33 ( .A(n199), .B(n38), .Y(n16) );
  INVX1 U34 ( .A(n16), .Y(n17) );
  AND2X2 U35 ( .A(n202), .B(n38), .Y(n18) );
  INVX1 U36 ( .A(n18), .Y(n19) );
  AND2X2 U37 ( .A(n105), .B(n38), .Y(n20) );
  INVX1 U38 ( .A(n20), .Y(n21) );
  AND2X2 U39 ( .A(n106), .B(n93), .Y(n22) );
  INVX1 U40 ( .A(n22), .Y(n23) );
  AND2X2 U41 ( .A(n103), .B(n93), .Y(n24) );
  INVX1 U42 ( .A(n24), .Y(n25) );
  AND2X2 U43 ( .A(n190), .B(n93), .Y(n26) );
  INVX1 U44 ( .A(n26), .Y(n27) );
  AND2X2 U45 ( .A(n193), .B(n93), .Y(n28) );
  INVX1 U46 ( .A(n28), .Y(n29) );
  AND2X2 U47 ( .A(n196), .B(n93), .Y(n30) );
  INVX1 U48 ( .A(n30), .Y(n31) );
  AND2X2 U49 ( .A(n199), .B(n93), .Y(n32) );
  INVX1 U50 ( .A(n32), .Y(n33) );
  AND2X2 U51 ( .A(n202), .B(n93), .Y(n34) );
  INVX1 U52 ( .A(n34), .Y(n35) );
  AND2X2 U53 ( .A(n105), .B(n93), .Y(n36) );
  INVX1 U54 ( .A(n36), .Y(n37) );
  INVX1 U55 ( .A(n154), .Y(n153) );
  INVX1 U56 ( .A(n156), .Y(n155) );
  INVX1 U57 ( .A(n152), .Y(n151) );
  AND2X2 U58 ( .A(\data_in<0> ), .B(n146), .Y(n38) );
  OR2X1 U59 ( .A(n153), .B(n155), .Y(n39) );
  INVX1 U60 ( .A(n39), .Y(n40) );
  AND2X2 U61 ( .A(n106), .B(n94), .Y(n41) );
  INVX1 U62 ( .A(n41), .Y(n42) );
  INVX1 U63 ( .A(n43), .Y(n44) );
  AND2X2 U64 ( .A(n190), .B(n94), .Y(n45) );
  INVX1 U65 ( .A(n45), .Y(n46) );
  AND2X2 U66 ( .A(n193), .B(n94), .Y(n47) );
  INVX1 U67 ( .A(n47), .Y(n48) );
  INVX1 U68 ( .A(n49), .Y(n50) );
  AND2X2 U69 ( .A(n199), .B(n94), .Y(n51) );
  INVX1 U70 ( .A(n51), .Y(n52) );
  AND2X2 U71 ( .A(n202), .B(n94), .Y(n53) );
  INVX1 U72 ( .A(n53), .Y(n54) );
  INVX1 U73 ( .A(n55), .Y(n56) );
  AND2X1 U74 ( .A(N17), .B(n150), .Y(n57) );
  INVX1 U75 ( .A(n160), .Y(n58) );
  INVX1 U76 ( .A(n58), .Y(n59) );
  AND2X1 U77 ( .A(n155), .B(n153), .Y(n60) );
  OR2X1 U78 ( .A(\addr<6> ), .B(\addr<7> ), .Y(n95) );
  INVX1 U79 ( .A(n95), .Y(n96) );
  BUFX2 U80 ( .A(n191), .Y(n97) );
  BUFX2 U81 ( .A(n194), .Y(n98) );
  BUFX2 U82 ( .A(n197), .Y(n99) );
  BUFX2 U83 ( .A(n200), .Y(n100) );
  BUFX2 U84 ( .A(n203), .Y(n101) );
  INVX1 U85 ( .A(n103), .Y(n102) );
  AND2X1 U86 ( .A(n152), .B(n60), .Y(n103) );
  INVX1 U87 ( .A(n105), .Y(n104) );
  AND2X2 U88 ( .A(n152), .B(n40), .Y(n105) );
  AND2X1 U89 ( .A(n151), .B(n60), .Y(n106) );
  INVX1 U90 ( .A(n106), .Y(n107) );
  AND2X1 U91 ( .A(\data_in<0> ), .B(n148), .Y(n109) );
  MUX2X1 U92 ( .B(n111), .A(n112), .S(n141), .Y(n110) );
  MUX2X1 U93 ( .B(n114), .A(n115), .S(n141), .Y(n113) );
  MUX2X1 U94 ( .B(n117), .A(n118), .S(n141), .Y(n116) );
  MUX2X1 U95 ( .B(n120), .A(n121), .S(n141), .Y(n119) );
  MUX2X1 U96 ( .B(n123), .A(n124), .S(n157), .Y(n122) );
  MUX2X1 U97 ( .B(n126), .A(n127), .S(n141), .Y(n125) );
  MUX2X1 U98 ( .B(n129), .A(n130), .S(n141), .Y(n128) );
  MUX2X1 U99 ( .B(n132), .A(n133), .S(n141), .Y(n131) );
  MUX2X1 U100 ( .B(n135), .A(n136), .S(n141), .Y(n134) );
  MUX2X1 U101 ( .B(n138), .A(n139), .S(n157), .Y(n137) );
  MUX2X1 U102 ( .B(\mem<30><0> ), .A(\mem<31><0> ), .S(n142), .Y(n112) );
  MUX2X1 U103 ( .B(\mem<28><0> ), .A(\mem<29><0> ), .S(n142), .Y(n111) );
  MUX2X1 U104 ( .B(\mem<26><0> ), .A(\mem<27><0> ), .S(n142), .Y(n115) );
  MUX2X1 U105 ( .B(\mem<24><0> ), .A(\mem<25><0> ), .S(n142), .Y(n114) );
  MUX2X1 U106 ( .B(n113), .A(n110), .S(n155), .Y(n124) );
  MUX2X1 U107 ( .B(\mem<22><0> ), .A(\mem<23><0> ), .S(n142), .Y(n118) );
  MUX2X1 U108 ( .B(\mem<20><0> ), .A(\mem<21><0> ), .S(n142), .Y(n117) );
  MUX2X1 U109 ( .B(\mem<18><0> ), .A(\mem<19><0> ), .S(n142), .Y(n121) );
  MUX2X1 U110 ( .B(\mem<16><0> ), .A(\mem<17><0> ), .S(n142), .Y(n120) );
  MUX2X1 U111 ( .B(n119), .A(n116), .S(n155), .Y(n123) );
  MUX2X1 U112 ( .B(\mem<14><0> ), .A(\mem<15><0> ), .S(n142), .Y(n127) );
  MUX2X1 U113 ( .B(\mem<12><0> ), .A(\mem<13><0> ), .S(n142), .Y(n126) );
  MUX2X1 U114 ( .B(\mem<10><0> ), .A(\mem<11><0> ), .S(n142), .Y(n130) );
  MUX2X1 U115 ( .B(\mem<8><0> ), .A(\mem<9><0> ), .S(n142), .Y(n129) );
  MUX2X1 U116 ( .B(n128), .A(n125), .S(n155), .Y(n139) );
  MUX2X1 U117 ( .B(\mem<6><0> ), .A(\mem<7><0> ), .S(n142), .Y(n133) );
  MUX2X1 U118 ( .B(\mem<4><0> ), .A(\mem<5><0> ), .S(n142), .Y(n132) );
  MUX2X1 U119 ( .B(\mem<2><0> ), .A(\mem<3><0> ), .S(n142), .Y(n136) );
  MUX2X1 U120 ( .B(\mem<0><0> ), .A(\mem<1><0> ), .S(n142), .Y(n135) );
  MUX2X1 U121 ( .B(n134), .A(n131), .S(n155), .Y(n138) );
  MUX2X1 U122 ( .B(n137), .A(n122), .S(N14), .Y(n140) );
  INVX8 U123 ( .A(n152), .Y(n142) );
  INVX1 U124 ( .A(N12), .Y(n156) );
  INVX1 U125 ( .A(n5), .Y(n144) );
  NOR3X1 U126 ( .A(N13), .B(n144), .C(N14), .Y(n143) );
  INVX1 U127 ( .A(N13), .Y(n158) );
  NOR3X1 U128 ( .A(n158), .B(n149), .C(N14), .Y(n145) );
  INVX1 U129 ( .A(N14), .Y(n159) );
  INVX1 U130 ( .A(n177), .Y(n146) );
  INVX1 U131 ( .A(n146), .Y(n147) );
  INVX1 U132 ( .A(N11), .Y(n154) );
  INVX1 U133 ( .A(N10), .Y(n152) );
  INVX1 U134 ( .A(n5), .Y(n149) );
  NOR3X1 U135 ( .A(n159), .B(n158), .C(n149), .Y(n148) );
  INVX2 U136 ( .A(n148), .Y(n168) );
  INVX1 U137 ( .A(n158), .Y(n157) );
  NAND3X1 U138 ( .A(n1), .B(n150), .C(n96), .Y(n160) );
  OAI21X1 U139 ( .A(n168), .B(n107), .C(\mem<31><0> ), .Y(n161) );
  OAI21X1 U140 ( .A(n108), .B(n107), .C(n161), .Y(n61) );
  OAI21X1 U141 ( .A(n102), .B(n168), .C(\mem<30><0> ), .Y(n162) );
  OAI21X1 U142 ( .A(n102), .B(n108), .C(n162), .Y(n62) );
  NAND3X1 U143 ( .A(n151), .B(n155), .C(n154), .Y(n191) );
  OAI21X1 U144 ( .A(n97), .B(n168), .C(\mem<29><0> ), .Y(n163) );
  OAI21X1 U145 ( .A(n97), .B(n108), .C(n163), .Y(n63) );
  NAND3X1 U146 ( .A(n155), .B(n154), .C(n152), .Y(n194) );
  OAI21X1 U147 ( .A(n98), .B(n168), .C(\mem<28><0> ), .Y(n164) );
  OAI21X1 U148 ( .A(n98), .B(n108), .C(n164), .Y(n64) );
  NAND3X1 U149 ( .A(n151), .B(n153), .C(n156), .Y(n197) );
  OAI21X1 U150 ( .A(n99), .B(n168), .C(\mem<27><0> ), .Y(n165) );
  OAI21X1 U151 ( .A(n99), .B(n108), .C(n165), .Y(n65) );
  NAND3X1 U152 ( .A(n156), .B(n153), .C(n152), .Y(n200) );
  OAI21X1 U153 ( .A(n100), .B(n168), .C(\mem<26><0> ), .Y(n166) );
  OAI21X1 U154 ( .A(n100), .B(n108), .C(n166), .Y(n66) );
  NAND3X1 U155 ( .A(n151), .B(n156), .C(n154), .Y(n203) );
  OAI21X1 U156 ( .A(n101), .B(n168), .C(\mem<25><0> ), .Y(n167) );
  OAI21X1 U157 ( .A(n101), .B(n108), .C(n167), .Y(n67) );
  OAI21X1 U158 ( .A(n104), .B(n168), .C(\mem<24><0> ), .Y(n169) );
  OAI21X1 U159 ( .A(n104), .B(n108), .C(n169), .Y(n68) );
  NAND3X1 U160 ( .A(N14), .B(n5), .C(n158), .Y(n177) );
  OAI21X1 U161 ( .A(n147), .B(n107), .C(\mem<23><0> ), .Y(n170) );
  NAND2X1 U162 ( .A(n7), .B(n170), .Y(n69) );
  OAI21X1 U163 ( .A(n147), .B(n102), .C(\mem<22><0> ), .Y(n171) );
  NAND2X1 U164 ( .A(n9), .B(n171), .Y(n70) );
  OAI21X1 U165 ( .A(n147), .B(n97), .C(\mem<21><0> ), .Y(n172) );
  NAND2X1 U166 ( .A(n11), .B(n172), .Y(n71) );
  OAI21X1 U167 ( .A(n147), .B(n98), .C(\mem<20><0> ), .Y(n173) );
  NAND2X1 U168 ( .A(n13), .B(n173), .Y(n72) );
  OAI21X1 U169 ( .A(n147), .B(n99), .C(\mem<19><0> ), .Y(n174) );
  NAND2X1 U170 ( .A(n15), .B(n174), .Y(n73) );
  OAI21X1 U171 ( .A(n147), .B(n100), .C(\mem<18><0> ), .Y(n175) );
  NAND2X1 U172 ( .A(n17), .B(n175), .Y(n74) );
  OAI21X1 U173 ( .A(n147), .B(n101), .C(\mem<17><0> ), .Y(n176) );
  NAND2X1 U174 ( .A(n19), .B(n176), .Y(n75) );
  OAI21X1 U175 ( .A(n147), .B(n104), .C(\mem<16><0> ), .Y(n178) );
  NAND2X1 U176 ( .A(n21), .B(n178), .Y(n76) );
  OAI21X1 U177 ( .A(n186), .B(n107), .C(\mem<15><0> ), .Y(n179) );
  NAND2X1 U178 ( .A(n23), .B(n179), .Y(n77) );
  OAI21X1 U179 ( .A(n186), .B(n102), .C(\mem<14><0> ), .Y(n180) );
  NAND2X1 U180 ( .A(n25), .B(n180), .Y(n78) );
  OAI21X1 U181 ( .A(n186), .B(n97), .C(\mem<13><0> ), .Y(n181) );
  NAND2X1 U182 ( .A(n27), .B(n181), .Y(n79) );
  OAI21X1 U183 ( .A(n186), .B(n98), .C(\mem<12><0> ), .Y(n182) );
  NAND2X1 U184 ( .A(n29), .B(n182), .Y(n80) );
  OAI21X1 U185 ( .A(n186), .B(n99), .C(\mem<11><0> ), .Y(n183) );
  NAND2X1 U186 ( .A(n31), .B(n183), .Y(n81) );
  OAI21X1 U187 ( .A(n186), .B(n100), .C(\mem<10><0> ), .Y(n184) );
  NAND2X1 U188 ( .A(n33), .B(n184), .Y(n82) );
  OAI21X1 U189 ( .A(n186), .B(n101), .C(\mem<9><0> ), .Y(n185) );
  NAND2X1 U190 ( .A(n35), .B(n185), .Y(n83) );
  OAI21X1 U191 ( .A(n186), .B(n104), .C(\mem<8><0> ), .Y(n187) );
  NAND2X1 U192 ( .A(n37), .B(n187), .Y(n84) );
  OAI21X1 U193 ( .A(n205), .B(n107), .C(\mem<7><0> ), .Y(n188) );
  NAND2X1 U194 ( .A(n42), .B(n188), .Y(n85) );
  OAI21X1 U195 ( .A(n205), .B(n102), .C(\mem<6><0> ), .Y(n189) );
  NAND2X1 U196 ( .A(n44), .B(n189), .Y(n86) );
  OAI21X1 U197 ( .A(n205), .B(n97), .C(\mem<5><0> ), .Y(n192) );
  NAND2X1 U198 ( .A(n46), .B(n192), .Y(n87) );
  OAI21X1 U199 ( .A(n205), .B(n98), .C(\mem<4><0> ), .Y(n195) );
  NAND2X1 U200 ( .A(n48), .B(n195), .Y(n88) );
  OAI21X1 U201 ( .A(n205), .B(n99), .C(\mem<3><0> ), .Y(n198) );
  NAND2X1 U202 ( .A(n50), .B(n198), .Y(n89) );
  OAI21X1 U203 ( .A(n205), .B(n100), .C(\mem<2><0> ), .Y(n201) );
  NAND2X1 U204 ( .A(n52), .B(n201), .Y(n90) );
  OAI21X1 U205 ( .A(n205), .B(n101), .C(\mem<1><0> ), .Y(n204) );
  NAND2X1 U206 ( .A(n54), .B(n204), .Y(n91) );
  OAI21X1 U207 ( .A(n205), .B(n104), .C(\mem<0><0> ), .Y(n206) );
  NAND2X1 U208 ( .A(n56), .B(n206), .Y(n92) );
endmodule


module memv ( data_out, .addr({\addr<7> , \addr<6> , \addr<5> , \addr<4> , 
        \addr<3> , \addr<2> , \addr<1> , \addr<0> }), data_in, write, clk, rst, 
        createdump, .file_id({\file_id<4> , \file_id<3> , \file_id<2> , 
        \file_id<1> , \file_id<0> }) );
  input \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> ,
         \addr<1> , \addr<0> , data_in, write, clk, rst, createdump,
         \file_id<4> , \file_id<3> , \file_id<2> , \file_id<1> , \file_id<0> ;
  output data_out;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \mem<0> , \mem<1> , \mem<2> ,
         \mem<3> , \mem<4> , \mem<5> , \mem<6> , \mem<7> , \mem<8> , \mem<9> ,
         \mem<10> , \mem<11> , \mem<12> , \mem<13> , \mem<14> , \mem<15> ,
         \mem<16> , \mem<17> , \mem<18> , \mem<19> , \mem<20> , \mem<21> ,
         \mem<22> , \mem<23> , \mem<24> , \mem<25> , \mem<26> , \mem<27> ,
         \mem<28> , \mem<29> , \mem<30> , \mem<31> , \mem<32> , \mem<33> ,
         \mem<34> , \mem<35> , \mem<36> , \mem<37> , \mem<38> , \mem<39> ,
         \mem<40> , \mem<41> , \mem<42> , \mem<43> , \mem<44> , \mem<45> ,
         \mem<46> , \mem<47> , \mem<48> , \mem<49> , \mem<50> , \mem<51> ,
         \mem<52> , \mem<53> , \mem<54> , \mem<55> , \mem<56> , \mem<57> ,
         \mem<58> , \mem<59> , \mem<60> , \mem<61> , \mem<62> , \mem<63> ,
         \mem<64> , \mem<65> , \mem<66> , \mem<67> , \mem<68> , \mem<69> ,
         \mem<70> , \mem<71> , \mem<72> , \mem<73> , \mem<74> , \mem<75> ,
         \mem<76> , \mem<77> , \mem<78> , \mem<79> , \mem<80> , \mem<81> ,
         \mem<82> , \mem<83> , \mem<84> , \mem<85> , \mem<86> , \mem<87> ,
         \mem<88> , \mem<89> , \mem<90> , \mem<91> , \mem<92> , \mem<93> ,
         \mem<94> , \mem<95> , \mem<96> , \mem<97> , \mem<98> , \mem<99> ,
         \mem<100> , \mem<101> , \mem<102> , \mem<103> , \mem<104> ,
         \mem<105> , \mem<106> , \mem<107> , \mem<108> , \mem<109> ,
         \mem<110> , \mem<111> , \mem<112> , \mem<113> , \mem<114> ,
         \mem<115> , \mem<116> , \mem<117> , \mem<118> , \mem<119> ,
         \mem<120> , \mem<121> , \mem<122> , \mem<123> , \mem<124> ,
         \mem<125> , \mem<126> , \mem<127> , \mem<128> , \mem<129> ,
         \mem<130> , \mem<131> , \mem<132> , \mem<133> , \mem<134> ,
         \mem<135> , \mem<136> , \mem<137> , \mem<138> , \mem<139> ,
         \mem<140> , \mem<141> , \mem<142> , \mem<143> , \mem<144> ,
         \mem<145> , \mem<146> , \mem<147> , \mem<148> , \mem<149> ,
         \mem<150> , \mem<151> , \mem<152> , \mem<153> , \mem<154> ,
         \mem<155> , \mem<156> , \mem<157> , \mem<158> , \mem<159> ,
         \mem<160> , \mem<161> , \mem<162> , \mem<163> , \mem<164> ,
         \mem<165> , \mem<166> , \mem<167> , \mem<168> , \mem<169> ,
         \mem<170> , \mem<171> , \mem<172> , \mem<173> , \mem<174> ,
         \mem<175> , \mem<176> , \mem<177> , \mem<178> , \mem<179> ,
         \mem<180> , \mem<181> , \mem<182> , \mem<183> , \mem<184> ,
         \mem<185> , \mem<186> , \mem<187> , \mem<188> , \mem<189> ,
         \mem<190> , \mem<191> , \mem<192> , \mem<193> , \mem<194> ,
         \mem<195> , \mem<196> , \mem<197> , \mem<198> , \mem<199> ,
         \mem<200> , \mem<201> , \mem<202> , \mem<203> , \mem<204> ,
         \mem<205> , \mem<206> , \mem<207> , \mem<208> , \mem<209> ,
         \mem<210> , \mem<211> , \mem<212> , \mem<213> , \mem<214> ,
         \mem<215> , \mem<216> , \mem<217> , \mem<218> , \mem<219> ,
         \mem<220> , \mem<221> , \mem<222> , \mem<223> , \mem<224> ,
         \mem<225> , \mem<226> , \mem<227> , \mem<228> , \mem<229> ,
         \mem<230> , \mem<231> , \mem<232> , \mem<233> , \mem<234> ,
         \mem<235> , \mem<236> , \mem<237> , \mem<238> , \mem<239> ,
         \mem<240> , \mem<241> , \mem<242> , \mem<243> , \mem<244> ,
         \mem<245> , \mem<246> , \mem<247> , \mem<248> , \mem<249> ,
         \mem<250> , \mem<251> , \mem<252> , \mem<253> , \mem<254> ,
         \mem<255> , N28, n42, n46, n49, n52, n55, n58, n61, n64, n67, n70,
         n73, n76, n79, n82, n85, n88, n90, n91, n92, n94, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n113, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n132, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n151, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n170, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n188, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n206, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n224,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n243, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n261, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n279, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n297, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n316, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n334, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n352, n355, n356, n357, n358, n359, n361, n363, n364, n365,
         n366, n367, n368, n370, n371, n372, n373, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n43, n44, n45, n47, n48, n50, n51, n53, n54, n56, n57, n59, n60, n62,
         n63, n65, n66, n68, n69, n71, n72, n74, n75, n77, n78, n80, n81, n83,
         n84, n86, n87, n89, n93, n95, n112, n114, n130, n131, n133, n149,
         n150, n152, n169, n171, n187, n189, n205, n207, n223, n225, n241,
         n242, n244, n260, n262, n278, n280, n296, n298, n314, n315, n317,
         n333, n335, n351, n353, n354, n360, n362, n369, n374, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999;
  assign N18 = \addr<0> ;
  assign N19 = \addr<1> ;
  assign N20 = \addr<2> ;
  assign N21 = \addr<3> ;
  assign N22 = \addr<4> ;
  assign N23 = \addr<5> ;
  assign N24 = \addr<6> ;
  assign N25 = \addr<7> ;

  DFFPOSX1 \mem_reg<0>  ( .D(n633), .CLK(clk), .Q(\mem<0> ) );
  DFFPOSX1 \mem_reg<1>  ( .D(n632), .CLK(clk), .Q(\mem<1> ) );
  DFFPOSX1 \mem_reg<2>  ( .D(n631), .CLK(clk), .Q(\mem<2> ) );
  DFFPOSX1 \mem_reg<3>  ( .D(n630), .CLK(clk), .Q(\mem<3> ) );
  DFFPOSX1 \mem_reg<4>  ( .D(n629), .CLK(clk), .Q(\mem<4> ) );
  DFFPOSX1 \mem_reg<5>  ( .D(n628), .CLK(clk), .Q(\mem<5> ) );
  DFFPOSX1 \mem_reg<6>  ( .D(n627), .CLK(clk), .Q(\mem<6> ) );
  DFFPOSX1 \mem_reg<7>  ( .D(n626), .CLK(clk), .Q(\mem<7> ) );
  DFFPOSX1 \mem_reg<8>  ( .D(n625), .CLK(clk), .Q(\mem<8> ) );
  DFFPOSX1 \mem_reg<9>  ( .D(n624), .CLK(clk), .Q(\mem<9> ) );
  DFFPOSX1 \mem_reg<10>  ( .D(n623), .CLK(clk), .Q(\mem<10> ) );
  DFFPOSX1 \mem_reg<11>  ( .D(n622), .CLK(clk), .Q(\mem<11> ) );
  DFFPOSX1 \mem_reg<12>  ( .D(n621), .CLK(clk), .Q(\mem<12> ) );
  DFFPOSX1 \mem_reg<13>  ( .D(n620), .CLK(clk), .Q(\mem<13> ) );
  DFFPOSX1 \mem_reg<14>  ( .D(n619), .CLK(clk), .Q(\mem<14> ) );
  DFFPOSX1 \mem_reg<15>  ( .D(n618), .CLK(clk), .Q(\mem<15> ) );
  DFFPOSX1 \mem_reg<16>  ( .D(n617), .CLK(clk), .Q(\mem<16> ) );
  DFFPOSX1 \mem_reg<17>  ( .D(n616), .CLK(clk), .Q(\mem<17> ) );
  DFFPOSX1 \mem_reg<18>  ( .D(n615), .CLK(clk), .Q(\mem<18> ) );
  DFFPOSX1 \mem_reg<19>  ( .D(n614), .CLK(clk), .Q(\mem<19> ) );
  DFFPOSX1 \mem_reg<20>  ( .D(n613), .CLK(clk), .Q(\mem<20> ) );
  DFFPOSX1 \mem_reg<21>  ( .D(n612), .CLK(clk), .Q(\mem<21> ) );
  DFFPOSX1 \mem_reg<22>  ( .D(n611), .CLK(clk), .Q(\mem<22> ) );
  DFFPOSX1 \mem_reg<23>  ( .D(n610), .CLK(clk), .Q(\mem<23> ) );
  DFFPOSX1 \mem_reg<24>  ( .D(n609), .CLK(clk), .Q(\mem<24> ) );
  DFFPOSX1 \mem_reg<25>  ( .D(n608), .CLK(clk), .Q(\mem<25> ) );
  DFFPOSX1 \mem_reg<26>  ( .D(n607), .CLK(clk), .Q(\mem<26> ) );
  DFFPOSX1 \mem_reg<27>  ( .D(n606), .CLK(clk), .Q(\mem<27> ) );
  DFFPOSX1 \mem_reg<28>  ( .D(n605), .CLK(clk), .Q(\mem<28> ) );
  DFFPOSX1 \mem_reg<29>  ( .D(n604), .CLK(clk), .Q(\mem<29> ) );
  DFFPOSX1 \mem_reg<30>  ( .D(n603), .CLK(clk), .Q(\mem<30> ) );
  DFFPOSX1 \mem_reg<31>  ( .D(n602), .CLK(clk), .Q(\mem<31> ) );
  DFFPOSX1 \mem_reg<32>  ( .D(n601), .CLK(clk), .Q(\mem<32> ) );
  DFFPOSX1 \mem_reg<33>  ( .D(n600), .CLK(clk), .Q(\mem<33> ) );
  DFFPOSX1 \mem_reg<34>  ( .D(n599), .CLK(clk), .Q(\mem<34> ) );
  DFFPOSX1 \mem_reg<35>  ( .D(n598), .CLK(clk), .Q(\mem<35> ) );
  DFFPOSX1 \mem_reg<36>  ( .D(n597), .CLK(clk), .Q(\mem<36> ) );
  DFFPOSX1 \mem_reg<37>  ( .D(n596), .CLK(clk), .Q(\mem<37> ) );
  DFFPOSX1 \mem_reg<38>  ( .D(n595), .CLK(clk), .Q(\mem<38> ) );
  DFFPOSX1 \mem_reg<39>  ( .D(n594), .CLK(clk), .Q(\mem<39> ) );
  DFFPOSX1 \mem_reg<40>  ( .D(n593), .CLK(clk), .Q(\mem<40> ) );
  DFFPOSX1 \mem_reg<41>  ( .D(n592), .CLK(clk), .Q(\mem<41> ) );
  DFFPOSX1 \mem_reg<42>  ( .D(n591), .CLK(clk), .Q(\mem<42> ) );
  DFFPOSX1 \mem_reg<43>  ( .D(n590), .CLK(clk), .Q(\mem<43> ) );
  DFFPOSX1 \mem_reg<44>  ( .D(n589), .CLK(clk), .Q(\mem<44> ) );
  DFFPOSX1 \mem_reg<45>  ( .D(n588), .CLK(clk), .Q(\mem<45> ) );
  DFFPOSX1 \mem_reg<46>  ( .D(n587), .CLK(clk), .Q(\mem<46> ) );
  DFFPOSX1 \mem_reg<47>  ( .D(n586), .CLK(clk), .Q(\mem<47> ) );
  DFFPOSX1 \mem_reg<48>  ( .D(n585), .CLK(clk), .Q(\mem<48> ) );
  DFFPOSX1 \mem_reg<49>  ( .D(n584), .CLK(clk), .Q(\mem<49> ) );
  DFFPOSX1 \mem_reg<50>  ( .D(n583), .CLK(clk), .Q(\mem<50> ) );
  DFFPOSX1 \mem_reg<51>  ( .D(n582), .CLK(clk), .Q(\mem<51> ) );
  DFFPOSX1 \mem_reg<52>  ( .D(n581), .CLK(clk), .Q(\mem<52> ) );
  DFFPOSX1 \mem_reg<53>  ( .D(n580), .CLK(clk), .Q(\mem<53> ) );
  DFFPOSX1 \mem_reg<54>  ( .D(n579), .CLK(clk), .Q(\mem<54> ) );
  DFFPOSX1 \mem_reg<55>  ( .D(n578), .CLK(clk), .Q(\mem<55> ) );
  DFFPOSX1 \mem_reg<56>  ( .D(n577), .CLK(clk), .Q(\mem<56> ) );
  DFFPOSX1 \mem_reg<57>  ( .D(n576), .CLK(clk), .Q(\mem<57> ) );
  DFFPOSX1 \mem_reg<58>  ( .D(n575), .CLK(clk), .Q(\mem<58> ) );
  DFFPOSX1 \mem_reg<59>  ( .D(n574), .CLK(clk), .Q(\mem<59> ) );
  DFFPOSX1 \mem_reg<60>  ( .D(n573), .CLK(clk), .Q(\mem<60> ) );
  DFFPOSX1 \mem_reg<61>  ( .D(n572), .CLK(clk), .Q(\mem<61> ) );
  DFFPOSX1 \mem_reg<62>  ( .D(n571), .CLK(clk), .Q(\mem<62> ) );
  DFFPOSX1 \mem_reg<63>  ( .D(n570), .CLK(clk), .Q(\mem<63> ) );
  DFFPOSX1 \mem_reg<64>  ( .D(n569), .CLK(clk), .Q(\mem<64> ) );
  DFFPOSX1 \mem_reg<65>  ( .D(n568), .CLK(clk), .Q(\mem<65> ) );
  DFFPOSX1 \mem_reg<66>  ( .D(n567), .CLK(clk), .Q(\mem<66> ) );
  DFFPOSX1 \mem_reg<67>  ( .D(n566), .CLK(clk), .Q(\mem<67> ) );
  DFFPOSX1 \mem_reg<68>  ( .D(n565), .CLK(clk), .Q(\mem<68> ) );
  DFFPOSX1 \mem_reg<69>  ( .D(n564), .CLK(clk), .Q(\mem<69> ) );
  DFFPOSX1 \mem_reg<70>  ( .D(n563), .CLK(clk), .Q(\mem<70> ) );
  DFFPOSX1 \mem_reg<71>  ( .D(n562), .CLK(clk), .Q(\mem<71> ) );
  DFFPOSX1 \mem_reg<72>  ( .D(n561), .CLK(clk), .Q(\mem<72> ) );
  DFFPOSX1 \mem_reg<73>  ( .D(n560), .CLK(clk), .Q(\mem<73> ) );
  DFFPOSX1 \mem_reg<74>  ( .D(n559), .CLK(clk), .Q(\mem<74> ) );
  DFFPOSX1 \mem_reg<75>  ( .D(n558), .CLK(clk), .Q(\mem<75> ) );
  DFFPOSX1 \mem_reg<76>  ( .D(n557), .CLK(clk), .Q(\mem<76> ) );
  DFFPOSX1 \mem_reg<77>  ( .D(n556), .CLK(clk), .Q(\mem<77> ) );
  DFFPOSX1 \mem_reg<78>  ( .D(n555), .CLK(clk), .Q(\mem<78> ) );
  DFFPOSX1 \mem_reg<79>  ( .D(n554), .CLK(clk), .Q(\mem<79> ) );
  DFFPOSX1 \mem_reg<80>  ( .D(n553), .CLK(clk), .Q(\mem<80> ) );
  DFFPOSX1 \mem_reg<81>  ( .D(n552), .CLK(clk), .Q(\mem<81> ) );
  DFFPOSX1 \mem_reg<82>  ( .D(n551), .CLK(clk), .Q(\mem<82> ) );
  DFFPOSX1 \mem_reg<83>  ( .D(n550), .CLK(clk), .Q(\mem<83> ) );
  DFFPOSX1 \mem_reg<84>  ( .D(n549), .CLK(clk), .Q(\mem<84> ) );
  DFFPOSX1 \mem_reg<85>  ( .D(n548), .CLK(clk), .Q(\mem<85> ) );
  DFFPOSX1 \mem_reg<86>  ( .D(n547), .CLK(clk), .Q(\mem<86> ) );
  DFFPOSX1 \mem_reg<87>  ( .D(n546), .CLK(clk), .Q(\mem<87> ) );
  DFFPOSX1 \mem_reg<88>  ( .D(n545), .CLK(clk), .Q(\mem<88> ) );
  DFFPOSX1 \mem_reg<89>  ( .D(n544), .CLK(clk), .Q(\mem<89> ) );
  DFFPOSX1 \mem_reg<90>  ( .D(n543), .CLK(clk), .Q(\mem<90> ) );
  DFFPOSX1 \mem_reg<91>  ( .D(n542), .CLK(clk), .Q(\mem<91> ) );
  DFFPOSX1 \mem_reg<92>  ( .D(n541), .CLK(clk), .Q(\mem<92> ) );
  DFFPOSX1 \mem_reg<93>  ( .D(n540), .CLK(clk), .Q(\mem<93> ) );
  DFFPOSX1 \mem_reg<94>  ( .D(n539), .CLK(clk), .Q(\mem<94> ) );
  DFFPOSX1 \mem_reg<95>  ( .D(n538), .CLK(clk), .Q(\mem<95> ) );
  DFFPOSX1 \mem_reg<96>  ( .D(n537), .CLK(clk), .Q(\mem<96> ) );
  DFFPOSX1 \mem_reg<97>  ( .D(n536), .CLK(clk), .Q(\mem<97> ) );
  DFFPOSX1 \mem_reg<98>  ( .D(n535), .CLK(clk), .Q(\mem<98> ) );
  DFFPOSX1 \mem_reg<99>  ( .D(n534), .CLK(clk), .Q(\mem<99> ) );
  DFFPOSX1 \mem_reg<100>  ( .D(n533), .CLK(clk), .Q(\mem<100> ) );
  DFFPOSX1 \mem_reg<101>  ( .D(n532), .CLK(clk), .Q(\mem<101> ) );
  DFFPOSX1 \mem_reg<102>  ( .D(n531), .CLK(clk), .Q(\mem<102> ) );
  DFFPOSX1 \mem_reg<103>  ( .D(n530), .CLK(clk), .Q(\mem<103> ) );
  DFFPOSX1 \mem_reg<104>  ( .D(n529), .CLK(clk), .Q(\mem<104> ) );
  DFFPOSX1 \mem_reg<105>  ( .D(n528), .CLK(clk), .Q(\mem<105> ) );
  DFFPOSX1 \mem_reg<106>  ( .D(n527), .CLK(clk), .Q(\mem<106> ) );
  DFFPOSX1 \mem_reg<107>  ( .D(n526), .CLK(clk), .Q(\mem<107> ) );
  DFFPOSX1 \mem_reg<108>  ( .D(n525), .CLK(clk), .Q(\mem<108> ) );
  DFFPOSX1 \mem_reg<109>  ( .D(n524), .CLK(clk), .Q(\mem<109> ) );
  DFFPOSX1 \mem_reg<110>  ( .D(n523), .CLK(clk), .Q(\mem<110> ) );
  DFFPOSX1 \mem_reg<111>  ( .D(n522), .CLK(clk), .Q(\mem<111> ) );
  DFFPOSX1 \mem_reg<112>  ( .D(n521), .CLK(clk), .Q(\mem<112> ) );
  DFFPOSX1 \mem_reg<113>  ( .D(n520), .CLK(clk), .Q(\mem<113> ) );
  DFFPOSX1 \mem_reg<114>  ( .D(n519), .CLK(clk), .Q(\mem<114> ) );
  DFFPOSX1 \mem_reg<115>  ( .D(n518), .CLK(clk), .Q(\mem<115> ) );
  DFFPOSX1 \mem_reg<116>  ( .D(n517), .CLK(clk), .Q(\mem<116> ) );
  DFFPOSX1 \mem_reg<117>  ( .D(n516), .CLK(clk), .Q(\mem<117> ) );
  DFFPOSX1 \mem_reg<118>  ( .D(n515), .CLK(clk), .Q(\mem<118> ) );
  DFFPOSX1 \mem_reg<119>  ( .D(n514), .CLK(clk), .Q(\mem<119> ) );
  DFFPOSX1 \mem_reg<120>  ( .D(n513), .CLK(clk), .Q(\mem<120> ) );
  DFFPOSX1 \mem_reg<121>  ( .D(n512), .CLK(clk), .Q(\mem<121> ) );
  DFFPOSX1 \mem_reg<122>  ( .D(n511), .CLK(clk), .Q(\mem<122> ) );
  DFFPOSX1 \mem_reg<123>  ( .D(n510), .CLK(clk), .Q(\mem<123> ) );
  DFFPOSX1 \mem_reg<124>  ( .D(n509), .CLK(clk), .Q(\mem<124> ) );
  DFFPOSX1 \mem_reg<125>  ( .D(n508), .CLK(clk), .Q(\mem<125> ) );
  DFFPOSX1 \mem_reg<126>  ( .D(n507), .CLK(clk), .Q(\mem<126> ) );
  DFFPOSX1 \mem_reg<127>  ( .D(n506), .CLK(clk), .Q(\mem<127> ) );
  DFFPOSX1 \mem_reg<128>  ( .D(n505), .CLK(clk), .Q(\mem<128> ) );
  DFFPOSX1 \mem_reg<129>  ( .D(n504), .CLK(clk), .Q(\mem<129> ) );
  DFFPOSX1 \mem_reg<130>  ( .D(n503), .CLK(clk), .Q(\mem<130> ) );
  DFFPOSX1 \mem_reg<131>  ( .D(n502), .CLK(clk), .Q(\mem<131> ) );
  DFFPOSX1 \mem_reg<132>  ( .D(n501), .CLK(clk), .Q(\mem<132> ) );
  DFFPOSX1 \mem_reg<133>  ( .D(n500), .CLK(clk), .Q(\mem<133> ) );
  DFFPOSX1 \mem_reg<134>  ( .D(n499), .CLK(clk), .Q(\mem<134> ) );
  DFFPOSX1 \mem_reg<135>  ( .D(n498), .CLK(clk), .Q(\mem<135> ) );
  DFFPOSX1 \mem_reg<136>  ( .D(n497), .CLK(clk), .Q(\mem<136> ) );
  DFFPOSX1 \mem_reg<137>  ( .D(n496), .CLK(clk), .Q(\mem<137> ) );
  DFFPOSX1 \mem_reg<138>  ( .D(n495), .CLK(clk), .Q(\mem<138> ) );
  DFFPOSX1 \mem_reg<139>  ( .D(n494), .CLK(clk), .Q(\mem<139> ) );
  DFFPOSX1 \mem_reg<140>  ( .D(n493), .CLK(clk), .Q(\mem<140> ) );
  DFFPOSX1 \mem_reg<141>  ( .D(n492), .CLK(clk), .Q(\mem<141> ) );
  DFFPOSX1 \mem_reg<142>  ( .D(n491), .CLK(clk), .Q(\mem<142> ) );
  DFFPOSX1 \mem_reg<143>  ( .D(n490), .CLK(clk), .Q(\mem<143> ) );
  DFFPOSX1 \mem_reg<144>  ( .D(n489), .CLK(clk), .Q(\mem<144> ) );
  DFFPOSX1 \mem_reg<145>  ( .D(n488), .CLK(clk), .Q(\mem<145> ) );
  DFFPOSX1 \mem_reg<146>  ( .D(n487), .CLK(clk), .Q(\mem<146> ) );
  DFFPOSX1 \mem_reg<147>  ( .D(n486), .CLK(clk), .Q(\mem<147> ) );
  DFFPOSX1 \mem_reg<148>  ( .D(n485), .CLK(clk), .Q(\mem<148> ) );
  DFFPOSX1 \mem_reg<149>  ( .D(n484), .CLK(clk), .Q(\mem<149> ) );
  DFFPOSX1 \mem_reg<150>  ( .D(n483), .CLK(clk), .Q(\mem<150> ) );
  DFFPOSX1 \mem_reg<151>  ( .D(n482), .CLK(clk), .Q(\mem<151> ) );
  DFFPOSX1 \mem_reg<152>  ( .D(n481), .CLK(clk), .Q(\mem<152> ) );
  DFFPOSX1 \mem_reg<153>  ( .D(n480), .CLK(clk), .Q(\mem<153> ) );
  DFFPOSX1 \mem_reg<154>  ( .D(n479), .CLK(clk), .Q(\mem<154> ) );
  DFFPOSX1 \mem_reg<155>  ( .D(n478), .CLK(clk), .Q(\mem<155> ) );
  DFFPOSX1 \mem_reg<156>  ( .D(n477), .CLK(clk), .Q(\mem<156> ) );
  DFFPOSX1 \mem_reg<157>  ( .D(n476), .CLK(clk), .Q(\mem<157> ) );
  DFFPOSX1 \mem_reg<158>  ( .D(n475), .CLK(clk), .Q(\mem<158> ) );
  DFFPOSX1 \mem_reg<159>  ( .D(n474), .CLK(clk), .Q(\mem<159> ) );
  DFFPOSX1 \mem_reg<160>  ( .D(n473), .CLK(clk), .Q(\mem<160> ) );
  DFFPOSX1 \mem_reg<161>  ( .D(n472), .CLK(clk), .Q(\mem<161> ) );
  DFFPOSX1 \mem_reg<162>  ( .D(n471), .CLK(clk), .Q(\mem<162> ) );
  DFFPOSX1 \mem_reg<163>  ( .D(n470), .CLK(clk), .Q(\mem<163> ) );
  DFFPOSX1 \mem_reg<164>  ( .D(n469), .CLK(clk), .Q(\mem<164> ) );
  DFFPOSX1 \mem_reg<165>  ( .D(n468), .CLK(clk), .Q(\mem<165> ) );
  DFFPOSX1 \mem_reg<166>  ( .D(n467), .CLK(clk), .Q(\mem<166> ) );
  DFFPOSX1 \mem_reg<167>  ( .D(n466), .CLK(clk), .Q(\mem<167> ) );
  DFFPOSX1 \mem_reg<168>  ( .D(n465), .CLK(clk), .Q(\mem<168> ) );
  DFFPOSX1 \mem_reg<169>  ( .D(n464), .CLK(clk), .Q(\mem<169> ) );
  DFFPOSX1 \mem_reg<170>  ( .D(n463), .CLK(clk), .Q(\mem<170> ) );
  DFFPOSX1 \mem_reg<171>  ( .D(n462), .CLK(clk), .Q(\mem<171> ) );
  DFFPOSX1 \mem_reg<172>  ( .D(n461), .CLK(clk), .Q(\mem<172> ) );
  DFFPOSX1 \mem_reg<173>  ( .D(n460), .CLK(clk), .Q(\mem<173> ) );
  DFFPOSX1 \mem_reg<174>  ( .D(n459), .CLK(clk), .Q(\mem<174> ) );
  DFFPOSX1 \mem_reg<175>  ( .D(n458), .CLK(clk), .Q(\mem<175> ) );
  DFFPOSX1 \mem_reg<176>  ( .D(n457), .CLK(clk), .Q(\mem<176> ) );
  DFFPOSX1 \mem_reg<177>  ( .D(n456), .CLK(clk), .Q(\mem<177> ) );
  DFFPOSX1 \mem_reg<178>  ( .D(n455), .CLK(clk), .Q(\mem<178> ) );
  DFFPOSX1 \mem_reg<179>  ( .D(n454), .CLK(clk), .Q(\mem<179> ) );
  DFFPOSX1 \mem_reg<180>  ( .D(n453), .CLK(clk), .Q(\mem<180> ) );
  DFFPOSX1 \mem_reg<181>  ( .D(n452), .CLK(clk), .Q(\mem<181> ) );
  DFFPOSX1 \mem_reg<182>  ( .D(n451), .CLK(clk), .Q(\mem<182> ) );
  DFFPOSX1 \mem_reg<183>  ( .D(n450), .CLK(clk), .Q(\mem<183> ) );
  DFFPOSX1 \mem_reg<184>  ( .D(n449), .CLK(clk), .Q(\mem<184> ) );
  DFFPOSX1 \mem_reg<185>  ( .D(n448), .CLK(clk), .Q(\mem<185> ) );
  DFFPOSX1 \mem_reg<186>  ( .D(n447), .CLK(clk), .Q(\mem<186> ) );
  DFFPOSX1 \mem_reg<187>  ( .D(n446), .CLK(clk), .Q(\mem<187> ) );
  DFFPOSX1 \mem_reg<188>  ( .D(n445), .CLK(clk), .Q(\mem<188> ) );
  DFFPOSX1 \mem_reg<189>  ( .D(n444), .CLK(clk), .Q(\mem<189> ) );
  DFFPOSX1 \mem_reg<190>  ( .D(n443), .CLK(clk), .Q(\mem<190> ) );
  DFFPOSX1 \mem_reg<191>  ( .D(n442), .CLK(clk), .Q(\mem<191> ) );
  DFFPOSX1 \mem_reg<192>  ( .D(n441), .CLK(clk), .Q(\mem<192> ) );
  DFFPOSX1 \mem_reg<193>  ( .D(n440), .CLK(clk), .Q(\mem<193> ) );
  DFFPOSX1 \mem_reg<194>  ( .D(n439), .CLK(clk), .Q(\mem<194> ) );
  DFFPOSX1 \mem_reg<195>  ( .D(n438), .CLK(clk), .Q(\mem<195> ) );
  DFFPOSX1 \mem_reg<196>  ( .D(n437), .CLK(clk), .Q(\mem<196> ) );
  DFFPOSX1 \mem_reg<197>  ( .D(n436), .CLK(clk), .Q(\mem<197> ) );
  DFFPOSX1 \mem_reg<198>  ( .D(n435), .CLK(clk), .Q(\mem<198> ) );
  DFFPOSX1 \mem_reg<199>  ( .D(n434), .CLK(clk), .Q(\mem<199> ) );
  DFFPOSX1 \mem_reg<200>  ( .D(n433), .CLK(clk), .Q(\mem<200> ) );
  DFFPOSX1 \mem_reg<201>  ( .D(n432), .CLK(clk), .Q(\mem<201> ) );
  DFFPOSX1 \mem_reg<202>  ( .D(n431), .CLK(clk), .Q(\mem<202> ) );
  DFFPOSX1 \mem_reg<203>  ( .D(n430), .CLK(clk), .Q(\mem<203> ) );
  DFFPOSX1 \mem_reg<204>  ( .D(n429), .CLK(clk), .Q(\mem<204> ) );
  DFFPOSX1 \mem_reg<205>  ( .D(n428), .CLK(clk), .Q(\mem<205> ) );
  DFFPOSX1 \mem_reg<206>  ( .D(n427), .CLK(clk), .Q(\mem<206> ) );
  DFFPOSX1 \mem_reg<207>  ( .D(n426), .CLK(clk), .Q(\mem<207> ) );
  DFFPOSX1 \mem_reg<208>  ( .D(n425), .CLK(clk), .Q(\mem<208> ) );
  DFFPOSX1 \mem_reg<209>  ( .D(n424), .CLK(clk), .Q(\mem<209> ) );
  DFFPOSX1 \mem_reg<210>  ( .D(n423), .CLK(clk), .Q(\mem<210> ) );
  DFFPOSX1 \mem_reg<211>  ( .D(n422), .CLK(clk), .Q(\mem<211> ) );
  DFFPOSX1 \mem_reg<212>  ( .D(n421), .CLK(clk), .Q(\mem<212> ) );
  DFFPOSX1 \mem_reg<213>  ( .D(n420), .CLK(clk), .Q(\mem<213> ) );
  DFFPOSX1 \mem_reg<214>  ( .D(n419), .CLK(clk), .Q(\mem<214> ) );
  DFFPOSX1 \mem_reg<215>  ( .D(n418), .CLK(clk), .Q(\mem<215> ) );
  DFFPOSX1 \mem_reg<216>  ( .D(n417), .CLK(clk), .Q(\mem<216> ) );
  DFFPOSX1 \mem_reg<217>  ( .D(n416), .CLK(clk), .Q(\mem<217> ) );
  DFFPOSX1 \mem_reg<218>  ( .D(n415), .CLK(clk), .Q(\mem<218> ) );
  DFFPOSX1 \mem_reg<219>  ( .D(n414), .CLK(clk), .Q(\mem<219> ) );
  DFFPOSX1 \mem_reg<220>  ( .D(n413), .CLK(clk), .Q(\mem<220> ) );
  DFFPOSX1 \mem_reg<221>  ( .D(n412), .CLK(clk), .Q(\mem<221> ) );
  DFFPOSX1 \mem_reg<222>  ( .D(n411), .CLK(clk), .Q(\mem<222> ) );
  DFFPOSX1 \mem_reg<223>  ( .D(n410), .CLK(clk), .Q(\mem<223> ) );
  DFFPOSX1 \mem_reg<224>  ( .D(n409), .CLK(clk), .Q(\mem<224> ) );
  DFFPOSX1 \mem_reg<225>  ( .D(n408), .CLK(clk), .Q(\mem<225> ) );
  DFFPOSX1 \mem_reg<226>  ( .D(n407), .CLK(clk), .Q(\mem<226> ) );
  DFFPOSX1 \mem_reg<227>  ( .D(n406), .CLK(clk), .Q(\mem<227> ) );
  DFFPOSX1 \mem_reg<228>  ( .D(n405), .CLK(clk), .Q(\mem<228> ) );
  DFFPOSX1 \mem_reg<229>  ( .D(n404), .CLK(clk), .Q(\mem<229> ) );
  DFFPOSX1 \mem_reg<230>  ( .D(n403), .CLK(clk), .Q(\mem<230> ) );
  DFFPOSX1 \mem_reg<231>  ( .D(n402), .CLK(clk), .Q(\mem<231> ) );
  DFFPOSX1 \mem_reg<232>  ( .D(n401), .CLK(clk), .Q(\mem<232> ) );
  DFFPOSX1 \mem_reg<233>  ( .D(n400), .CLK(clk), .Q(\mem<233> ) );
  DFFPOSX1 \mem_reg<234>  ( .D(n399), .CLK(clk), .Q(\mem<234> ) );
  DFFPOSX1 \mem_reg<235>  ( .D(n398), .CLK(clk), .Q(\mem<235> ) );
  DFFPOSX1 \mem_reg<236>  ( .D(n397), .CLK(clk), .Q(\mem<236> ) );
  DFFPOSX1 \mem_reg<237>  ( .D(n396), .CLK(clk), .Q(\mem<237> ) );
  DFFPOSX1 \mem_reg<238>  ( .D(n395), .CLK(clk), .Q(\mem<238> ) );
  DFFPOSX1 \mem_reg<239>  ( .D(n394), .CLK(clk), .Q(\mem<239> ) );
  DFFPOSX1 \mem_reg<240>  ( .D(n393), .CLK(clk), .Q(\mem<240> ) );
  DFFPOSX1 \mem_reg<241>  ( .D(n392), .CLK(clk), .Q(\mem<241> ) );
  DFFPOSX1 \mem_reg<242>  ( .D(n391), .CLK(clk), .Q(\mem<242> ) );
  DFFPOSX1 \mem_reg<243>  ( .D(n390), .CLK(clk), .Q(\mem<243> ) );
  DFFPOSX1 \mem_reg<244>  ( .D(n389), .CLK(clk), .Q(\mem<244> ) );
  DFFPOSX1 \mem_reg<245>  ( .D(n388), .CLK(clk), .Q(\mem<245> ) );
  DFFPOSX1 \mem_reg<246>  ( .D(n387), .CLK(clk), .Q(\mem<246> ) );
  DFFPOSX1 \mem_reg<247>  ( .D(n386), .CLK(clk), .Q(\mem<247> ) );
  DFFPOSX1 \mem_reg<248>  ( .D(n385), .CLK(clk), .Q(\mem<248> ) );
  DFFPOSX1 \mem_reg<249>  ( .D(n384), .CLK(clk), .Q(\mem<249> ) );
  DFFPOSX1 \mem_reg<250>  ( .D(n383), .CLK(clk), .Q(\mem<250> ) );
  DFFPOSX1 \mem_reg<251>  ( .D(n382), .CLK(clk), .Q(\mem<251> ) );
  DFFPOSX1 \mem_reg<252>  ( .D(n381), .CLK(clk), .Q(\mem<252> ) );
  DFFPOSX1 \mem_reg<253>  ( .D(n380), .CLK(clk), .Q(\mem<253> ) );
  DFFPOSX1 \mem_reg<254>  ( .D(n379), .CLK(clk), .Q(\mem<254> ) );
  DFFPOSX1 \mem_reg<255>  ( .D(n378), .CLK(clk), .Q(\mem<255> ) );
  AND2X2 U6 ( .A(N21), .B(n905), .Y(n355) );
  AND2X2 U7 ( .A(N21), .B(n995), .Y(n364) );
  AND2X2 U8 ( .A(n993), .B(n915), .Y(n356) );
  AND2X2 U9 ( .A(n993), .B(n992), .Y(n358) );
  OAI21X1 U49 ( .A(n81), .B(n988), .C(n42), .Y(n378) );
  OAI21X1 U50 ( .A(n32), .B(n986), .C(\mem<255> ), .Y(n42) );
  OAI21X1 U51 ( .A(n989), .B(n78), .C(n46), .Y(n379) );
  OAI21X1 U52 ( .A(n987), .B(n30), .C(\mem<254> ), .Y(n46) );
  OAI21X1 U53 ( .A(n989), .B(n938), .C(n49), .Y(n380) );
  OAI21X1 U54 ( .A(n987), .B(n28), .C(\mem<253> ), .Y(n49) );
  OAI21X1 U55 ( .A(n989), .B(n937), .C(n52), .Y(n381) );
  OAI21X1 U56 ( .A(n987), .B(n26), .C(\mem<252> ), .Y(n52) );
  OAI21X1 U57 ( .A(n989), .B(n75), .C(n55), .Y(n382) );
  OAI21X1 U58 ( .A(n987), .B(n24), .C(\mem<251> ), .Y(n55) );
  OAI21X1 U59 ( .A(n989), .B(n72), .C(n58), .Y(n383) );
  OAI21X1 U60 ( .A(n987), .B(n22), .C(\mem<250> ), .Y(n58) );
  OAI21X1 U61 ( .A(n989), .B(n69), .C(n61), .Y(n384) );
  OAI21X1 U62 ( .A(n987), .B(n20), .C(\mem<249> ), .Y(n61) );
  OAI21X1 U63 ( .A(n989), .B(n66), .C(n64), .Y(n385) );
  OAI21X1 U64 ( .A(n987), .B(n18), .C(\mem<248> ), .Y(n64) );
  OAI21X1 U65 ( .A(n989), .B(n936), .C(n67), .Y(n386) );
  OAI21X1 U66 ( .A(n987), .B(n16), .C(\mem<247> ), .Y(n67) );
  OAI21X1 U67 ( .A(n988), .B(n935), .C(n70), .Y(n387) );
  OAI21X1 U68 ( .A(n986), .B(n14), .C(\mem<246> ), .Y(n70) );
  OAI21X1 U69 ( .A(n988), .B(n934), .C(n73), .Y(n388) );
  OAI21X1 U70 ( .A(n986), .B(n12), .C(\mem<245> ), .Y(n73) );
  OAI21X1 U71 ( .A(n988), .B(n933), .C(n76), .Y(n389) );
  OAI21X1 U72 ( .A(n986), .B(n10), .C(\mem<244> ), .Y(n76) );
  OAI21X1 U73 ( .A(n988), .B(n932), .C(n79), .Y(n390) );
  OAI21X1 U74 ( .A(n986), .B(n8), .C(\mem<243> ), .Y(n79) );
  OAI21X1 U75 ( .A(n988), .B(n931), .C(n82), .Y(n391) );
  OAI21X1 U76 ( .A(n986), .B(n6), .C(\mem<242> ), .Y(n82) );
  OAI21X1 U77 ( .A(n988), .B(n930), .C(n85), .Y(n392) );
  OAI21X1 U78 ( .A(n986), .B(n4), .C(\mem<241> ), .Y(n85) );
  OAI21X1 U79 ( .A(n988), .B(n924), .C(n88), .Y(n393) );
  OAI21X1 U80 ( .A(n986), .B(n2), .C(\mem<240> ), .Y(n88) );
  OAI21X1 U83 ( .A(n81), .B(n985), .C(n94), .Y(n394) );
  OAI21X1 U84 ( .A(n32), .B(n983), .C(\mem<239> ), .Y(n94) );
  OAI21X1 U85 ( .A(n78), .B(n985), .C(n96), .Y(n395) );
  OAI21X1 U86 ( .A(n30), .B(n983), .C(\mem<238> ), .Y(n96) );
  OAI21X1 U87 ( .A(n938), .B(n985), .C(n97), .Y(n396) );
  OAI21X1 U88 ( .A(n28), .B(n983), .C(\mem<237> ), .Y(n97) );
  OAI21X1 U89 ( .A(n937), .B(n985), .C(n98), .Y(n397) );
  OAI21X1 U90 ( .A(n26), .B(n983), .C(\mem<236> ), .Y(n98) );
  OAI21X1 U91 ( .A(n75), .B(n985), .C(n99), .Y(n398) );
  OAI21X1 U92 ( .A(n24), .B(n983), .C(\mem<235> ), .Y(n99) );
  OAI21X1 U93 ( .A(n72), .B(n985), .C(n100), .Y(n399) );
  OAI21X1 U94 ( .A(n22), .B(n983), .C(\mem<234> ), .Y(n100) );
  OAI21X1 U95 ( .A(n69), .B(n985), .C(n101), .Y(n400) );
  OAI21X1 U96 ( .A(n20), .B(n983), .C(\mem<233> ), .Y(n101) );
  OAI21X1 U97 ( .A(n66), .B(n985), .C(n102), .Y(n401) );
  OAI21X1 U98 ( .A(n18), .B(n983), .C(\mem<232> ), .Y(n102) );
  OAI21X1 U99 ( .A(n936), .B(n984), .C(n103), .Y(n402) );
  OAI21X1 U100 ( .A(n16), .B(n982), .C(\mem<231> ), .Y(n103) );
  OAI21X1 U101 ( .A(n935), .B(n984), .C(n104), .Y(n403) );
  OAI21X1 U102 ( .A(n14), .B(n982), .C(\mem<230> ), .Y(n104) );
  OAI21X1 U103 ( .A(n934), .B(n984), .C(n105), .Y(n404) );
  OAI21X1 U104 ( .A(n12), .B(n982), .C(\mem<229> ), .Y(n105) );
  OAI21X1 U105 ( .A(n933), .B(n984), .C(n106), .Y(n405) );
  OAI21X1 U106 ( .A(n10), .B(n982), .C(\mem<228> ), .Y(n106) );
  OAI21X1 U107 ( .A(n932), .B(n984), .C(n107), .Y(n406) );
  OAI21X1 U108 ( .A(n8), .B(n982), .C(\mem<227> ), .Y(n107) );
  OAI21X1 U109 ( .A(n931), .B(n984), .C(n108), .Y(n407) );
  OAI21X1 U110 ( .A(n6), .B(n982), .C(\mem<226> ), .Y(n108) );
  OAI21X1 U111 ( .A(n930), .B(n984), .C(n109), .Y(n408) );
  OAI21X1 U112 ( .A(n4), .B(n982), .C(\mem<225> ), .Y(n109) );
  OAI21X1 U113 ( .A(n924), .B(n984), .C(n110), .Y(n409) );
  OAI21X1 U114 ( .A(n2), .B(n982), .C(\mem<224> ), .Y(n110) );
  OAI21X1 U117 ( .A(n81), .B(n981), .C(n113), .Y(n410) );
  OAI21X1 U118 ( .A(n32), .B(n979), .C(\mem<223> ), .Y(n113) );
  OAI21X1 U119 ( .A(n78), .B(n981), .C(n115), .Y(n411) );
  OAI21X1 U120 ( .A(n30), .B(n979), .C(\mem<222> ), .Y(n115) );
  OAI21X1 U121 ( .A(n938), .B(n981), .C(n116), .Y(n412) );
  OAI21X1 U122 ( .A(n28), .B(n979), .C(\mem<221> ), .Y(n116) );
  OAI21X1 U123 ( .A(n937), .B(n981), .C(n117), .Y(n413) );
  OAI21X1 U124 ( .A(n26), .B(n979), .C(\mem<220> ), .Y(n117) );
  OAI21X1 U125 ( .A(n75), .B(n981), .C(n118), .Y(n414) );
  OAI21X1 U126 ( .A(n24), .B(n979), .C(\mem<219> ), .Y(n118) );
  OAI21X1 U127 ( .A(n72), .B(n981), .C(n119), .Y(n415) );
  OAI21X1 U128 ( .A(n22), .B(n979), .C(\mem<218> ), .Y(n119) );
  OAI21X1 U129 ( .A(n69), .B(n981), .C(n120), .Y(n416) );
  OAI21X1 U130 ( .A(n20), .B(n979), .C(\mem<217> ), .Y(n120) );
  OAI21X1 U131 ( .A(n66), .B(n981), .C(n121), .Y(n417) );
  OAI21X1 U132 ( .A(n18), .B(n979), .C(\mem<216> ), .Y(n121) );
  OAI21X1 U133 ( .A(n936), .B(n980), .C(n122), .Y(n418) );
  OAI21X1 U134 ( .A(n16), .B(n979), .C(\mem<215> ), .Y(n122) );
  OAI21X1 U135 ( .A(n935), .B(n980), .C(n123), .Y(n419) );
  OAI21X1 U136 ( .A(n14), .B(n979), .C(\mem<214> ), .Y(n123) );
  OAI21X1 U137 ( .A(n934), .B(n980), .C(n124), .Y(n420) );
  OAI21X1 U138 ( .A(n12), .B(n979), .C(\mem<213> ), .Y(n124) );
  OAI21X1 U139 ( .A(n933), .B(n980), .C(n125), .Y(n421) );
  OAI21X1 U140 ( .A(n10), .B(n979), .C(\mem<212> ), .Y(n125) );
  OAI21X1 U141 ( .A(n932), .B(n980), .C(n126), .Y(n422) );
  OAI21X1 U142 ( .A(n8), .B(n979), .C(\mem<211> ), .Y(n126) );
  OAI21X1 U143 ( .A(n931), .B(n980), .C(n127), .Y(n423) );
  OAI21X1 U144 ( .A(n6), .B(n979), .C(\mem<210> ), .Y(n127) );
  OAI21X1 U145 ( .A(n930), .B(n980), .C(n128), .Y(n424) );
  OAI21X1 U146 ( .A(n4), .B(n979), .C(\mem<209> ), .Y(n128) );
  OAI21X1 U147 ( .A(n924), .B(n980), .C(n129), .Y(n425) );
  OAI21X1 U148 ( .A(n2), .B(n979), .C(\mem<208> ), .Y(n129) );
  OAI21X1 U151 ( .A(n81), .B(n978), .C(n132), .Y(n426) );
  OAI21X1 U152 ( .A(n32), .B(n976), .C(\mem<207> ), .Y(n132) );
  OAI21X1 U153 ( .A(n78), .B(n978), .C(n134), .Y(n427) );
  OAI21X1 U154 ( .A(n30), .B(n976), .C(\mem<206> ), .Y(n134) );
  OAI21X1 U155 ( .A(n938), .B(n978), .C(n135), .Y(n428) );
  OAI21X1 U156 ( .A(n28), .B(n976), .C(\mem<205> ), .Y(n135) );
  OAI21X1 U157 ( .A(n937), .B(n978), .C(n136), .Y(n429) );
  OAI21X1 U158 ( .A(n26), .B(n976), .C(\mem<204> ), .Y(n136) );
  OAI21X1 U159 ( .A(n75), .B(n978), .C(n137), .Y(n430) );
  OAI21X1 U160 ( .A(n24), .B(n976), .C(\mem<203> ), .Y(n137) );
  OAI21X1 U161 ( .A(n72), .B(n978), .C(n138), .Y(n431) );
  OAI21X1 U162 ( .A(n22), .B(n976), .C(\mem<202> ), .Y(n138) );
  OAI21X1 U163 ( .A(n69), .B(n978), .C(n139), .Y(n432) );
  OAI21X1 U164 ( .A(n20), .B(n976), .C(\mem<201> ), .Y(n139) );
  OAI21X1 U165 ( .A(n66), .B(n978), .C(n140), .Y(n433) );
  OAI21X1 U166 ( .A(n18), .B(n976), .C(\mem<200> ), .Y(n140) );
  OAI21X1 U167 ( .A(n936), .B(n977), .C(n141), .Y(n434) );
  OAI21X1 U168 ( .A(n16), .B(n976), .C(\mem<199> ), .Y(n141) );
  OAI21X1 U169 ( .A(n935), .B(n977), .C(n142), .Y(n435) );
  OAI21X1 U170 ( .A(n14), .B(n976), .C(\mem<198> ), .Y(n142) );
  OAI21X1 U171 ( .A(n934), .B(n977), .C(n143), .Y(n436) );
  OAI21X1 U172 ( .A(n12), .B(n976), .C(\mem<197> ), .Y(n143) );
  OAI21X1 U173 ( .A(n933), .B(n977), .C(n144), .Y(n437) );
  OAI21X1 U174 ( .A(n10), .B(n976), .C(\mem<196> ), .Y(n144) );
  OAI21X1 U175 ( .A(n932), .B(n977), .C(n145), .Y(n438) );
  OAI21X1 U176 ( .A(n8), .B(n976), .C(\mem<195> ), .Y(n145) );
  OAI21X1 U177 ( .A(n931), .B(n977), .C(n146), .Y(n439) );
  OAI21X1 U178 ( .A(n6), .B(n976), .C(\mem<194> ), .Y(n146) );
  OAI21X1 U179 ( .A(n930), .B(n977), .C(n147), .Y(n440) );
  OAI21X1 U180 ( .A(n4), .B(n976), .C(\mem<193> ), .Y(n147) );
  OAI21X1 U181 ( .A(n924), .B(n977), .C(n148), .Y(n441) );
  OAI21X1 U182 ( .A(n2), .B(n976), .C(\mem<192> ), .Y(n148) );
  OAI21X1 U185 ( .A(n81), .B(n975), .C(n151), .Y(n442) );
  OAI21X1 U186 ( .A(n32), .B(n973), .C(\mem<191> ), .Y(n151) );
  OAI21X1 U187 ( .A(n78), .B(n975), .C(n153), .Y(n443) );
  OAI21X1 U188 ( .A(n30), .B(n973), .C(\mem<190> ), .Y(n153) );
  OAI21X1 U189 ( .A(n938), .B(n975), .C(n154), .Y(n444) );
  OAI21X1 U190 ( .A(n28), .B(n973), .C(\mem<189> ), .Y(n154) );
  OAI21X1 U191 ( .A(n937), .B(n975), .C(n155), .Y(n445) );
  OAI21X1 U192 ( .A(n26), .B(n973), .C(\mem<188> ), .Y(n155) );
  OAI21X1 U193 ( .A(n75), .B(n975), .C(n156), .Y(n446) );
  OAI21X1 U194 ( .A(n24), .B(n973), .C(\mem<187> ), .Y(n156) );
  OAI21X1 U195 ( .A(n72), .B(n975), .C(n157), .Y(n447) );
  OAI21X1 U196 ( .A(n22), .B(n973), .C(\mem<186> ), .Y(n157) );
  OAI21X1 U197 ( .A(n69), .B(n975), .C(n158), .Y(n448) );
  OAI21X1 U198 ( .A(n20), .B(n973), .C(\mem<185> ), .Y(n158) );
  OAI21X1 U199 ( .A(n66), .B(n975), .C(n159), .Y(n449) );
  OAI21X1 U200 ( .A(n18), .B(n973), .C(\mem<184> ), .Y(n159) );
  OAI21X1 U201 ( .A(n936), .B(n974), .C(n160), .Y(n450) );
  OAI21X1 U202 ( .A(n16), .B(n972), .C(\mem<183> ), .Y(n160) );
  OAI21X1 U203 ( .A(n935), .B(n974), .C(n161), .Y(n451) );
  OAI21X1 U204 ( .A(n14), .B(n972), .C(\mem<182> ), .Y(n161) );
  OAI21X1 U205 ( .A(n934), .B(n974), .C(n162), .Y(n452) );
  OAI21X1 U206 ( .A(n12), .B(n972), .C(\mem<181> ), .Y(n162) );
  OAI21X1 U207 ( .A(n933), .B(n974), .C(n163), .Y(n453) );
  OAI21X1 U208 ( .A(n10), .B(n972), .C(\mem<180> ), .Y(n163) );
  OAI21X1 U209 ( .A(n932), .B(n974), .C(n164), .Y(n454) );
  OAI21X1 U210 ( .A(n8), .B(n972), .C(\mem<179> ), .Y(n164) );
  OAI21X1 U211 ( .A(n931), .B(n974), .C(n165), .Y(n455) );
  OAI21X1 U212 ( .A(n6), .B(n972), .C(\mem<178> ), .Y(n165) );
  OAI21X1 U213 ( .A(n930), .B(n974), .C(n166), .Y(n456) );
  OAI21X1 U214 ( .A(n4), .B(n972), .C(\mem<177> ), .Y(n166) );
  OAI21X1 U215 ( .A(n924), .B(n974), .C(n167), .Y(n457) );
  OAI21X1 U216 ( .A(n2), .B(n972), .C(\mem<176> ), .Y(n167) );
  OAI21X1 U219 ( .A(n81), .B(n971), .C(n170), .Y(n458) );
  OAI21X1 U220 ( .A(n32), .B(n969), .C(\mem<175> ), .Y(n170) );
  OAI21X1 U221 ( .A(n78), .B(n971), .C(n172), .Y(n459) );
  OAI21X1 U222 ( .A(n30), .B(n969), .C(\mem<174> ), .Y(n172) );
  OAI21X1 U223 ( .A(n938), .B(n971), .C(n173), .Y(n460) );
  OAI21X1 U224 ( .A(n28), .B(n969), .C(\mem<173> ), .Y(n173) );
  OAI21X1 U225 ( .A(n937), .B(n971), .C(n174), .Y(n461) );
  OAI21X1 U226 ( .A(n26), .B(n969), .C(\mem<172> ), .Y(n174) );
  OAI21X1 U227 ( .A(n75), .B(n971), .C(n175), .Y(n462) );
  OAI21X1 U228 ( .A(n24), .B(n969), .C(\mem<171> ), .Y(n175) );
  OAI21X1 U229 ( .A(n72), .B(n971), .C(n176), .Y(n463) );
  OAI21X1 U230 ( .A(n22), .B(n969), .C(\mem<170> ), .Y(n176) );
  OAI21X1 U231 ( .A(n69), .B(n971), .C(n177), .Y(n464) );
  OAI21X1 U232 ( .A(n20), .B(n969), .C(\mem<169> ), .Y(n177) );
  OAI21X1 U233 ( .A(n66), .B(n971), .C(n178), .Y(n465) );
  OAI21X1 U234 ( .A(n18), .B(n969), .C(\mem<168> ), .Y(n178) );
  OAI21X1 U235 ( .A(n936), .B(n970), .C(n179), .Y(n466) );
  OAI21X1 U236 ( .A(n16), .B(n968), .C(\mem<167> ), .Y(n179) );
  OAI21X1 U237 ( .A(n935), .B(n970), .C(n180), .Y(n467) );
  OAI21X1 U238 ( .A(n14), .B(n968), .C(\mem<166> ), .Y(n180) );
  OAI21X1 U239 ( .A(n934), .B(n970), .C(n181), .Y(n468) );
  OAI21X1 U240 ( .A(n12), .B(n968), .C(\mem<165> ), .Y(n181) );
  OAI21X1 U241 ( .A(n933), .B(n970), .C(n182), .Y(n469) );
  OAI21X1 U242 ( .A(n10), .B(n968), .C(\mem<164> ), .Y(n182) );
  OAI21X1 U243 ( .A(n932), .B(n970), .C(n183), .Y(n470) );
  OAI21X1 U244 ( .A(n8), .B(n968), .C(\mem<163> ), .Y(n183) );
  OAI21X1 U245 ( .A(n931), .B(n970), .C(n184), .Y(n471) );
  OAI21X1 U246 ( .A(n6), .B(n968), .C(\mem<162> ), .Y(n184) );
  OAI21X1 U247 ( .A(n930), .B(n970), .C(n185), .Y(n472) );
  OAI21X1 U248 ( .A(n4), .B(n968), .C(\mem<161> ), .Y(n185) );
  OAI21X1 U249 ( .A(n924), .B(n970), .C(n186), .Y(n473) );
  OAI21X1 U250 ( .A(n2), .B(n968), .C(\mem<160> ), .Y(n186) );
  OAI21X1 U253 ( .A(n81), .B(n967), .C(n188), .Y(n474) );
  OAI21X1 U254 ( .A(n32), .B(n965), .C(\mem<159> ), .Y(n188) );
  OAI21X1 U255 ( .A(n78), .B(n967), .C(n190), .Y(n475) );
  OAI21X1 U256 ( .A(n30), .B(n965), .C(\mem<158> ), .Y(n190) );
  OAI21X1 U257 ( .A(n938), .B(n967), .C(n191), .Y(n476) );
  OAI21X1 U258 ( .A(n28), .B(n965), .C(\mem<157> ), .Y(n191) );
  OAI21X1 U259 ( .A(n937), .B(n967), .C(n192), .Y(n477) );
  OAI21X1 U260 ( .A(n26), .B(n965), .C(\mem<156> ), .Y(n192) );
  OAI21X1 U261 ( .A(n75), .B(n967), .C(n193), .Y(n478) );
  OAI21X1 U262 ( .A(n24), .B(n965), .C(\mem<155> ), .Y(n193) );
  OAI21X1 U263 ( .A(n72), .B(n967), .C(n194), .Y(n479) );
  OAI21X1 U264 ( .A(n22), .B(n965), .C(\mem<154> ), .Y(n194) );
  OAI21X1 U265 ( .A(n69), .B(n967), .C(n195), .Y(n480) );
  OAI21X1 U266 ( .A(n20), .B(n965), .C(\mem<153> ), .Y(n195) );
  OAI21X1 U267 ( .A(n66), .B(n967), .C(n196), .Y(n481) );
  OAI21X1 U268 ( .A(n18), .B(n965), .C(\mem<152> ), .Y(n196) );
  OAI21X1 U269 ( .A(n936), .B(n966), .C(n197), .Y(n482) );
  OAI21X1 U270 ( .A(n16), .B(n964), .C(\mem<151> ), .Y(n197) );
  OAI21X1 U271 ( .A(n935), .B(n966), .C(n198), .Y(n483) );
  OAI21X1 U272 ( .A(n14), .B(n964), .C(\mem<150> ), .Y(n198) );
  OAI21X1 U273 ( .A(n934), .B(n966), .C(n199), .Y(n484) );
  OAI21X1 U274 ( .A(n12), .B(n964), .C(\mem<149> ), .Y(n199) );
  OAI21X1 U275 ( .A(n933), .B(n966), .C(n200), .Y(n485) );
  OAI21X1 U276 ( .A(n10), .B(n964), .C(\mem<148> ), .Y(n200) );
  OAI21X1 U277 ( .A(n932), .B(n966), .C(n201), .Y(n486) );
  OAI21X1 U278 ( .A(n8), .B(n964), .C(\mem<147> ), .Y(n201) );
  OAI21X1 U279 ( .A(n931), .B(n966), .C(n202), .Y(n487) );
  OAI21X1 U280 ( .A(n6), .B(n964), .C(\mem<146> ), .Y(n202) );
  OAI21X1 U281 ( .A(n930), .B(n966), .C(n203), .Y(n488) );
  OAI21X1 U282 ( .A(n4), .B(n964), .C(\mem<145> ), .Y(n203) );
  OAI21X1 U283 ( .A(n924), .B(n966), .C(n204), .Y(n489) );
  OAI21X1 U284 ( .A(n2), .B(n964), .C(\mem<144> ), .Y(n204) );
  OAI21X1 U287 ( .A(n81), .B(n963), .C(n206), .Y(n490) );
  OAI21X1 U288 ( .A(n32), .B(n961), .C(\mem<143> ), .Y(n206) );
  OAI21X1 U289 ( .A(n78), .B(n963), .C(n208), .Y(n491) );
  OAI21X1 U290 ( .A(n30), .B(n961), .C(\mem<142> ), .Y(n208) );
  OAI21X1 U291 ( .A(n938), .B(n963), .C(n209), .Y(n492) );
  OAI21X1 U292 ( .A(n28), .B(n961), .C(\mem<141> ), .Y(n209) );
  OAI21X1 U293 ( .A(n937), .B(n963), .C(n210), .Y(n493) );
  OAI21X1 U294 ( .A(n26), .B(n961), .C(\mem<140> ), .Y(n210) );
  OAI21X1 U295 ( .A(n75), .B(n963), .C(n211), .Y(n494) );
  OAI21X1 U296 ( .A(n24), .B(n961), .C(\mem<139> ), .Y(n211) );
  OAI21X1 U297 ( .A(n72), .B(n963), .C(n212), .Y(n495) );
  OAI21X1 U298 ( .A(n22), .B(n961), .C(\mem<138> ), .Y(n212) );
  OAI21X1 U299 ( .A(n69), .B(n963), .C(n213), .Y(n496) );
  OAI21X1 U300 ( .A(n20), .B(n961), .C(\mem<137> ), .Y(n213) );
  OAI21X1 U301 ( .A(n66), .B(n963), .C(n214), .Y(n497) );
  OAI21X1 U302 ( .A(n18), .B(n961), .C(\mem<136> ), .Y(n214) );
  OAI21X1 U303 ( .A(n936), .B(n962), .C(n215), .Y(n498) );
  OAI21X1 U304 ( .A(n16), .B(n960), .C(\mem<135> ), .Y(n215) );
  OAI21X1 U305 ( .A(n935), .B(n962), .C(n216), .Y(n499) );
  OAI21X1 U306 ( .A(n14), .B(n960), .C(\mem<134> ), .Y(n216) );
  OAI21X1 U307 ( .A(n934), .B(n962), .C(n217), .Y(n500) );
  OAI21X1 U308 ( .A(n12), .B(n960), .C(\mem<133> ), .Y(n217) );
  OAI21X1 U309 ( .A(n933), .B(n962), .C(n218), .Y(n501) );
  OAI21X1 U310 ( .A(n10), .B(n960), .C(\mem<132> ), .Y(n218) );
  OAI21X1 U311 ( .A(n932), .B(n962), .C(n219), .Y(n502) );
  OAI21X1 U312 ( .A(n8), .B(n960), .C(\mem<131> ), .Y(n219) );
  OAI21X1 U313 ( .A(n931), .B(n962), .C(n220), .Y(n503) );
  OAI21X1 U314 ( .A(n6), .B(n960), .C(\mem<130> ), .Y(n220) );
  OAI21X1 U315 ( .A(n930), .B(n962), .C(n221), .Y(n504) );
  OAI21X1 U316 ( .A(n4), .B(n960), .C(\mem<129> ), .Y(n221) );
  OAI21X1 U317 ( .A(n924), .B(n962), .C(n222), .Y(n505) );
  OAI21X1 U318 ( .A(n2), .B(n960), .C(\mem<128> ), .Y(n222) );
  OAI21X1 U321 ( .A(n81), .B(n959), .C(n224), .Y(n506) );
  OAI21X1 U322 ( .A(n32), .B(n957), .C(\mem<127> ), .Y(n224) );
  OAI21X1 U323 ( .A(n78), .B(n959), .C(n226), .Y(n507) );
  OAI21X1 U324 ( .A(n30), .B(n957), .C(\mem<126> ), .Y(n226) );
  OAI21X1 U325 ( .A(n938), .B(n959), .C(n227), .Y(n508) );
  OAI21X1 U326 ( .A(n28), .B(n957), .C(\mem<125> ), .Y(n227) );
  OAI21X1 U327 ( .A(n937), .B(n959), .C(n228), .Y(n509) );
  OAI21X1 U328 ( .A(n26), .B(n957), .C(\mem<124> ), .Y(n228) );
  OAI21X1 U329 ( .A(n75), .B(n959), .C(n229), .Y(n510) );
  OAI21X1 U330 ( .A(n24), .B(n957), .C(\mem<123> ), .Y(n229) );
  OAI21X1 U331 ( .A(n72), .B(n959), .C(n230), .Y(n511) );
  OAI21X1 U332 ( .A(n22), .B(n957), .C(\mem<122> ), .Y(n230) );
  OAI21X1 U333 ( .A(n69), .B(n959), .C(n231), .Y(n512) );
  OAI21X1 U334 ( .A(n20), .B(n957), .C(\mem<121> ), .Y(n231) );
  OAI21X1 U335 ( .A(n66), .B(n959), .C(n232), .Y(n513) );
  OAI21X1 U336 ( .A(n18), .B(n957), .C(\mem<120> ), .Y(n232) );
  OAI21X1 U337 ( .A(n936), .B(n958), .C(n233), .Y(n514) );
  OAI21X1 U338 ( .A(n16), .B(n957), .C(\mem<119> ), .Y(n233) );
  OAI21X1 U339 ( .A(n935), .B(n958), .C(n234), .Y(n515) );
  OAI21X1 U340 ( .A(n14), .B(n957), .C(\mem<118> ), .Y(n234) );
  OAI21X1 U341 ( .A(n934), .B(n958), .C(n235), .Y(n516) );
  OAI21X1 U342 ( .A(n12), .B(n957), .C(\mem<117> ), .Y(n235) );
  OAI21X1 U343 ( .A(n933), .B(n958), .C(n236), .Y(n517) );
  OAI21X1 U344 ( .A(n10), .B(n957), .C(\mem<116> ), .Y(n236) );
  OAI21X1 U345 ( .A(n932), .B(n958), .C(n237), .Y(n518) );
  OAI21X1 U346 ( .A(n8), .B(n957), .C(\mem<115> ), .Y(n237) );
  OAI21X1 U347 ( .A(n931), .B(n958), .C(n238), .Y(n519) );
  OAI21X1 U348 ( .A(n6), .B(n957), .C(\mem<114> ), .Y(n238) );
  OAI21X1 U349 ( .A(n930), .B(n958), .C(n239), .Y(n520) );
  OAI21X1 U350 ( .A(n4), .B(n957), .C(\mem<113> ), .Y(n239) );
  OAI21X1 U351 ( .A(n924), .B(n958), .C(n240), .Y(n521) );
  OAI21X1 U352 ( .A(n2), .B(n957), .C(\mem<112> ), .Y(n240) );
  OAI21X1 U355 ( .A(n81), .B(n956), .C(n243), .Y(n522) );
  OAI21X1 U356 ( .A(n32), .B(n954), .C(\mem<111> ), .Y(n243) );
  OAI21X1 U357 ( .A(n78), .B(n956), .C(n245), .Y(n523) );
  OAI21X1 U358 ( .A(n30), .B(n954), .C(\mem<110> ), .Y(n245) );
  OAI21X1 U359 ( .A(n938), .B(n956), .C(n246), .Y(n524) );
  OAI21X1 U360 ( .A(n28), .B(n954), .C(\mem<109> ), .Y(n246) );
  OAI21X1 U361 ( .A(n937), .B(n956), .C(n247), .Y(n525) );
  OAI21X1 U362 ( .A(n26), .B(n954), .C(\mem<108> ), .Y(n247) );
  OAI21X1 U363 ( .A(n75), .B(n956), .C(n248), .Y(n526) );
  OAI21X1 U364 ( .A(n24), .B(n954), .C(\mem<107> ), .Y(n248) );
  OAI21X1 U365 ( .A(n72), .B(n956), .C(n249), .Y(n527) );
  OAI21X1 U366 ( .A(n22), .B(n954), .C(\mem<106> ), .Y(n249) );
  OAI21X1 U367 ( .A(n69), .B(n956), .C(n250), .Y(n528) );
  OAI21X1 U368 ( .A(n20), .B(n954), .C(\mem<105> ), .Y(n250) );
  OAI21X1 U369 ( .A(n66), .B(n956), .C(n251), .Y(n529) );
  OAI21X1 U370 ( .A(n18), .B(n954), .C(\mem<104> ), .Y(n251) );
  OAI21X1 U371 ( .A(n936), .B(n955), .C(n252), .Y(n530) );
  OAI21X1 U372 ( .A(n16), .B(n954), .C(\mem<103> ), .Y(n252) );
  OAI21X1 U373 ( .A(n935), .B(n955), .C(n253), .Y(n531) );
  OAI21X1 U374 ( .A(n14), .B(n954), .C(\mem<102> ), .Y(n253) );
  OAI21X1 U375 ( .A(n934), .B(n955), .C(n254), .Y(n532) );
  OAI21X1 U376 ( .A(n12), .B(n954), .C(\mem<101> ), .Y(n254) );
  OAI21X1 U377 ( .A(n933), .B(n955), .C(n255), .Y(n533) );
  OAI21X1 U378 ( .A(n10), .B(n954), .C(\mem<100> ), .Y(n255) );
  OAI21X1 U379 ( .A(n932), .B(n955), .C(n256), .Y(n534) );
  OAI21X1 U380 ( .A(n8), .B(n954), .C(\mem<99> ), .Y(n256) );
  OAI21X1 U381 ( .A(n931), .B(n955), .C(n257), .Y(n535) );
  OAI21X1 U382 ( .A(n6), .B(n954), .C(\mem<98> ), .Y(n257) );
  OAI21X1 U383 ( .A(n930), .B(n955), .C(n258), .Y(n536) );
  OAI21X1 U384 ( .A(n4), .B(n954), .C(\mem<97> ), .Y(n258) );
  OAI21X1 U385 ( .A(n924), .B(n955), .C(n259), .Y(n537) );
  OAI21X1 U386 ( .A(n2), .B(n954), .C(\mem<96> ), .Y(n259) );
  OAI21X1 U389 ( .A(n81), .B(n953), .C(n261), .Y(n538) );
  OAI21X1 U390 ( .A(n32), .B(n951), .C(\mem<95> ), .Y(n261) );
  OAI21X1 U391 ( .A(n78), .B(n953), .C(n263), .Y(n539) );
  OAI21X1 U392 ( .A(n30), .B(n951), .C(\mem<94> ), .Y(n263) );
  OAI21X1 U393 ( .A(n938), .B(n953), .C(n264), .Y(n540) );
  OAI21X1 U394 ( .A(n28), .B(n951), .C(\mem<93> ), .Y(n264) );
  OAI21X1 U395 ( .A(n937), .B(n953), .C(n265), .Y(n541) );
  OAI21X1 U396 ( .A(n26), .B(n951), .C(\mem<92> ), .Y(n265) );
  OAI21X1 U397 ( .A(n75), .B(n953), .C(n266), .Y(n542) );
  OAI21X1 U398 ( .A(n24), .B(n951), .C(\mem<91> ), .Y(n266) );
  OAI21X1 U399 ( .A(n72), .B(n953), .C(n267), .Y(n543) );
  OAI21X1 U400 ( .A(n22), .B(n951), .C(\mem<90> ), .Y(n267) );
  OAI21X1 U401 ( .A(n69), .B(n953), .C(n268), .Y(n544) );
  OAI21X1 U402 ( .A(n20), .B(n951), .C(\mem<89> ), .Y(n268) );
  OAI21X1 U403 ( .A(n66), .B(n953), .C(n269), .Y(n545) );
  OAI21X1 U404 ( .A(n18), .B(n951), .C(\mem<88> ), .Y(n269) );
  OAI21X1 U405 ( .A(n936), .B(n952), .C(n270), .Y(n546) );
  OAI21X1 U406 ( .A(n16), .B(n951), .C(\mem<87> ), .Y(n270) );
  OAI21X1 U407 ( .A(n935), .B(n952), .C(n271), .Y(n547) );
  OAI21X1 U408 ( .A(n14), .B(n951), .C(\mem<86> ), .Y(n271) );
  OAI21X1 U409 ( .A(n934), .B(n952), .C(n272), .Y(n548) );
  OAI21X1 U410 ( .A(n12), .B(n951), .C(\mem<85> ), .Y(n272) );
  OAI21X1 U411 ( .A(n933), .B(n952), .C(n273), .Y(n549) );
  OAI21X1 U412 ( .A(n10), .B(n951), .C(\mem<84> ), .Y(n273) );
  OAI21X1 U413 ( .A(n932), .B(n952), .C(n274), .Y(n550) );
  OAI21X1 U414 ( .A(n8), .B(n951), .C(\mem<83> ), .Y(n274) );
  OAI21X1 U415 ( .A(n931), .B(n952), .C(n275), .Y(n551) );
  OAI21X1 U416 ( .A(n6), .B(n951), .C(\mem<82> ), .Y(n275) );
  OAI21X1 U417 ( .A(n930), .B(n952), .C(n276), .Y(n552) );
  OAI21X1 U418 ( .A(n4), .B(n951), .C(\mem<81> ), .Y(n276) );
  OAI21X1 U419 ( .A(n924), .B(n952), .C(n277), .Y(n553) );
  OAI21X1 U420 ( .A(n2), .B(n951), .C(\mem<80> ), .Y(n277) );
  OAI21X1 U423 ( .A(n81), .B(n950), .C(n279), .Y(n554) );
  OAI21X1 U424 ( .A(n32), .B(n948), .C(\mem<79> ), .Y(n279) );
  OAI21X1 U425 ( .A(n78), .B(n950), .C(n281), .Y(n555) );
  OAI21X1 U426 ( .A(n30), .B(n948), .C(\mem<78> ), .Y(n281) );
  OAI21X1 U427 ( .A(n938), .B(n950), .C(n282), .Y(n556) );
  OAI21X1 U428 ( .A(n28), .B(n948), .C(\mem<77> ), .Y(n282) );
  OAI21X1 U429 ( .A(n937), .B(n950), .C(n283), .Y(n557) );
  OAI21X1 U430 ( .A(n26), .B(n948), .C(\mem<76> ), .Y(n283) );
  OAI21X1 U431 ( .A(n75), .B(n950), .C(n284), .Y(n558) );
  OAI21X1 U432 ( .A(n24), .B(n948), .C(\mem<75> ), .Y(n284) );
  OAI21X1 U433 ( .A(n72), .B(n950), .C(n285), .Y(n559) );
  OAI21X1 U434 ( .A(n22), .B(n948), .C(\mem<74> ), .Y(n285) );
  OAI21X1 U435 ( .A(n69), .B(n950), .C(n286), .Y(n560) );
  OAI21X1 U436 ( .A(n20), .B(n948), .C(\mem<73> ), .Y(n286) );
  OAI21X1 U437 ( .A(n66), .B(n950), .C(n287), .Y(n561) );
  OAI21X1 U438 ( .A(n18), .B(n948), .C(\mem<72> ), .Y(n287) );
  OAI21X1 U439 ( .A(n936), .B(n949), .C(n288), .Y(n562) );
  OAI21X1 U440 ( .A(n16), .B(n948), .C(\mem<71> ), .Y(n288) );
  OAI21X1 U441 ( .A(n935), .B(n949), .C(n289), .Y(n563) );
  OAI21X1 U442 ( .A(n14), .B(n948), .C(\mem<70> ), .Y(n289) );
  OAI21X1 U443 ( .A(n934), .B(n949), .C(n290), .Y(n564) );
  OAI21X1 U444 ( .A(n12), .B(n948), .C(\mem<69> ), .Y(n290) );
  OAI21X1 U445 ( .A(n933), .B(n949), .C(n291), .Y(n565) );
  OAI21X1 U446 ( .A(n10), .B(n948), .C(\mem<68> ), .Y(n291) );
  OAI21X1 U447 ( .A(n932), .B(n949), .C(n292), .Y(n566) );
  OAI21X1 U448 ( .A(n8), .B(n948), .C(\mem<67> ), .Y(n292) );
  OAI21X1 U449 ( .A(n931), .B(n949), .C(n293), .Y(n567) );
  OAI21X1 U450 ( .A(n6), .B(n948), .C(\mem<66> ), .Y(n293) );
  OAI21X1 U451 ( .A(n930), .B(n949), .C(n294), .Y(n568) );
  OAI21X1 U452 ( .A(n4), .B(n948), .C(\mem<65> ), .Y(n294) );
  OAI21X1 U453 ( .A(n924), .B(n949), .C(n295), .Y(n569) );
  OAI21X1 U454 ( .A(n2), .B(n948), .C(\mem<64> ), .Y(n295) );
  OAI21X1 U458 ( .A(n81), .B(n947), .C(n297), .Y(n570) );
  OAI21X1 U459 ( .A(n32), .B(n945), .C(\mem<63> ), .Y(n297) );
  OAI21X1 U460 ( .A(n78), .B(n947), .C(n299), .Y(n571) );
  OAI21X1 U461 ( .A(n30), .B(n945), .C(\mem<62> ), .Y(n299) );
  OAI21X1 U462 ( .A(n938), .B(n947), .C(n300), .Y(n572) );
  OAI21X1 U463 ( .A(n28), .B(n945), .C(\mem<61> ), .Y(n300) );
  OAI21X1 U464 ( .A(n937), .B(n947), .C(n301), .Y(n573) );
  OAI21X1 U465 ( .A(n26), .B(n945), .C(\mem<60> ), .Y(n301) );
  OAI21X1 U466 ( .A(n75), .B(n947), .C(n302), .Y(n574) );
  OAI21X1 U467 ( .A(n24), .B(n945), .C(\mem<59> ), .Y(n302) );
  OAI21X1 U468 ( .A(n72), .B(n947), .C(n303), .Y(n575) );
  OAI21X1 U469 ( .A(n22), .B(n945), .C(\mem<58> ), .Y(n303) );
  OAI21X1 U470 ( .A(n69), .B(n947), .C(n304), .Y(n576) );
  OAI21X1 U471 ( .A(n20), .B(n945), .C(\mem<57> ), .Y(n304) );
  OAI21X1 U472 ( .A(n66), .B(n947), .C(n305), .Y(n577) );
  OAI21X1 U473 ( .A(n18), .B(n945), .C(\mem<56> ), .Y(n305) );
  OAI21X1 U474 ( .A(n936), .B(n946), .C(n306), .Y(n578) );
  OAI21X1 U475 ( .A(n16), .B(n945), .C(\mem<55> ), .Y(n306) );
  OAI21X1 U476 ( .A(n935), .B(n946), .C(n307), .Y(n579) );
  OAI21X1 U477 ( .A(n14), .B(n945), .C(\mem<54> ), .Y(n307) );
  OAI21X1 U478 ( .A(n934), .B(n946), .C(n308), .Y(n580) );
  OAI21X1 U479 ( .A(n12), .B(n945), .C(\mem<53> ), .Y(n308) );
  OAI21X1 U480 ( .A(n933), .B(n946), .C(n309), .Y(n581) );
  OAI21X1 U481 ( .A(n10), .B(n945), .C(\mem<52> ), .Y(n309) );
  OAI21X1 U482 ( .A(n932), .B(n946), .C(n310), .Y(n582) );
  OAI21X1 U483 ( .A(n8), .B(n945), .C(\mem<51> ), .Y(n310) );
  OAI21X1 U484 ( .A(n931), .B(n946), .C(n311), .Y(n583) );
  OAI21X1 U485 ( .A(n6), .B(n945), .C(\mem<50> ), .Y(n311) );
  OAI21X1 U486 ( .A(n930), .B(n946), .C(n312), .Y(n584) );
  OAI21X1 U487 ( .A(n4), .B(n945), .C(\mem<49> ), .Y(n312) );
  OAI21X1 U488 ( .A(n924), .B(n946), .C(n313), .Y(n585) );
  OAI21X1 U489 ( .A(n2), .B(n945), .C(\mem<48> ), .Y(n313) );
  OAI21X1 U492 ( .A(n81), .B(n944), .C(n316), .Y(n586) );
  OAI21X1 U493 ( .A(n32), .B(n942), .C(\mem<47> ), .Y(n316) );
  OAI21X1 U494 ( .A(n78), .B(n944), .C(n318), .Y(n587) );
  OAI21X1 U495 ( .A(n30), .B(n942), .C(\mem<46> ), .Y(n318) );
  OAI21X1 U496 ( .A(n938), .B(n944), .C(n319), .Y(n588) );
  OAI21X1 U497 ( .A(n28), .B(n942), .C(\mem<45> ), .Y(n319) );
  OAI21X1 U498 ( .A(n937), .B(n944), .C(n320), .Y(n589) );
  OAI21X1 U499 ( .A(n26), .B(n942), .C(\mem<44> ), .Y(n320) );
  OAI21X1 U500 ( .A(n75), .B(n944), .C(n321), .Y(n590) );
  OAI21X1 U501 ( .A(n24), .B(n942), .C(\mem<43> ), .Y(n321) );
  OAI21X1 U502 ( .A(n72), .B(n944), .C(n322), .Y(n591) );
  OAI21X1 U503 ( .A(n22), .B(n942), .C(\mem<42> ), .Y(n322) );
  OAI21X1 U504 ( .A(n69), .B(n944), .C(n323), .Y(n592) );
  OAI21X1 U505 ( .A(n20), .B(n942), .C(\mem<41> ), .Y(n323) );
  OAI21X1 U506 ( .A(n66), .B(n944), .C(n324), .Y(n593) );
  OAI21X1 U507 ( .A(n18), .B(n942), .C(\mem<40> ), .Y(n324) );
  OAI21X1 U508 ( .A(n936), .B(n943), .C(n325), .Y(n594) );
  OAI21X1 U509 ( .A(n16), .B(n942), .C(\mem<39> ), .Y(n325) );
  OAI21X1 U510 ( .A(n935), .B(n943), .C(n326), .Y(n595) );
  OAI21X1 U511 ( .A(n14), .B(n942), .C(\mem<38> ), .Y(n326) );
  OAI21X1 U512 ( .A(n934), .B(n943), .C(n327), .Y(n596) );
  OAI21X1 U513 ( .A(n12), .B(n942), .C(\mem<37> ), .Y(n327) );
  OAI21X1 U514 ( .A(n933), .B(n943), .C(n328), .Y(n597) );
  OAI21X1 U515 ( .A(n10), .B(n942), .C(\mem<36> ), .Y(n328) );
  OAI21X1 U516 ( .A(n932), .B(n943), .C(n329), .Y(n598) );
  OAI21X1 U517 ( .A(n8), .B(n942), .C(\mem<35> ), .Y(n329) );
  OAI21X1 U518 ( .A(n931), .B(n943), .C(n330), .Y(n599) );
  OAI21X1 U519 ( .A(n6), .B(n942), .C(\mem<34> ), .Y(n330) );
  OAI21X1 U520 ( .A(n930), .B(n943), .C(n331), .Y(n600) );
  OAI21X1 U521 ( .A(n4), .B(n942), .C(\mem<33> ), .Y(n331) );
  OAI21X1 U522 ( .A(n924), .B(n943), .C(n332), .Y(n601) );
  OAI21X1 U523 ( .A(n2), .B(n942), .C(\mem<32> ), .Y(n332) );
  OAI21X1 U526 ( .A(n81), .B(n941), .C(n334), .Y(n602) );
  OAI21X1 U527 ( .A(n32), .B(n939), .C(\mem<31> ), .Y(n334) );
  OAI21X1 U528 ( .A(n78), .B(n941), .C(n336), .Y(n603) );
  OAI21X1 U529 ( .A(n30), .B(n939), .C(\mem<30> ), .Y(n336) );
  OAI21X1 U530 ( .A(n938), .B(n941), .C(n337), .Y(n604) );
  OAI21X1 U531 ( .A(n28), .B(n939), .C(\mem<29> ), .Y(n337) );
  OAI21X1 U532 ( .A(n937), .B(n941), .C(n338), .Y(n605) );
  OAI21X1 U533 ( .A(n26), .B(n939), .C(\mem<28> ), .Y(n338) );
  OAI21X1 U534 ( .A(n75), .B(n941), .C(n339), .Y(n606) );
  OAI21X1 U535 ( .A(n24), .B(n939), .C(\mem<27> ), .Y(n339) );
  OAI21X1 U536 ( .A(n72), .B(n941), .C(n340), .Y(n607) );
  OAI21X1 U537 ( .A(n22), .B(n939), .C(\mem<26> ), .Y(n340) );
  OAI21X1 U538 ( .A(n69), .B(n941), .C(n341), .Y(n608) );
  OAI21X1 U539 ( .A(n20), .B(n939), .C(\mem<25> ), .Y(n341) );
  OAI21X1 U540 ( .A(n66), .B(n941), .C(n342), .Y(n609) );
  OAI21X1 U541 ( .A(n18), .B(n939), .C(\mem<24> ), .Y(n342) );
  OAI21X1 U542 ( .A(n936), .B(n940), .C(n343), .Y(n610) );
  OAI21X1 U543 ( .A(n16), .B(n939), .C(\mem<23> ), .Y(n343) );
  OAI21X1 U544 ( .A(n935), .B(n940), .C(n344), .Y(n611) );
  OAI21X1 U545 ( .A(n14), .B(n939), .C(\mem<22> ), .Y(n344) );
  OAI21X1 U546 ( .A(n934), .B(n940), .C(n345), .Y(n612) );
  OAI21X1 U547 ( .A(n12), .B(n939), .C(\mem<21> ), .Y(n345) );
  OAI21X1 U548 ( .A(n933), .B(n940), .C(n346), .Y(n613) );
  OAI21X1 U549 ( .A(n10), .B(n939), .C(\mem<20> ), .Y(n346) );
  OAI21X1 U550 ( .A(n932), .B(n940), .C(n347), .Y(n614) );
  OAI21X1 U551 ( .A(n8), .B(n939), .C(\mem<19> ), .Y(n347) );
  OAI21X1 U552 ( .A(n931), .B(n940), .C(n348), .Y(n615) );
  OAI21X1 U553 ( .A(n6), .B(n939), .C(\mem<18> ), .Y(n348) );
  OAI21X1 U554 ( .A(n930), .B(n940), .C(n349), .Y(n616) );
  OAI21X1 U555 ( .A(n4), .B(n939), .C(\mem<17> ), .Y(n349) );
  OAI21X1 U556 ( .A(n924), .B(n940), .C(n350), .Y(n617) );
  OAI21X1 U557 ( .A(n2), .B(n939), .C(\mem<16> ), .Y(n350) );
  OAI21X1 U561 ( .A(n81), .B(n929), .C(n352), .Y(n618) );
  OAI21X1 U562 ( .A(n32), .B(n925), .C(\mem<15> ), .Y(n352) );
  OAI21X1 U565 ( .A(n78), .B(n929), .C(n357), .Y(n619) );
  OAI21X1 U566 ( .A(n30), .B(n925), .C(\mem<14> ), .Y(n357) );
  OAI21X1 U569 ( .A(n938), .B(n929), .C(n359), .Y(n620) );
  OAI21X1 U570 ( .A(n28), .B(n925), .C(\mem<13> ), .Y(n359) );
  OAI21X1 U573 ( .A(n937), .B(n929), .C(n361), .Y(n621) );
  OAI21X1 U574 ( .A(n26), .B(n925), .C(\mem<12> ), .Y(n361) );
  OAI21X1 U577 ( .A(n75), .B(n929), .C(n363), .Y(n622) );
  OAI21X1 U578 ( .A(n24), .B(n925), .C(\mem<11> ), .Y(n363) );
  OAI21X1 U581 ( .A(n72), .B(n929), .C(n365), .Y(n623) );
  OAI21X1 U582 ( .A(n22), .B(n925), .C(\mem<10> ), .Y(n365) );
  OAI21X1 U585 ( .A(n69), .B(n929), .C(n366), .Y(n624) );
  OAI21X1 U586 ( .A(n20), .B(n925), .C(\mem<9> ), .Y(n366) );
  OAI21X1 U589 ( .A(n66), .B(n929), .C(n367), .Y(n625) );
  OAI21X1 U590 ( .A(n18), .B(n925), .C(\mem<8> ), .Y(n367) );
  OAI21X1 U593 ( .A(n936), .B(n928), .C(n368), .Y(n626) );
  OAI21X1 U594 ( .A(n16), .B(n925), .C(\mem<7> ), .Y(n368) );
  OAI21X1 U597 ( .A(n935), .B(n928), .C(n370), .Y(n627) );
  OAI21X1 U598 ( .A(n14), .B(n925), .C(\mem<6> ), .Y(n370) );
  OAI21X1 U601 ( .A(n934), .B(n928), .C(n371), .Y(n628) );
  OAI21X1 U602 ( .A(n12), .B(n925), .C(\mem<5> ), .Y(n371) );
  OAI21X1 U605 ( .A(n933), .B(n928), .C(n372), .Y(n629) );
  OAI21X1 U606 ( .A(n10), .B(n925), .C(\mem<4> ), .Y(n372) );
  OAI21X1 U610 ( .A(n932), .B(n928), .C(n373), .Y(n630) );
  OAI21X1 U611 ( .A(n8), .B(n925), .C(\mem<3> ), .Y(n373) );
  OAI21X1 U614 ( .A(n931), .B(n928), .C(n375), .Y(n631) );
  OAI21X1 U615 ( .A(n6), .B(n925), .C(\mem<2> ), .Y(n375) );
  OAI21X1 U618 ( .A(n930), .B(n928), .C(n376), .Y(n632) );
  OAI21X1 U619 ( .A(n4), .B(n925), .C(\mem<1> ), .Y(n376) );
  OAI21X1 U623 ( .A(n924), .B(n928), .C(n377), .Y(n633) );
  OAI21X1 U624 ( .A(n2), .B(n925), .C(\mem<0> ), .Y(n377) );
  NOR3X1 U634 ( .A(rst), .B(write), .C(n998), .Y(data_out) );
  INVX2 U2 ( .A(n993), .Y(n908) );
  INVX2 U3 ( .A(n995), .Y(n906) );
  INVX1 U4 ( .A(N21), .Y(n902) );
  INVX2 U5 ( .A(n995), .Y(n907) );
  INVX1 U10 ( .A(n902), .Y(n903) );
  INVX1 U11 ( .A(n902), .Y(n904) );
  AND2X1 U12 ( .A(N25), .B(n999), .Y(n168) );
  INVX1 U13 ( .A(N24), .Y(n999) );
  AND2X1 U14 ( .A(data_in), .B(n927), .Y(n90) );
  INVX1 U15 ( .A(n994), .Y(n993) );
  AND2X1 U16 ( .A(N25), .B(N24), .Y(n91) );
  BUFX2 U17 ( .A(n90), .Y(n991) );
  AND2X1 U18 ( .A(N23), .B(N22), .Y(n92) );
  AND2X1 U19 ( .A(N23), .B(n996), .Y(n111) );
  BUFX2 U20 ( .A(n90), .Y(n990) );
  INVX1 U21 ( .A(N28), .Y(n998) );
  BUFX2 U22 ( .A(n60), .Y(n927) );
  BUFX2 U23 ( .A(n60), .Y(n926) );
  BUFX2 U24 ( .A(n362), .Y(n989) );
  BUFX2 U25 ( .A(n354), .Y(n986) );
  BUFX2 U26 ( .A(n362), .Y(n988) );
  BUFX2 U27 ( .A(n351), .Y(n985) );
  BUFX2 U28 ( .A(n317), .Y(n982) );
  BUFX2 U29 ( .A(n351), .Y(n984) );
  BUFX2 U30 ( .A(n315), .Y(n981) );
  BUFX2 U31 ( .A(n315), .Y(n980) );
  BUFX2 U32 ( .A(n298), .Y(n978) );
  BUFX2 U33 ( .A(n298), .Y(n977) );
  BUFX2 U34 ( .A(n280), .Y(n975) );
  BUFX2 U35 ( .A(n262), .Y(n972) );
  BUFX2 U36 ( .A(n280), .Y(n974) );
  BUFX2 U37 ( .A(n244), .Y(n971) );
  BUFX2 U38 ( .A(n241), .Y(n968) );
  BUFX2 U39 ( .A(n244), .Y(n970) );
  BUFX2 U40 ( .A(n223), .Y(n967) );
  BUFX2 U41 ( .A(n205), .Y(n964) );
  BUFX2 U42 ( .A(n223), .Y(n966) );
  BUFX2 U43 ( .A(n187), .Y(n963) );
  BUFX2 U44 ( .A(n169), .Y(n960) );
  BUFX2 U45 ( .A(n187), .Y(n962) );
  BUFX2 U46 ( .A(n150), .Y(n959) );
  BUFX2 U47 ( .A(n150), .Y(n958) );
  BUFX2 U48 ( .A(n133), .Y(n956) );
  BUFX2 U81 ( .A(n133), .Y(n955) );
  BUFX2 U82 ( .A(n130), .Y(n953) );
  BUFX2 U115 ( .A(n130), .Y(n952) );
  BUFX2 U116 ( .A(n112), .Y(n950) );
  BUFX2 U149 ( .A(n112), .Y(n949) );
  BUFX2 U150 ( .A(n93), .Y(n947) );
  BUFX2 U183 ( .A(n93), .Y(n946) );
  BUFX2 U184 ( .A(n87), .Y(n944) );
  BUFX2 U217 ( .A(n87), .Y(n943) );
  BUFX2 U218 ( .A(n84), .Y(n941) );
  BUFX2 U251 ( .A(n84), .Y(n940) );
  BUFX2 U252 ( .A(n63), .Y(n929) );
  BUFX2 U285 ( .A(n63), .Y(n928) );
  INVX4 U286 ( .A(n992), .Y(n923) );
  INVX2 U319 ( .A(n923), .Y(n913) );
  INVX1 U320 ( .A(n50), .Y(n948) );
  INVX1 U353 ( .A(n51), .Y(n951) );
  INVX1 U354 ( .A(n53), .Y(n954) );
  INVX1 U387 ( .A(n54), .Y(n957) );
  INVX2 U388 ( .A(n995), .Y(n905) );
  INVX1 U421 ( .A(n34), .Y(n925) );
  INVX1 U422 ( .A(n45), .Y(n939) );
  INVX1 U455 ( .A(n56), .Y(n976) );
  INVX1 U456 ( .A(n57), .Y(n979) );
  INVX1 U457 ( .A(n47), .Y(n942) );
  INVX1 U490 ( .A(n48), .Y(n945) );
  BUFX2 U491 ( .A(n169), .Y(n961) );
  BUFX2 U524 ( .A(n205), .Y(n965) );
  BUFX2 U525 ( .A(n241), .Y(n969) );
  BUFX2 U558 ( .A(n262), .Y(n973) );
  BUFX2 U559 ( .A(n317), .Y(n983) );
  BUFX2 U560 ( .A(n354), .Y(n987) );
  INVX1 U563 ( .A(n33), .Y(n924) );
  INVX1 U564 ( .A(n35), .Y(n930) );
  INVX1 U567 ( .A(n36), .Y(n931) );
  INVX1 U568 ( .A(n37), .Y(n932) );
  INVX1 U571 ( .A(n38), .Y(n933) );
  INVX1 U572 ( .A(n39), .Y(n934) );
  INVX1 U575 ( .A(n40), .Y(n935) );
  INVX1 U576 ( .A(n41), .Y(n936) );
  INVX1 U579 ( .A(n43), .Y(n937) );
  INVX1 U580 ( .A(n44), .Y(n938) );
  INVX1 U583 ( .A(N22), .Y(n996) );
  AND2X1 U584 ( .A(n33), .B(n926), .Y(n1) );
  INVX1 U587 ( .A(n1), .Y(n2) );
  AND2X1 U588 ( .A(n35), .B(n926), .Y(n3) );
  INVX1 U591 ( .A(n3), .Y(n4) );
  AND2X1 U592 ( .A(n36), .B(n926), .Y(n5) );
  INVX1 U595 ( .A(n5), .Y(n6) );
  AND2X1 U596 ( .A(n37), .B(n926), .Y(n7) );
  INVX1 U599 ( .A(n7), .Y(n8) );
  AND2X1 U600 ( .A(n38), .B(n926), .Y(n9) );
  INVX1 U603 ( .A(n9), .Y(n10) );
  AND2X1 U604 ( .A(n39), .B(n926), .Y(n11) );
  INVX1 U607 ( .A(n11), .Y(n12) );
  AND2X1 U608 ( .A(n40), .B(n926), .Y(n13) );
  INVX1 U609 ( .A(n13), .Y(n14) );
  AND2X1 U612 ( .A(n41), .B(n926), .Y(n15) );
  INVX1 U613 ( .A(n15), .Y(n16) );
  AND2X1 U616 ( .A(n65), .B(n927), .Y(n17) );
  INVX1 U617 ( .A(n17), .Y(n18) );
  AND2X1 U620 ( .A(n68), .B(n927), .Y(n19) );
  INVX1 U621 ( .A(n19), .Y(n20) );
  AND2X1 U622 ( .A(n71), .B(n927), .Y(n21) );
  INVX1 U625 ( .A(n21), .Y(n22) );
  AND2X1 U626 ( .A(n74), .B(n927), .Y(n23) );
  INVX1 U627 ( .A(n23), .Y(n24) );
  AND2X1 U628 ( .A(n43), .B(n927), .Y(n25) );
  INVX1 U629 ( .A(n25), .Y(n26) );
  AND2X1 U630 ( .A(n44), .B(n927), .Y(n27) );
  INVX1 U631 ( .A(n27), .Y(n28) );
  AND2X1 U632 ( .A(n77), .B(n927), .Y(n29) );
  INVX1 U633 ( .A(n29), .Y(n30) );
  AND2X1 U635 ( .A(n80), .B(n927), .Y(n31) );
  INVX1 U636 ( .A(n31), .Y(n32) );
  AND2X1 U637 ( .A(n641), .B(n374), .Y(n33) );
  AND2X1 U638 ( .A(n643), .B(n635), .Y(n34) );
  AND2X1 U639 ( .A(n641), .B(n637), .Y(n35) );
  AND2X1 U640 ( .A(n641), .B(n358), .Y(n36) );
  AND2X1 U641 ( .A(n641), .B(n356), .Y(n37) );
  AND2X1 U642 ( .A(n645), .B(n374), .Y(n38) );
  AND2X1 U643 ( .A(n645), .B(n637), .Y(n39) );
  AND2X1 U644 ( .A(n645), .B(n358), .Y(n40) );
  AND2X1 U645 ( .A(n645), .B(n356), .Y(n41) );
  AND2X1 U646 ( .A(n374), .B(n355), .Y(n43) );
  AND2X1 U647 ( .A(n637), .B(n355), .Y(n44) );
  AND2X1 U648 ( .A(n643), .B(n639), .Y(n45) );
  AND2X1 U649 ( .A(n643), .B(n111), .Y(n47) );
  AND2X1 U650 ( .A(n643), .B(n92), .Y(n48) );
  AND2X1 U651 ( .A(n647), .B(n635), .Y(n50) );
  AND2X1 U652 ( .A(n647), .B(n639), .Y(n51) );
  AND2X1 U653 ( .A(n647), .B(n111), .Y(n53) );
  AND2X1 U654 ( .A(n647), .B(n92), .Y(n54) );
  AND2X1 U655 ( .A(n635), .B(n91), .Y(n56) );
  AND2X1 U656 ( .A(n639), .B(n91), .Y(n57) );
  OR2X1 U657 ( .A(n997), .B(rst), .Y(n59) );
  INVX1 U658 ( .A(n59), .Y(n60) );
  AND2X1 U659 ( .A(n34), .B(n990), .Y(n62) );
  INVX1 U660 ( .A(n62), .Y(n63) );
  AND2X1 U661 ( .A(n364), .B(n374), .Y(n65) );
  INVX1 U662 ( .A(n65), .Y(n66) );
  AND2X1 U663 ( .A(n364), .B(n637), .Y(n68) );
  INVX1 U664 ( .A(n68), .Y(n69) );
  AND2X1 U665 ( .A(n364), .B(n358), .Y(n71) );
  INVX1 U666 ( .A(n71), .Y(n72) );
  AND2X1 U667 ( .A(n364), .B(n356), .Y(n74) );
  INVX1 U668 ( .A(n74), .Y(n75) );
  AND2X1 U669 ( .A(n358), .B(n355), .Y(n77) );
  INVX1 U670 ( .A(n77), .Y(n78) );
  AND2X1 U671 ( .A(n355), .B(n356), .Y(n80) );
  INVX1 U672 ( .A(n80), .Y(n81) );
  AND2X1 U673 ( .A(n45), .B(n990), .Y(n83) );
  INVX1 U674 ( .A(n83), .Y(n84) );
  AND2X1 U675 ( .A(n47), .B(n990), .Y(n86) );
  INVX1 U676 ( .A(n86), .Y(n87) );
  AND2X1 U677 ( .A(n48), .B(n990), .Y(n89) );
  INVX1 U678 ( .A(n89), .Y(n93) );
  AND2X1 U679 ( .A(n50), .B(n990), .Y(n95) );
  INVX1 U680 ( .A(n95), .Y(n112) );
  AND2X1 U681 ( .A(n51), .B(n990), .Y(n114) );
  INVX1 U682 ( .A(n114), .Y(n130) );
  AND2X1 U683 ( .A(n53), .B(n990), .Y(n131) );
  INVX1 U684 ( .A(n131), .Y(n133) );
  AND2X1 U685 ( .A(n54), .B(n991), .Y(n149) );
  INVX1 U686 ( .A(n149), .Y(n150) );
  AND2X1 U687 ( .A(n168), .B(n635), .Y(n152) );
  INVX1 U688 ( .A(n152), .Y(n169) );
  AND2X1 U689 ( .A(n152), .B(n991), .Y(n171) );
  INVX1 U690 ( .A(n171), .Y(n187) );
  AND2X1 U691 ( .A(n168), .B(n639), .Y(n189) );
  INVX1 U692 ( .A(n189), .Y(n205) );
  AND2X1 U693 ( .A(n189), .B(n991), .Y(n207) );
  INVX1 U694 ( .A(n207), .Y(n223) );
  AND2X1 U695 ( .A(n168), .B(n111), .Y(n225) );
  INVX1 U696 ( .A(n225), .Y(n241) );
  AND2X1 U697 ( .A(n225), .B(n991), .Y(n242) );
  INVX1 U698 ( .A(n242), .Y(n244) );
  AND2X1 U699 ( .A(n168), .B(n92), .Y(n260) );
  INVX1 U700 ( .A(n260), .Y(n262) );
  AND2X1 U701 ( .A(n260), .B(n991), .Y(n278) );
  INVX1 U702 ( .A(n278), .Y(n280) );
  AND2X1 U703 ( .A(n56), .B(n991), .Y(n296) );
  INVX1 U704 ( .A(n296), .Y(n298) );
  AND2X1 U705 ( .A(n57), .B(n991), .Y(n314) );
  INVX1 U706 ( .A(n314), .Y(n315) );
  INVX1 U707 ( .A(n333), .Y(n317) );
  AND2X1 U708 ( .A(n111), .B(n91), .Y(n333) );
  AND2X1 U709 ( .A(n333), .B(n991), .Y(n335) );
  INVX1 U710 ( .A(n335), .Y(n351) );
  AND2X1 U711 ( .A(n91), .B(n92), .Y(n353) );
  INVX1 U712 ( .A(n353), .Y(n354) );
  AND2X1 U713 ( .A(n990), .B(n353), .Y(n360) );
  INVX1 U714 ( .A(n360), .Y(n362) );
  OR2X1 U715 ( .A(n915), .B(n993), .Y(n369) );
  INVX1 U716 ( .A(n369), .Y(n374) );
  OR2X1 U717 ( .A(N22), .B(N23), .Y(n634) );
  INVX1 U718 ( .A(n634), .Y(n635) );
  OR2X1 U719 ( .A(n992), .B(n993), .Y(n636) );
  INVX1 U720 ( .A(n636), .Y(n637) );
  OR2X1 U721 ( .A(n996), .B(N23), .Y(n638) );
  INVX1 U722 ( .A(n638), .Y(n639) );
  OR2X1 U723 ( .A(n905), .B(N21), .Y(n640) );
  INVX1 U724 ( .A(n640), .Y(n641) );
  OR2X1 U725 ( .A(N24), .B(N25), .Y(n642) );
  INVX1 U726 ( .A(n642), .Y(n643) );
  OR2X1 U727 ( .A(n995), .B(N21), .Y(n644) );
  INVX1 U728 ( .A(n644), .Y(n645) );
  OR2X1 U729 ( .A(n999), .B(N25), .Y(n646) );
  INVX1 U730 ( .A(n646), .Y(n647) );
  MUX2X1 U731 ( .B(n649), .A(n650), .S(n912), .Y(n648) );
  MUX2X1 U732 ( .B(n652), .A(n653), .S(n912), .Y(n651) );
  MUX2X1 U733 ( .B(n655), .A(n656), .S(n912), .Y(n654) );
  MUX2X1 U734 ( .B(n658), .A(n659), .S(n912), .Y(n657) );
  MUX2X1 U735 ( .B(n661), .A(n662), .S(n904), .Y(n660) );
  MUX2X1 U736 ( .B(n664), .A(n665), .S(n912), .Y(n663) );
  MUX2X1 U737 ( .B(n667), .A(n668), .S(n912), .Y(n666) );
  MUX2X1 U738 ( .B(n670), .A(n671), .S(n912), .Y(n669) );
  MUX2X1 U739 ( .B(n673), .A(n674), .S(n912), .Y(n672) );
  MUX2X1 U740 ( .B(n676), .A(n677), .S(n904), .Y(n675) );
  MUX2X1 U741 ( .B(n679), .A(n680), .S(n912), .Y(n678) );
  MUX2X1 U742 ( .B(n682), .A(n683), .S(n912), .Y(n681) );
  MUX2X1 U743 ( .B(n685), .A(n686), .S(n912), .Y(n684) );
  MUX2X1 U744 ( .B(n688), .A(n689), .S(n912), .Y(n687) );
  MUX2X1 U745 ( .B(n691), .A(n692), .S(n904), .Y(n690) );
  MUX2X1 U746 ( .B(n694), .A(n695), .S(n911), .Y(n693) );
  MUX2X1 U747 ( .B(n697), .A(n698), .S(n911), .Y(n696) );
  MUX2X1 U748 ( .B(n700), .A(n701), .S(n911), .Y(n699) );
  MUX2X1 U749 ( .B(n703), .A(n704), .S(n911), .Y(n702) );
  MUX2X1 U750 ( .B(n706), .A(n707), .S(n904), .Y(n705) );
  MUX2X1 U751 ( .B(n709), .A(n710), .S(N23), .Y(n708) );
  MUX2X1 U752 ( .B(n712), .A(n713), .S(n911), .Y(n711) );
  MUX2X1 U753 ( .B(n715), .A(n716), .S(n911), .Y(n714) );
  MUX2X1 U754 ( .B(n718), .A(n719), .S(n911), .Y(n717) );
  MUX2X1 U755 ( .B(n721), .A(n722), .S(n911), .Y(n720) );
  MUX2X1 U756 ( .B(n724), .A(n725), .S(n904), .Y(n723) );
  MUX2X1 U757 ( .B(n727), .A(n728), .S(n911), .Y(n726) );
  MUX2X1 U758 ( .B(n730), .A(n731), .S(n911), .Y(n729) );
  MUX2X1 U759 ( .B(n733), .A(n734), .S(n911), .Y(n732) );
  MUX2X1 U760 ( .B(n736), .A(n737), .S(n911), .Y(n735) );
  MUX2X1 U761 ( .B(n739), .A(n740), .S(n904), .Y(n738) );
  MUX2X1 U762 ( .B(n742), .A(n743), .S(n910), .Y(n741) );
  MUX2X1 U763 ( .B(n745), .A(n746), .S(n910), .Y(n744) );
  MUX2X1 U764 ( .B(n748), .A(n749), .S(n910), .Y(n747) );
  MUX2X1 U765 ( .B(n751), .A(n752), .S(n910), .Y(n750) );
  MUX2X1 U766 ( .B(n754), .A(n755), .S(n904), .Y(n753) );
  MUX2X1 U767 ( .B(n757), .A(n758), .S(n910), .Y(n756) );
  MUX2X1 U768 ( .B(n760), .A(n761), .S(n910), .Y(n759) );
  MUX2X1 U769 ( .B(n763), .A(n764), .S(n910), .Y(n762) );
  MUX2X1 U770 ( .B(n766), .A(n767), .S(n910), .Y(n765) );
  MUX2X1 U771 ( .B(n769), .A(n770), .S(n904), .Y(n768) );
  MUX2X1 U772 ( .B(n772), .A(n773), .S(N23), .Y(n771) );
  MUX2X1 U773 ( .B(n775), .A(n776), .S(n910), .Y(n774) );
  MUX2X1 U774 ( .B(n778), .A(n779), .S(n910), .Y(n777) );
  MUX2X1 U775 ( .B(n781), .A(n782), .S(n910), .Y(n780) );
  MUX2X1 U776 ( .B(n784), .A(n785), .S(n910), .Y(n783) );
  MUX2X1 U777 ( .B(n787), .A(n788), .S(n904), .Y(n786) );
  MUX2X1 U778 ( .B(n790), .A(n791), .S(n910), .Y(n789) );
  MUX2X1 U779 ( .B(n793), .A(n794), .S(n911), .Y(n792) );
  MUX2X1 U780 ( .B(n796), .A(n797), .S(n912), .Y(n795) );
  MUX2X1 U781 ( .B(n799), .A(n800), .S(n912), .Y(n798) );
  MUX2X1 U782 ( .B(n802), .A(n803), .S(n904), .Y(n801) );
  MUX2X1 U783 ( .B(n805), .A(n806), .S(n912), .Y(n804) );
  MUX2X1 U784 ( .B(n808), .A(n809), .S(n911), .Y(n807) );
  MUX2X1 U785 ( .B(n811), .A(n812), .S(n909), .Y(n810) );
  MUX2X1 U786 ( .B(n814), .A(n815), .S(n909), .Y(n813) );
  MUX2X1 U787 ( .B(n817), .A(n818), .S(n904), .Y(n816) );
  MUX2X1 U788 ( .B(n820), .A(n821), .S(n911), .Y(n819) );
  MUX2X1 U789 ( .B(n823), .A(n824), .S(n911), .Y(n822) );
  MUX2X1 U790 ( .B(n826), .A(n827), .S(n909), .Y(n825) );
  MUX2X1 U791 ( .B(n829), .A(n830), .S(n910), .Y(n828) );
  MUX2X1 U792 ( .B(n832), .A(n833), .S(n904), .Y(n831) );
  MUX2X1 U793 ( .B(n835), .A(n836), .S(N23), .Y(n834) );
  MUX2X1 U794 ( .B(n838), .A(n839), .S(n909), .Y(n837) );
  MUX2X1 U795 ( .B(n841), .A(n842), .S(n911), .Y(n840) );
  MUX2X1 U796 ( .B(n844), .A(n845), .S(n911), .Y(n843) );
  MUX2X1 U797 ( .B(n847), .A(n848), .S(n911), .Y(n846) );
  MUX2X1 U798 ( .B(n850), .A(n851), .S(n903), .Y(n849) );
  MUX2X1 U799 ( .B(n853), .A(n854), .S(n912), .Y(n852) );
  MUX2X1 U800 ( .B(n856), .A(n857), .S(n910), .Y(n855) );
  MUX2X1 U801 ( .B(n859), .A(n860), .S(n912), .Y(n858) );
  MUX2X1 U802 ( .B(n862), .A(n863), .S(n910), .Y(n861) );
  MUX2X1 U803 ( .B(n865), .A(n866), .S(n903), .Y(n864) );
  MUX2X1 U804 ( .B(n868), .A(n869), .S(n909), .Y(n867) );
  MUX2X1 U805 ( .B(n871), .A(n872), .S(n909), .Y(n870) );
  MUX2X1 U806 ( .B(n874), .A(n875), .S(n909), .Y(n873) );
  MUX2X1 U807 ( .B(n877), .A(n878), .S(n909), .Y(n876) );
  MUX2X1 U808 ( .B(n880), .A(n881), .S(n903), .Y(n879) );
  MUX2X1 U809 ( .B(n883), .A(n884), .S(n909), .Y(n882) );
  MUX2X1 U810 ( .B(n886), .A(n887), .S(n909), .Y(n885) );
  MUX2X1 U811 ( .B(n889), .A(n890), .S(n909), .Y(n888) );
  MUX2X1 U812 ( .B(n892), .A(n893), .S(n909), .Y(n891) );
  MUX2X1 U813 ( .B(n895), .A(n896), .S(n903), .Y(n894) );
  MUX2X1 U814 ( .B(n898), .A(n899), .S(N23), .Y(n897) );
  MUX2X1 U815 ( .B(n900), .A(n901), .S(N25), .Y(N28) );
  MUX2X1 U816 ( .B(\mem<254> ), .A(\mem<255> ), .S(n915), .Y(n650) );
  MUX2X1 U817 ( .B(\mem<252> ), .A(\mem<253> ), .S(n915), .Y(n649) );
  MUX2X1 U818 ( .B(\mem<250> ), .A(\mem<251> ), .S(n915), .Y(n653) );
  MUX2X1 U819 ( .B(\mem<248> ), .A(\mem<249> ), .S(n915), .Y(n652) );
  MUX2X1 U820 ( .B(n651), .A(n648), .S(n907), .Y(n662) );
  MUX2X1 U821 ( .B(\mem<246> ), .A(\mem<247> ), .S(n915), .Y(n656) );
  MUX2X1 U822 ( .B(\mem<244> ), .A(\mem<245> ), .S(n915), .Y(n655) );
  MUX2X1 U823 ( .B(\mem<242> ), .A(\mem<243> ), .S(n915), .Y(n659) );
  MUX2X1 U824 ( .B(\mem<240> ), .A(\mem<241> ), .S(n915), .Y(n658) );
  MUX2X1 U825 ( .B(n657), .A(n654), .S(n907), .Y(n661) );
  MUX2X1 U826 ( .B(\mem<238> ), .A(\mem<239> ), .S(n916), .Y(n665) );
  MUX2X1 U827 ( .B(\mem<236> ), .A(\mem<237> ), .S(n916), .Y(n664) );
  MUX2X1 U828 ( .B(\mem<234> ), .A(\mem<235> ), .S(n916), .Y(n668) );
  MUX2X1 U829 ( .B(\mem<232> ), .A(\mem<233> ), .S(n916), .Y(n667) );
  MUX2X1 U830 ( .B(n666), .A(n663), .S(n907), .Y(n677) );
  MUX2X1 U831 ( .B(\mem<230> ), .A(\mem<231> ), .S(n916), .Y(n671) );
  MUX2X1 U832 ( .B(\mem<228> ), .A(\mem<229> ), .S(n916), .Y(n670) );
  MUX2X1 U833 ( .B(\mem<226> ), .A(\mem<227> ), .S(n916), .Y(n674) );
  MUX2X1 U834 ( .B(\mem<224> ), .A(\mem<225> ), .S(n916), .Y(n673) );
  MUX2X1 U835 ( .B(n672), .A(n669), .S(n907), .Y(n676) );
  MUX2X1 U836 ( .B(n675), .A(n660), .S(N22), .Y(n710) );
  MUX2X1 U837 ( .B(\mem<222> ), .A(\mem<223> ), .S(n916), .Y(n680) );
  MUX2X1 U838 ( .B(\mem<220> ), .A(\mem<221> ), .S(n916), .Y(n679) );
  MUX2X1 U839 ( .B(\mem<218> ), .A(\mem<219> ), .S(n916), .Y(n683) );
  MUX2X1 U840 ( .B(\mem<216> ), .A(\mem<217> ), .S(n916), .Y(n682) );
  MUX2X1 U841 ( .B(n681), .A(n678), .S(n907), .Y(n692) );
  MUX2X1 U842 ( .B(\mem<214> ), .A(\mem<215> ), .S(n917), .Y(n686) );
  MUX2X1 U843 ( .B(\mem<212> ), .A(\mem<213> ), .S(n917), .Y(n685) );
  MUX2X1 U844 ( .B(\mem<210> ), .A(\mem<211> ), .S(n917), .Y(n689) );
  MUX2X1 U845 ( .B(\mem<208> ), .A(\mem<209> ), .S(n917), .Y(n688) );
  MUX2X1 U846 ( .B(n687), .A(n684), .S(n907), .Y(n691) );
  MUX2X1 U847 ( .B(\mem<206> ), .A(\mem<207> ), .S(n917), .Y(n695) );
  MUX2X1 U848 ( .B(\mem<204> ), .A(\mem<205> ), .S(n917), .Y(n694) );
  MUX2X1 U849 ( .B(\mem<202> ), .A(\mem<203> ), .S(n917), .Y(n698) );
  MUX2X1 U850 ( .B(\mem<200> ), .A(\mem<201> ), .S(n917), .Y(n697) );
  MUX2X1 U851 ( .B(n696), .A(n693), .S(n907), .Y(n707) );
  MUX2X1 U852 ( .B(\mem<198> ), .A(\mem<199> ), .S(n917), .Y(n701) );
  MUX2X1 U853 ( .B(\mem<196> ), .A(\mem<197> ), .S(n917), .Y(n700) );
  MUX2X1 U854 ( .B(\mem<194> ), .A(\mem<195> ), .S(n917), .Y(n704) );
  MUX2X1 U855 ( .B(\mem<192> ), .A(\mem<193> ), .S(n917), .Y(n703) );
  MUX2X1 U856 ( .B(n702), .A(n699), .S(n907), .Y(n706) );
  MUX2X1 U857 ( .B(n705), .A(n690), .S(N22), .Y(n709) );
  MUX2X1 U858 ( .B(\mem<190> ), .A(\mem<191> ), .S(n918), .Y(n713) );
  MUX2X1 U859 ( .B(\mem<188> ), .A(\mem<189> ), .S(n918), .Y(n712) );
  MUX2X1 U860 ( .B(\mem<186> ), .A(\mem<187> ), .S(n918), .Y(n716) );
  MUX2X1 U861 ( .B(\mem<184> ), .A(\mem<185> ), .S(n918), .Y(n715) );
  MUX2X1 U862 ( .B(n714), .A(n711), .S(n907), .Y(n725) );
  MUX2X1 U863 ( .B(\mem<182> ), .A(\mem<183> ), .S(n918), .Y(n719) );
  MUX2X1 U864 ( .B(\mem<180> ), .A(\mem<181> ), .S(n918), .Y(n718) );
  MUX2X1 U865 ( .B(\mem<178> ), .A(\mem<179> ), .S(n918), .Y(n722) );
  MUX2X1 U866 ( .B(\mem<176> ), .A(\mem<177> ), .S(n918), .Y(n721) );
  MUX2X1 U867 ( .B(n720), .A(n717), .S(n907), .Y(n724) );
  MUX2X1 U868 ( .B(\mem<174> ), .A(\mem<175> ), .S(n918), .Y(n728) );
  MUX2X1 U869 ( .B(\mem<172> ), .A(\mem<173> ), .S(n918), .Y(n727) );
  MUX2X1 U870 ( .B(\mem<170> ), .A(\mem<171> ), .S(n918), .Y(n731) );
  MUX2X1 U871 ( .B(\mem<168> ), .A(\mem<169> ), .S(n918), .Y(n730) );
  MUX2X1 U872 ( .B(n729), .A(n726), .S(n907), .Y(n740) );
  MUX2X1 U873 ( .B(\mem<166> ), .A(\mem<167> ), .S(n917), .Y(n734) );
  MUX2X1 U874 ( .B(\mem<164> ), .A(\mem<165> ), .S(n918), .Y(n733) );
  MUX2X1 U875 ( .B(\mem<162> ), .A(\mem<163> ), .S(n920), .Y(n737) );
  MUX2X1 U876 ( .B(\mem<160> ), .A(\mem<161> ), .S(n915), .Y(n736) );
  MUX2X1 U877 ( .B(n735), .A(n732), .S(n907), .Y(n739) );
  MUX2X1 U878 ( .B(n738), .A(n723), .S(N22), .Y(n773) );
  MUX2X1 U879 ( .B(\mem<158> ), .A(\mem<159> ), .S(n918), .Y(n743) );
  MUX2X1 U880 ( .B(\mem<156> ), .A(\mem<157> ), .S(n917), .Y(n742) );
  MUX2X1 U881 ( .B(\mem<154> ), .A(\mem<155> ), .S(n916), .Y(n746) );
  MUX2X1 U882 ( .B(\mem<152> ), .A(\mem<153> ), .S(n921), .Y(n745) );
  MUX2X1 U883 ( .B(n744), .A(n741), .S(n906), .Y(n755) );
  MUX2X1 U884 ( .B(\mem<150> ), .A(\mem<151> ), .S(n915), .Y(n749) );
  MUX2X1 U885 ( .B(\mem<148> ), .A(\mem<149> ), .S(n916), .Y(n748) );
  MUX2X1 U886 ( .B(\mem<146> ), .A(\mem<147> ), .S(n916), .Y(n752) );
  MUX2X1 U887 ( .B(\mem<144> ), .A(\mem<145> ), .S(n917), .Y(n751) );
  MUX2X1 U888 ( .B(n750), .A(n747), .S(n906), .Y(n754) );
  MUX2X1 U889 ( .B(\mem<142> ), .A(\mem<143> ), .S(n917), .Y(n758) );
  MUX2X1 U890 ( .B(\mem<140> ), .A(\mem<141> ), .S(n918), .Y(n757) );
  MUX2X1 U891 ( .B(\mem<138> ), .A(\mem<139> ), .S(n918), .Y(n761) );
  MUX2X1 U892 ( .B(\mem<136> ), .A(\mem<137> ), .S(n917), .Y(n760) );
  MUX2X1 U893 ( .B(n759), .A(n756), .S(n906), .Y(n770) );
  MUX2X1 U894 ( .B(\mem<134> ), .A(\mem<135> ), .S(n915), .Y(n764) );
  MUX2X1 U895 ( .B(\mem<132> ), .A(\mem<133> ), .S(n918), .Y(n763) );
  MUX2X1 U896 ( .B(\mem<130> ), .A(\mem<131> ), .S(n918), .Y(n767) );
  MUX2X1 U897 ( .B(\mem<128> ), .A(\mem<129> ), .S(n915), .Y(n766) );
  MUX2X1 U898 ( .B(n765), .A(n762), .S(n906), .Y(n769) );
  MUX2X1 U899 ( .B(n768), .A(n753), .S(N22), .Y(n772) );
  MUX2X1 U900 ( .B(n771), .A(n708), .S(N24), .Y(n901) );
  MUX2X1 U901 ( .B(\mem<126> ), .A(\mem<127> ), .S(n915), .Y(n776) );
  MUX2X1 U902 ( .B(\mem<124> ), .A(\mem<125> ), .S(n918), .Y(n775) );
  MUX2X1 U903 ( .B(\mem<122> ), .A(\mem<123> ), .S(n921), .Y(n779) );
  MUX2X1 U904 ( .B(\mem<120> ), .A(\mem<121> ), .S(n916), .Y(n778) );
  MUX2X1 U905 ( .B(n777), .A(n774), .S(n906), .Y(n788) );
  MUX2X1 U906 ( .B(\mem<118> ), .A(\mem<119> ), .S(n919), .Y(n782) );
  MUX2X1 U907 ( .B(\mem<116> ), .A(\mem<117> ), .S(n919), .Y(n781) );
  MUX2X1 U908 ( .B(\mem<114> ), .A(\mem<115> ), .S(n919), .Y(n785) );
  MUX2X1 U909 ( .B(\mem<112> ), .A(\mem<113> ), .S(n919), .Y(n784) );
  MUX2X1 U910 ( .B(n783), .A(n780), .S(n906), .Y(n787) );
  MUX2X1 U911 ( .B(\mem<110> ), .A(\mem<111> ), .S(n919), .Y(n791) );
  MUX2X1 U912 ( .B(\mem<108> ), .A(\mem<109> ), .S(n919), .Y(n790) );
  MUX2X1 U913 ( .B(\mem<106> ), .A(\mem<107> ), .S(n919), .Y(n794) );
  MUX2X1 U914 ( .B(\mem<104> ), .A(\mem<105> ), .S(n919), .Y(n793) );
  MUX2X1 U915 ( .B(n792), .A(n789), .S(n906), .Y(n803) );
  MUX2X1 U916 ( .B(\mem<102> ), .A(\mem<103> ), .S(n919), .Y(n797) );
  MUX2X1 U917 ( .B(\mem<100> ), .A(\mem<101> ), .S(n919), .Y(n796) );
  MUX2X1 U918 ( .B(\mem<98> ), .A(\mem<99> ), .S(n919), .Y(n800) );
  MUX2X1 U919 ( .B(\mem<96> ), .A(\mem<97> ), .S(n919), .Y(n799) );
  MUX2X1 U920 ( .B(n798), .A(n795), .S(n906), .Y(n802) );
  MUX2X1 U921 ( .B(n801), .A(n786), .S(N22), .Y(n836) );
  MUX2X1 U922 ( .B(\mem<94> ), .A(\mem<95> ), .S(n920), .Y(n806) );
  MUX2X1 U923 ( .B(\mem<92> ), .A(\mem<93> ), .S(n920), .Y(n805) );
  MUX2X1 U924 ( .B(\mem<90> ), .A(\mem<91> ), .S(n920), .Y(n809) );
  MUX2X1 U925 ( .B(\mem<88> ), .A(\mem<89> ), .S(n920), .Y(n808) );
  MUX2X1 U926 ( .B(n807), .A(n804), .S(n906), .Y(n818) );
  MUX2X1 U927 ( .B(\mem<86> ), .A(\mem<87> ), .S(n920), .Y(n812) );
  MUX2X1 U928 ( .B(\mem<84> ), .A(\mem<85> ), .S(n920), .Y(n811) );
  MUX2X1 U929 ( .B(\mem<82> ), .A(\mem<83> ), .S(n920), .Y(n815) );
  MUX2X1 U930 ( .B(\mem<80> ), .A(\mem<81> ), .S(n920), .Y(n814) );
  MUX2X1 U931 ( .B(n813), .A(n810), .S(n906), .Y(n817) );
  MUX2X1 U932 ( .B(\mem<78> ), .A(\mem<79> ), .S(n920), .Y(n821) );
  MUX2X1 U933 ( .B(\mem<76> ), .A(\mem<77> ), .S(n920), .Y(n820) );
  MUX2X1 U934 ( .B(\mem<74> ), .A(\mem<75> ), .S(n920), .Y(n824) );
  MUX2X1 U935 ( .B(\mem<72> ), .A(\mem<73> ), .S(n920), .Y(n823) );
  MUX2X1 U936 ( .B(n822), .A(n819), .S(n906), .Y(n833) );
  MUX2X1 U937 ( .B(\mem<70> ), .A(\mem<71> ), .S(n921), .Y(n827) );
  MUX2X1 U938 ( .B(\mem<68> ), .A(\mem<69> ), .S(n921), .Y(n826) );
  MUX2X1 U939 ( .B(\mem<66> ), .A(\mem<67> ), .S(n921), .Y(n830) );
  MUX2X1 U940 ( .B(\mem<64> ), .A(\mem<65> ), .S(n921), .Y(n829) );
  MUX2X1 U941 ( .B(n828), .A(n825), .S(n906), .Y(n832) );
  MUX2X1 U942 ( .B(n831), .A(n816), .S(N22), .Y(n835) );
  MUX2X1 U943 ( .B(\mem<62> ), .A(\mem<63> ), .S(n921), .Y(n839) );
  MUX2X1 U944 ( .B(\mem<60> ), .A(\mem<61> ), .S(n921), .Y(n838) );
  MUX2X1 U945 ( .B(\mem<58> ), .A(\mem<59> ), .S(n921), .Y(n842) );
  MUX2X1 U946 ( .B(\mem<56> ), .A(\mem<57> ), .S(n921), .Y(n841) );
  MUX2X1 U947 ( .B(n840), .A(n837), .S(n905), .Y(n851) );
  MUX2X1 U948 ( .B(\mem<54> ), .A(\mem<55> ), .S(n921), .Y(n845) );
  MUX2X1 U949 ( .B(\mem<52> ), .A(\mem<53> ), .S(n921), .Y(n844) );
  MUX2X1 U950 ( .B(\mem<50> ), .A(\mem<51> ), .S(n921), .Y(n848) );
  MUX2X1 U951 ( .B(\mem<48> ), .A(\mem<49> ), .S(n921), .Y(n847) );
  MUX2X1 U952 ( .B(n846), .A(n843), .S(n905), .Y(n850) );
  MUX2X1 U953 ( .B(\mem<46> ), .A(\mem<47> ), .S(n922), .Y(n854) );
  MUX2X1 U954 ( .B(\mem<44> ), .A(\mem<45> ), .S(n922), .Y(n853) );
  MUX2X1 U955 ( .B(\mem<42> ), .A(\mem<43> ), .S(n922), .Y(n857) );
  MUX2X1 U956 ( .B(\mem<40> ), .A(\mem<41> ), .S(n922), .Y(n856) );
  MUX2X1 U957 ( .B(n855), .A(n852), .S(n905), .Y(n866) );
  MUX2X1 U958 ( .B(\mem<38> ), .A(\mem<39> ), .S(n922), .Y(n860) );
  MUX2X1 U959 ( .B(\mem<36> ), .A(\mem<37> ), .S(n922), .Y(n859) );
  MUX2X1 U960 ( .B(\mem<34> ), .A(\mem<35> ), .S(n922), .Y(n863) );
  MUX2X1 U961 ( .B(\mem<32> ), .A(\mem<33> ), .S(n922), .Y(n862) );
  MUX2X1 U962 ( .B(n861), .A(n858), .S(n905), .Y(n865) );
  MUX2X1 U963 ( .B(n864), .A(n849), .S(N22), .Y(n899) );
  MUX2X1 U964 ( .B(\mem<30> ), .A(\mem<31> ), .S(n922), .Y(n869) );
  MUX2X1 U965 ( .B(\mem<28> ), .A(\mem<29> ), .S(n922), .Y(n868) );
  MUX2X1 U966 ( .B(\mem<26> ), .A(\mem<27> ), .S(n922), .Y(n872) );
  MUX2X1 U967 ( .B(\mem<24> ), .A(\mem<25> ), .S(n922), .Y(n871) );
  MUX2X1 U968 ( .B(n870), .A(n867), .S(n905), .Y(n881) );
  MUX2X1 U969 ( .B(\mem<22> ), .A(\mem<23> ), .S(n916), .Y(n875) );
  MUX2X1 U970 ( .B(\mem<20> ), .A(\mem<21> ), .S(n923), .Y(n874) );
  MUX2X1 U971 ( .B(\mem<18> ), .A(\mem<19> ), .S(n915), .Y(n878) );
  MUX2X1 U972 ( .B(\mem<16> ), .A(\mem<17> ), .S(n919), .Y(n877) );
  MUX2X1 U973 ( .B(n876), .A(n873), .S(n905), .Y(n880) );
  MUX2X1 U974 ( .B(\mem<14> ), .A(\mem<15> ), .S(n918), .Y(n884) );
  MUX2X1 U975 ( .B(\mem<12> ), .A(\mem<13> ), .S(n916), .Y(n883) );
  MUX2X1 U976 ( .B(\mem<10> ), .A(\mem<11> ), .S(n923), .Y(n887) );
  MUX2X1 U977 ( .B(\mem<8> ), .A(\mem<9> ), .S(n916), .Y(n886) );
  MUX2X1 U978 ( .B(n885), .A(n882), .S(n905), .Y(n896) );
  MUX2X1 U979 ( .B(\mem<6> ), .A(\mem<7> ), .S(n915), .Y(n890) );
  MUX2X1 U980 ( .B(\mem<4> ), .A(\mem<5> ), .S(n922), .Y(n889) );
  MUX2X1 U981 ( .B(\mem<2> ), .A(\mem<3> ), .S(n917), .Y(n893) );
  MUX2X1 U982 ( .B(\mem<0> ), .A(\mem<1> ), .S(n915), .Y(n892) );
  MUX2X1 U983 ( .B(n891), .A(n888), .S(n905), .Y(n895) );
  MUX2X1 U984 ( .B(n894), .A(n879), .S(N22), .Y(n898) );
  MUX2X1 U985 ( .B(n897), .A(n834), .S(N24), .Y(n900) );
  INVX8 U986 ( .A(n908), .Y(n909) );
  INVX8 U987 ( .A(n908), .Y(n910) );
  INVX8 U988 ( .A(n908), .Y(n911) );
  INVX8 U989 ( .A(n908), .Y(n912) );
  INVX8 U990 ( .A(n923), .Y(n914) );
  INVX8 U991 ( .A(n914), .Y(n915) );
  INVX8 U992 ( .A(n914), .Y(n916) );
  INVX8 U993 ( .A(n914), .Y(n917) );
  INVX8 U994 ( .A(n914), .Y(n918) );
  INVX8 U995 ( .A(n913), .Y(n919) );
  INVX8 U996 ( .A(n914), .Y(n920) );
  INVX8 U997 ( .A(n914), .Y(n921) );
  INVX8 U998 ( .A(n913), .Y(n922) );
  INVX1 U999 ( .A(N20), .Y(n995) );
  INVX1 U1000 ( .A(N19), .Y(n994) );
  INVX1 U1001 ( .A(write), .Y(n997) );
  INVX1 U1002 ( .A(N18), .Y(n992) );
endmodule


module final_memory_3 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1050, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n373, n374, n375, n376, n377, n378, n380,
         n382, n383, n384, n385, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n403, n404, n405, n406, n407,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n584, n585, n586, n587,
         n588, n589, n590, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n50, n150, n189, n289, n348, n372, n379, n381, n386, n387,
         n401, n402, n409, n421, n422, n434, n435, n447, n448, n460, n461,
         n473, n474, n486, n487, n507, n508, n522, n523, n537, n538, n552,
         n553, n567, n568, n582, n583, n591, n592, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n870), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n869), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n868), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n867), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n866), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n865), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n864), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n863), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n862), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n861), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n860), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n859), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n858), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n857), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n856), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n855), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n854), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n853), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n852), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n851), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n850), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n849), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n848), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n847), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n846), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n845), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n844), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n843), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n842), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n841), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n840), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n839), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n838), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n837), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n836), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n835), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n834), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n833), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n832), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n831), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n830), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n829), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n828), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n827), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n826), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n825), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n824), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n823), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n822), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n821), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n820), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n819), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n818), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n817), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n816), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n815), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n814), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n813), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n812), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n811), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n810), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n809), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n808), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n807), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n806), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n805), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n804), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n803), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n802), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n801), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n800), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n799), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n798), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n797), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n796), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n795), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n794), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n793), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n792), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n791), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n790), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n789), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n788), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n787), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n786), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n785), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n784), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n783), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n782), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n781), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n780), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n779), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n778), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n777), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n776), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n775), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n774), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n773), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n772), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n771), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n770), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n769), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n768), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n767), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n766), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n765), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n764), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n763), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n762), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n761), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n760), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n759), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n758), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n757), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n756), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n755), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n754), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n753), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n752), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n751), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n750), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n749), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n748), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n747), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n746), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n745), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n744), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n743), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n742), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n741), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n740), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n739), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n738), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n737), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n736), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n735), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n734), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n733), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n732), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n731), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n730), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n729), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n728), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n727), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n726), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n725), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n724), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n723), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n722), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n721), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n720), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n719), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n718), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n717), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n716), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n715), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n714), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n713), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n712), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n711), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n710), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n709), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n708), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n707), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n706), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n705), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n704), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n703), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n702), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n701), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n700), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n699), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n698), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n697), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n696), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n695), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n694), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n693), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n692), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n691), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n690), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n689), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n688), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n687), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n686), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n685), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n684), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n683), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n682), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n681), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n680), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n679), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n678), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n677), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n676), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n675), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n674), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n673), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n672), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n671), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n670), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n669), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n668), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n667), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n666), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n665), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n664), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n663), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n662), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n661), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n660), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n659), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n658), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n657), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n656), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n655), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n654), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n653), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n652), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n651), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n650), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n649), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n648), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n647), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n646), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n645), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n644), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n643), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n642), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n641), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n640), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n639), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n638), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n637), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n636), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n635), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n634), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n633), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n632), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n631), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n630), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n629), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n628), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n627), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n626), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n625), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n624), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n623), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n622), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n621), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n620), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n619), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n618), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n617), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n616), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n615), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n614), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n613), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n612), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n611), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n610), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n609), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n608), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n607), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n413), .B(n414), .Y(n412) );
  AND2X2 U10 ( .A(n418), .B(n419), .Y(n417) );
  AND2X2 U11 ( .A(n426), .B(n427), .Y(n425) );
  AND2X2 U12 ( .A(n431), .B(n432), .Y(n430) );
  AND2X2 U13 ( .A(n439), .B(n440), .Y(n438) );
  AND2X2 U14 ( .A(n444), .B(n445), .Y(n443) );
  AND2X2 U15 ( .A(n452), .B(n453), .Y(n451) );
  AND2X2 U16 ( .A(n457), .B(n458), .Y(n456) );
  AND2X2 U17 ( .A(n465), .B(n466), .Y(n464) );
  AND2X2 U18 ( .A(n470), .B(n471), .Y(n469) );
  AND2X2 U19 ( .A(n478), .B(n479), .Y(n477) );
  AND2X2 U20 ( .A(n483), .B(n484), .Y(n482) );
  AND2X2 U21 ( .A(n491), .B(n492), .Y(n490) );
  AND2X2 U22 ( .A(n496), .B(n497), .Y(n495) );
  AND2X2 U30 ( .A(n588), .B(n1030), .Y(n248) );
  AND2X2 U31 ( .A(n589), .B(n1030), .Y(n91) );
  AND2X2 U32 ( .A(n588), .B(\addr_1c<0> ), .Y(n228) );
  AND2X2 U33 ( .A(n589), .B(\addr_1c<0> ), .Y(n71) );
  AND2X2 U34 ( .A(n596), .B(n597), .Y(n595) );
  AND2X2 U45 ( .A(n603), .B(n604), .Y(n602) );
  NOR3X1 U94 ( .A(n1018), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1019), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1042), .C(n40), .Y(n607) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n40) );
  OAI21X1 U98 ( .A(n1011), .B(n1043), .C(n41), .Y(n608) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n41) );
  OAI21X1 U100 ( .A(n1011), .B(n1044), .C(n42), .Y(n609) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n42) );
  OAI21X1 U102 ( .A(n1011), .B(n1045), .C(n43), .Y(n610) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n43) );
  OAI21X1 U104 ( .A(n1011), .B(n1046), .C(n44), .Y(n611) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n44) );
  OAI21X1 U106 ( .A(n1011), .B(n1047), .C(n45), .Y(n612) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n45) );
  OAI21X1 U108 ( .A(n1011), .B(n1048), .C(n46), .Y(n613) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n46) );
  OAI21X1 U110 ( .A(n1011), .B(n1049), .C(n47), .Y(n614) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n47) );
  NAND3X1 U112 ( .A(n1012), .B(n49), .C(n965), .Y(n39) );
  OAI21X1 U113 ( .A(n6), .B(n1034), .C(n51), .Y(n615) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n51) );
  OAI21X1 U115 ( .A(n6), .B(n1035), .C(n52), .Y(n616) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n52) );
  OAI21X1 U117 ( .A(n6), .B(n1036), .C(n53), .Y(n617) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n53) );
  OAI21X1 U119 ( .A(n6), .B(n1037), .C(n54), .Y(n618) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n54) );
  OAI21X1 U121 ( .A(n6), .B(n1038), .C(n55), .Y(n619) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n55) );
  OAI21X1 U123 ( .A(n6), .B(n1039), .C(n56), .Y(n620) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n56) );
  OAI21X1 U125 ( .A(n6), .B(n1040), .C(n57), .Y(n621) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n57) );
  OAI21X1 U127 ( .A(n6), .B(n1041), .C(n58), .Y(n622) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n58) );
  OAI21X1 U130 ( .A(n1042), .B(n1010), .C(n62), .Y(n623) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n62) );
  OAI21X1 U132 ( .A(n1043), .B(n1009), .C(n63), .Y(n624) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n63) );
  OAI21X1 U134 ( .A(n1044), .B(n1009), .C(n64), .Y(n625) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n64) );
  OAI21X1 U136 ( .A(n1045), .B(n1009), .C(n65), .Y(n626) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n65) );
  OAI21X1 U138 ( .A(n1046), .B(n1009), .C(n66), .Y(n627) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n66) );
  OAI21X1 U140 ( .A(n1047), .B(n1009), .C(n67), .Y(n628) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n67) );
  OAI21X1 U142 ( .A(n1048), .B(n1009), .C(n68), .Y(n629) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n68) );
  OAI21X1 U144 ( .A(n1049), .B(n1009), .C(n69), .Y(n630) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n69) );
  NAND3X1 U146 ( .A(n70), .B(n48), .C(n71), .Y(n61) );
  OAI21X1 U147 ( .A(n1034), .B(n1008), .C(n73), .Y(n631) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n73) );
  OAI21X1 U149 ( .A(n1035), .B(n1008), .C(n74), .Y(n632) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n74) );
  OAI21X1 U151 ( .A(n1036), .B(n1008), .C(n75), .Y(n633) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n75) );
  OAI21X1 U153 ( .A(n1037), .B(n1008), .C(n76), .Y(n634) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n76) );
  OAI21X1 U155 ( .A(n1038), .B(n1008), .C(n77), .Y(n635) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n77) );
  OAI21X1 U157 ( .A(n1039), .B(n1008), .C(n78), .Y(n636) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n78) );
  OAI21X1 U159 ( .A(n1040), .B(n1008), .C(n79), .Y(n637) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n79) );
  OAI21X1 U161 ( .A(n1041), .B(n1008), .C(n80), .Y(n638) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n80) );
  NAND3X1 U163 ( .A(n973), .B(n1013), .C(n81), .Y(n72) );
  OAI21X1 U164 ( .A(n1042), .B(n1007), .C(n83), .Y(n639) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n83) );
  OAI21X1 U166 ( .A(n1043), .B(n1006), .C(n84), .Y(n640) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n84) );
  OAI21X1 U168 ( .A(n1044), .B(n1006), .C(n85), .Y(n641) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n85) );
  OAI21X1 U170 ( .A(n1045), .B(n1006), .C(n86), .Y(n642) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n86) );
  OAI21X1 U172 ( .A(n1046), .B(n1006), .C(n87), .Y(n643) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n87) );
  OAI21X1 U174 ( .A(n1047), .B(n1006), .C(n88), .Y(n644) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n88) );
  OAI21X1 U176 ( .A(n1048), .B(n1006), .C(n89), .Y(n645) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n89) );
  OAI21X1 U178 ( .A(n1049), .B(n1006), .C(n90), .Y(n646) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n90) );
  NAND3X1 U180 ( .A(n70), .B(n48), .C(n91), .Y(n82) );
  OAI21X1 U181 ( .A(n1034), .B(n1005), .C(n93), .Y(n647) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n93) );
  OAI21X1 U183 ( .A(n1035), .B(n1005), .C(n94), .Y(n648) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n94) );
  OAI21X1 U185 ( .A(n1036), .B(n1005), .C(n95), .Y(n649) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n95) );
  OAI21X1 U187 ( .A(n1037), .B(n1005), .C(n96), .Y(n650) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n96) );
  OAI21X1 U189 ( .A(n1038), .B(n1005), .C(n97), .Y(n651) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n97) );
  OAI21X1 U191 ( .A(n1039), .B(n1005), .C(n98), .Y(n652) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n98) );
  OAI21X1 U193 ( .A(n1040), .B(n1005), .C(n99), .Y(n653) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n99) );
  OAI21X1 U195 ( .A(n1041), .B(n1005), .C(n100), .Y(n654) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n100) );
  NAND3X1 U197 ( .A(n973), .B(n1012), .C(n101), .Y(n92) );
  OAI21X1 U198 ( .A(n1042), .B(n1004), .C(n103), .Y(n655) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n103) );
  OAI21X1 U200 ( .A(n1043), .B(n1003), .C(n104), .Y(n656) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n104) );
  OAI21X1 U202 ( .A(n1044), .B(n1003), .C(n105), .Y(n657) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n105) );
  OAI21X1 U204 ( .A(n1045), .B(n1003), .C(n106), .Y(n658) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n106) );
  OAI21X1 U206 ( .A(n1046), .B(n1003), .C(n107), .Y(n659) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n107) );
  OAI21X1 U208 ( .A(n1047), .B(n1003), .C(n108), .Y(n660) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n108) );
  OAI21X1 U210 ( .A(n1048), .B(n1003), .C(n109), .Y(n661) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n109) );
  OAI21X1 U212 ( .A(n1049), .B(n1003), .C(n110), .Y(n662) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n110) );
  NAND3X1 U214 ( .A(n71), .B(n1013), .C(n111), .Y(n102) );
  OAI21X1 U215 ( .A(n1034), .B(n1002), .C(n113), .Y(n663) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n113) );
  OAI21X1 U217 ( .A(n1035), .B(n1002), .C(n114), .Y(n664) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n114) );
  OAI21X1 U219 ( .A(n1036), .B(n1002), .C(n115), .Y(n665) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n115) );
  OAI21X1 U221 ( .A(n1037), .B(n1002), .C(n116), .Y(n666) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n116) );
  OAI21X1 U223 ( .A(n1038), .B(n1002), .C(n117), .Y(n667) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n117) );
  OAI21X1 U225 ( .A(n1039), .B(n1002), .C(n118), .Y(n668) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n118) );
  OAI21X1 U227 ( .A(n1040), .B(n1002), .C(n119), .Y(n669) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n119) );
  OAI21X1 U229 ( .A(n1041), .B(n1002), .C(n120), .Y(n670) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n120) );
  NAND3X1 U231 ( .A(n973), .B(n1013), .C(n121), .Y(n112) );
  OAI21X1 U232 ( .A(n1042), .B(n1001), .C(n123), .Y(n671) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n123) );
  OAI21X1 U234 ( .A(n1043), .B(n1000), .C(n124), .Y(n672) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n124) );
  OAI21X1 U236 ( .A(n1044), .B(n1000), .C(n125), .Y(n673) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n125) );
  OAI21X1 U238 ( .A(n1045), .B(n1000), .C(n126), .Y(n674) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n126) );
  OAI21X1 U240 ( .A(n1046), .B(n1000), .C(n127), .Y(n675) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n127) );
  OAI21X1 U242 ( .A(n1047), .B(n1000), .C(n128), .Y(n676) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n128) );
  OAI21X1 U244 ( .A(n1048), .B(n1000), .C(n129), .Y(n677) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n129) );
  OAI21X1 U246 ( .A(n1049), .B(n1000), .C(n130), .Y(n678) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n130) );
  NAND3X1 U248 ( .A(n91), .B(n1013), .C(n111), .Y(n122) );
  OAI21X1 U249 ( .A(n1034), .B(n999), .C(n132), .Y(n679) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n132) );
  OAI21X1 U251 ( .A(n1035), .B(n999), .C(n133), .Y(n680) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n133) );
  OAI21X1 U253 ( .A(n1036), .B(n999), .C(n134), .Y(n681) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n134) );
  OAI21X1 U255 ( .A(n1037), .B(n999), .C(n135), .Y(n682) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n135) );
  OAI21X1 U257 ( .A(n1038), .B(n999), .C(n136), .Y(n683) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n136) );
  OAI21X1 U259 ( .A(n1039), .B(n999), .C(n137), .Y(n684) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n137) );
  OAI21X1 U261 ( .A(n1040), .B(n999), .C(n138), .Y(n685) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n138) );
  OAI21X1 U263 ( .A(n1041), .B(n999), .C(n139), .Y(n686) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n139) );
  NAND3X1 U265 ( .A(n973), .B(n1013), .C(n140), .Y(n131) );
  OAI21X1 U266 ( .A(n1042), .B(n998), .C(n142), .Y(n687) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n142) );
  OAI21X1 U268 ( .A(n1043), .B(n998), .C(n143), .Y(n688) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n143) );
  OAI21X1 U270 ( .A(n1044), .B(n998), .C(n144), .Y(n689) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n144) );
  OAI21X1 U272 ( .A(n1045), .B(n998), .C(n145), .Y(n690) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n145) );
  OAI21X1 U274 ( .A(n1046), .B(n998), .C(n146), .Y(n691) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n146) );
  OAI21X1 U276 ( .A(n1047), .B(n998), .C(n147), .Y(n692) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n147) );
  OAI21X1 U278 ( .A(n1048), .B(n998), .C(n148), .Y(n693) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n148) );
  OAI21X1 U280 ( .A(n1049), .B(n998), .C(n149), .Y(n694) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n149) );
  NAND3X1 U282 ( .A(n71), .B(n1013), .C(n969), .Y(n141) );
  OAI21X1 U283 ( .A(n1034), .B(n997), .C(n152), .Y(n695) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n152) );
  OAI21X1 U285 ( .A(n1035), .B(n997), .C(n153), .Y(n696) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n153) );
  OAI21X1 U287 ( .A(n1036), .B(n997), .C(n154), .Y(n697) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n154) );
  OAI21X1 U289 ( .A(n1037), .B(n997), .C(n155), .Y(n698) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n155) );
  OAI21X1 U291 ( .A(n1038), .B(n997), .C(n156), .Y(n699) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n156) );
  OAI21X1 U293 ( .A(n1039), .B(n997), .C(n157), .Y(n700) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n157) );
  OAI21X1 U295 ( .A(n1040), .B(n997), .C(n158), .Y(n701) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n158) );
  OAI21X1 U297 ( .A(n1041), .B(n997), .C(n159), .Y(n702) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n159) );
  NAND3X1 U299 ( .A(n973), .B(n1013), .C(n160), .Y(n151) );
  OAI21X1 U300 ( .A(n1042), .B(n996), .C(n162), .Y(n703) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n162) );
  OAI21X1 U302 ( .A(n1043), .B(n996), .C(n163), .Y(n704) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n163) );
  OAI21X1 U304 ( .A(n1044), .B(n996), .C(n164), .Y(n705) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n164) );
  OAI21X1 U306 ( .A(n1045), .B(n996), .C(n165), .Y(n706) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n165) );
  OAI21X1 U308 ( .A(n1046), .B(n996), .C(n166), .Y(n707) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n166) );
  OAI21X1 U310 ( .A(n1047), .B(n996), .C(n167), .Y(n708) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n167) );
  OAI21X1 U312 ( .A(n1048), .B(n996), .C(n168), .Y(n709) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n168) );
  OAI21X1 U314 ( .A(n1049), .B(n996), .C(n169), .Y(n710) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n169) );
  NAND3X1 U316 ( .A(n91), .B(n1013), .C(n969), .Y(n161) );
  OAI21X1 U317 ( .A(n1034), .B(n995), .C(n171), .Y(n711) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n171) );
  OAI21X1 U319 ( .A(n1035), .B(n995), .C(n172), .Y(n712) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n172) );
  OAI21X1 U321 ( .A(n1036), .B(n995), .C(n173), .Y(n713) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n173) );
  OAI21X1 U323 ( .A(n1037), .B(n995), .C(n174), .Y(n714) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n174) );
  OAI21X1 U325 ( .A(n1038), .B(n995), .C(n175), .Y(n715) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n175) );
  OAI21X1 U327 ( .A(n1039), .B(n995), .C(n176), .Y(n716) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n176) );
  OAI21X1 U329 ( .A(n1040), .B(n995), .C(n177), .Y(n717) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n177) );
  OAI21X1 U331 ( .A(n1041), .B(n995), .C(n178), .Y(n718) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n178) );
  NAND3X1 U333 ( .A(n973), .B(n1013), .C(n179), .Y(n170) );
  OAI21X1 U334 ( .A(n1042), .B(n994), .C(n181), .Y(n719) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n181) );
  OAI21X1 U336 ( .A(n1043), .B(n994), .C(n182), .Y(n720) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n182) );
  OAI21X1 U338 ( .A(n1044), .B(n994), .C(n183), .Y(n721) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n183) );
  OAI21X1 U340 ( .A(n1045), .B(n994), .C(n184), .Y(n722) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n184) );
  OAI21X1 U342 ( .A(n1046), .B(n994), .C(n185), .Y(n723) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n185) );
  OAI21X1 U344 ( .A(n1047), .B(n994), .C(n186), .Y(n724) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n186) );
  OAI21X1 U346 ( .A(n1048), .B(n994), .C(n187), .Y(n725) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n187) );
  OAI21X1 U348 ( .A(n1049), .B(n994), .C(n188), .Y(n726) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n188) );
  NAND3X1 U350 ( .A(n71), .B(n1013), .C(n967), .Y(n180) );
  OAI21X1 U351 ( .A(n1034), .B(n993), .C(n191), .Y(n727) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n191) );
  OAI21X1 U353 ( .A(n1035), .B(n993), .C(n192), .Y(n728) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n192) );
  OAI21X1 U355 ( .A(n1036), .B(n993), .C(n193), .Y(n729) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n193) );
  OAI21X1 U357 ( .A(n1037), .B(n993), .C(n194), .Y(n730) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n194) );
  OAI21X1 U359 ( .A(n1038), .B(n993), .C(n195), .Y(n731) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n195) );
  OAI21X1 U361 ( .A(n1039), .B(n993), .C(n196), .Y(n732) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n196) );
  OAI21X1 U363 ( .A(n1040), .B(n993), .C(n197), .Y(n733) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n197) );
  OAI21X1 U365 ( .A(n1041), .B(n993), .C(n198), .Y(n734) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n198) );
  NAND3X1 U367 ( .A(n973), .B(n1013), .C(n199), .Y(n190) );
  OAI21X1 U368 ( .A(n1042), .B(n992), .C(n201), .Y(n735) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n201) );
  OAI21X1 U370 ( .A(n1043), .B(n992), .C(n202), .Y(n736) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n202) );
  OAI21X1 U372 ( .A(n1044), .B(n992), .C(n203), .Y(n737) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n203) );
  OAI21X1 U374 ( .A(n1045), .B(n992), .C(n204), .Y(n738) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n204) );
  OAI21X1 U376 ( .A(n1046), .B(n992), .C(n205), .Y(n739) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n205) );
  OAI21X1 U378 ( .A(n1047), .B(n992), .C(n206), .Y(n740) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n206) );
  OAI21X1 U380 ( .A(n1048), .B(n992), .C(n207), .Y(n741) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n207) );
  OAI21X1 U382 ( .A(n1049), .B(n992), .C(n208), .Y(n742) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n208) );
  NAND3X1 U384 ( .A(n91), .B(n1013), .C(n967), .Y(n200) );
  OAI21X1 U385 ( .A(n1034), .B(n991), .C(n210), .Y(n743) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n210) );
  OAI21X1 U387 ( .A(n1035), .B(n991), .C(n211), .Y(n744) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n211) );
  OAI21X1 U389 ( .A(n1036), .B(n991), .C(n212), .Y(n745) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n212) );
  OAI21X1 U391 ( .A(n1037), .B(n991), .C(n213), .Y(n746) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n213) );
  OAI21X1 U393 ( .A(n1038), .B(n991), .C(n214), .Y(n747) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n214) );
  OAI21X1 U395 ( .A(n1039), .B(n991), .C(n215), .Y(n748) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n215) );
  OAI21X1 U397 ( .A(n1040), .B(n991), .C(n216), .Y(n749) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n216) );
  OAI21X1 U399 ( .A(n1041), .B(n991), .C(n217), .Y(n750) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n217) );
  NAND3X1 U401 ( .A(n973), .B(n1013), .C(n218), .Y(n209) );
  OAI21X1 U402 ( .A(n1042), .B(n990), .C(n220), .Y(n751) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n220) );
  OAI21X1 U404 ( .A(n1043), .B(n989), .C(n221), .Y(n752) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n221) );
  OAI21X1 U406 ( .A(n1044), .B(n989), .C(n222), .Y(n753) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n222) );
  OAI21X1 U408 ( .A(n1045), .B(n989), .C(n223), .Y(n754) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n223) );
  OAI21X1 U410 ( .A(n1046), .B(n989), .C(n224), .Y(n755) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n224) );
  OAI21X1 U412 ( .A(n1047), .B(n989), .C(n225), .Y(n756) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n225) );
  OAI21X1 U414 ( .A(n1048), .B(n989), .C(n226), .Y(n757) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n226) );
  OAI21X1 U416 ( .A(n1049), .B(n989), .C(n227), .Y(n758) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n227) );
  NAND3X1 U418 ( .A(n70), .B(n1012), .C(n228), .Y(n219) );
  OAI21X1 U419 ( .A(n1034), .B(n988), .C(n230), .Y(n759) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n230) );
  OAI21X1 U421 ( .A(n1035), .B(n988), .C(n231), .Y(n760) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n231) );
  OAI21X1 U423 ( .A(n1036), .B(n988), .C(n232), .Y(n761) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n232) );
  OAI21X1 U425 ( .A(n1037), .B(n988), .C(n233), .Y(n762) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n233) );
  OAI21X1 U427 ( .A(n1038), .B(n988), .C(n234), .Y(n763) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n234) );
  OAI21X1 U429 ( .A(n1039), .B(n988), .C(n235), .Y(n764) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n235) );
  OAI21X1 U431 ( .A(n1040), .B(n988), .C(n236), .Y(n765) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n236) );
  OAI21X1 U433 ( .A(n1041), .B(n988), .C(n237), .Y(n766) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n237) );
  NAND3X1 U435 ( .A(n973), .B(n1012), .C(n238), .Y(n229) );
  OAI21X1 U436 ( .A(n1042), .B(n987), .C(n240), .Y(n767) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n240) );
  OAI21X1 U438 ( .A(n1043), .B(n986), .C(n241), .Y(n768) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n241) );
  OAI21X1 U440 ( .A(n1044), .B(n986), .C(n242), .Y(n769) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n242) );
  OAI21X1 U442 ( .A(n1045), .B(n986), .C(n243), .Y(n770) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n243) );
  OAI21X1 U444 ( .A(n1046), .B(n986), .C(n244), .Y(n771) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n244) );
  OAI21X1 U446 ( .A(n1047), .B(n986), .C(n245), .Y(n772) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n245) );
  OAI21X1 U448 ( .A(n1048), .B(n986), .C(n246), .Y(n773) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n246) );
  OAI21X1 U450 ( .A(n1049), .B(n986), .C(n247), .Y(n774) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n247) );
  NAND3X1 U452 ( .A(n70), .B(n1012), .C(n248), .Y(n239) );
  OAI21X1 U453 ( .A(n1034), .B(n985), .C(n251), .Y(n775) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n251) );
  OAI21X1 U455 ( .A(n1035), .B(n985), .C(n252), .Y(n776) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n252) );
  OAI21X1 U457 ( .A(n1036), .B(n985), .C(n253), .Y(n777) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n253) );
  OAI21X1 U459 ( .A(n1037), .B(n985), .C(n254), .Y(n778) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n254) );
  OAI21X1 U461 ( .A(n1038), .B(n985), .C(n255), .Y(n779) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n255) );
  OAI21X1 U463 ( .A(n1039), .B(n985), .C(n256), .Y(n780) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n256) );
  OAI21X1 U465 ( .A(n1040), .B(n985), .C(n257), .Y(n781) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n257) );
  OAI21X1 U467 ( .A(n1041), .B(n985), .C(n258), .Y(n782) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n258) );
  NAND3X1 U469 ( .A(n973), .B(n1012), .C(n259), .Y(n250) );
  OAI21X1 U470 ( .A(n1042), .B(n984), .C(n261), .Y(n783) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n261) );
  OAI21X1 U472 ( .A(n1043), .B(n983), .C(n262), .Y(n784) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n262) );
  OAI21X1 U474 ( .A(n1044), .B(n983), .C(n263), .Y(n785) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n263) );
  OAI21X1 U476 ( .A(n1045), .B(n983), .C(n264), .Y(n786) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n264) );
  OAI21X1 U478 ( .A(n1046), .B(n983), .C(n265), .Y(n787) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n265) );
  OAI21X1 U480 ( .A(n1047), .B(n983), .C(n266), .Y(n788) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n266) );
  OAI21X1 U482 ( .A(n1048), .B(n983), .C(n267), .Y(n789) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n267) );
  OAI21X1 U484 ( .A(n1049), .B(n983), .C(n268), .Y(n790) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n268) );
  NAND3X1 U486 ( .A(n111), .B(n1012), .C(n228), .Y(n260) );
  OAI21X1 U487 ( .A(n1034), .B(n982), .C(n270), .Y(n791) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n270) );
  OAI21X1 U489 ( .A(n1035), .B(n982), .C(n271), .Y(n792) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n271) );
  OAI21X1 U491 ( .A(n1036), .B(n982), .C(n272), .Y(n793) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n272) );
  OAI21X1 U493 ( .A(n1037), .B(n982), .C(n273), .Y(n794) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n273) );
  OAI21X1 U495 ( .A(n1038), .B(n982), .C(n274), .Y(n795) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n274) );
  OAI21X1 U497 ( .A(n1039), .B(n982), .C(n275), .Y(n796) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n275) );
  OAI21X1 U499 ( .A(n1040), .B(n982), .C(n276), .Y(n797) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n276) );
  OAI21X1 U501 ( .A(n1041), .B(n982), .C(n277), .Y(n798) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n277) );
  NAND3X1 U503 ( .A(n973), .B(n1012), .C(n278), .Y(n269) );
  OAI21X1 U504 ( .A(n1042), .B(n981), .C(n280), .Y(n799) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n280) );
  OAI21X1 U506 ( .A(n1043), .B(n980), .C(n281), .Y(n800) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n281) );
  OAI21X1 U508 ( .A(n1044), .B(n980), .C(n282), .Y(n801) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n282) );
  OAI21X1 U510 ( .A(n1045), .B(n980), .C(n283), .Y(n802) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n283) );
  OAI21X1 U512 ( .A(n1046), .B(n980), .C(n284), .Y(n803) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n284) );
  OAI21X1 U514 ( .A(n1047), .B(n980), .C(n285), .Y(n804) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n285) );
  OAI21X1 U516 ( .A(n1048), .B(n980), .C(n286), .Y(n805) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n286) );
  OAI21X1 U518 ( .A(n1049), .B(n980), .C(n287), .Y(n806) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n287) );
  NAND3X1 U520 ( .A(n111), .B(n1012), .C(n248), .Y(n279) );
  OAI21X1 U521 ( .A(n1034), .B(n979), .C(n291), .Y(n807) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n291) );
  OAI21X1 U523 ( .A(n1035), .B(n979), .C(n292), .Y(n808) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n292) );
  OAI21X1 U525 ( .A(n1036), .B(n979), .C(n293), .Y(n809) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n293) );
  OAI21X1 U527 ( .A(n1037), .B(n979), .C(n294), .Y(n810) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n294) );
  OAI21X1 U529 ( .A(n1038), .B(n979), .C(n295), .Y(n811) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n295) );
  OAI21X1 U531 ( .A(n1039), .B(n979), .C(n296), .Y(n812) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n296) );
  OAI21X1 U533 ( .A(n1040), .B(n979), .C(n297), .Y(n813) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n297) );
  OAI21X1 U535 ( .A(n1041), .B(n979), .C(n298), .Y(n814) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n298) );
  NAND3X1 U537 ( .A(n973), .B(n1012), .C(n299), .Y(n290) );
  OAI21X1 U538 ( .A(n1042), .B(n978), .C(n301), .Y(n815) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n301) );
  OAI21X1 U540 ( .A(n1043), .B(n978), .C(n302), .Y(n816) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n302) );
  OAI21X1 U542 ( .A(n1044), .B(n978), .C(n303), .Y(n817) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n303) );
  OAI21X1 U544 ( .A(n1045), .B(n978), .C(n304), .Y(n818) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n304) );
  OAI21X1 U546 ( .A(n1046), .B(n978), .C(n305), .Y(n819) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n305) );
  OAI21X1 U548 ( .A(n1047), .B(n978), .C(n306), .Y(n820) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n306) );
  OAI21X1 U550 ( .A(n1048), .B(n978), .C(n307), .Y(n821) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n307) );
  OAI21X1 U552 ( .A(n1049), .B(n978), .C(n308), .Y(n822) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n308) );
  NAND3X1 U554 ( .A(n969), .B(n1012), .C(n228), .Y(n300) );
  OAI21X1 U555 ( .A(n1034), .B(n977), .C(n310), .Y(n823) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n310) );
  OAI21X1 U557 ( .A(n1035), .B(n977), .C(n311), .Y(n824) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n311) );
  OAI21X1 U559 ( .A(n1036), .B(n977), .C(n312), .Y(n825) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n312) );
  OAI21X1 U561 ( .A(n1037), .B(n977), .C(n313), .Y(n826) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n313) );
  OAI21X1 U563 ( .A(n1038), .B(n977), .C(n314), .Y(n827) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n314) );
  OAI21X1 U565 ( .A(n1039), .B(n977), .C(n315), .Y(n828) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n315) );
  OAI21X1 U567 ( .A(n1040), .B(n977), .C(n316), .Y(n829) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n316) );
  OAI21X1 U569 ( .A(n1041), .B(n977), .C(n317), .Y(n830) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n317) );
  NAND3X1 U571 ( .A(n973), .B(n1012), .C(n318), .Y(n309) );
  OAI21X1 U572 ( .A(n1042), .B(n976), .C(n320), .Y(n831) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n320) );
  OAI21X1 U574 ( .A(n1043), .B(n976), .C(n321), .Y(n832) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n321) );
  OAI21X1 U576 ( .A(n1044), .B(n976), .C(n322), .Y(n833) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n322) );
  OAI21X1 U578 ( .A(n1045), .B(n976), .C(n323), .Y(n834) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n323) );
  OAI21X1 U580 ( .A(n1046), .B(n976), .C(n324), .Y(n835) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n324) );
  OAI21X1 U582 ( .A(n1047), .B(n976), .C(n325), .Y(n836) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n325) );
  OAI21X1 U584 ( .A(n1048), .B(n976), .C(n326), .Y(n837) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n326) );
  OAI21X1 U586 ( .A(n1049), .B(n976), .C(n327), .Y(n838) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n327) );
  NAND3X1 U588 ( .A(n969), .B(n1012), .C(n248), .Y(n319) );
  OAI21X1 U590 ( .A(n1034), .B(n975), .C(n330), .Y(n839) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n330) );
  OAI21X1 U592 ( .A(n1035), .B(n975), .C(n331), .Y(n840) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n331) );
  OAI21X1 U594 ( .A(n1036), .B(n975), .C(n332), .Y(n841) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n332) );
  OAI21X1 U596 ( .A(n1037), .B(n975), .C(n333), .Y(n842) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n333) );
  OAI21X1 U598 ( .A(n1038), .B(n975), .C(n334), .Y(n843) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n334) );
  OAI21X1 U600 ( .A(n1039), .B(n975), .C(n335), .Y(n844) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n335) );
  OAI21X1 U602 ( .A(n1040), .B(n975), .C(n336), .Y(n845) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n336) );
  OAI21X1 U604 ( .A(n1041), .B(n975), .C(n337), .Y(n846) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n337) );
  NAND3X1 U606 ( .A(n973), .B(n1012), .C(n338), .Y(n329) );
  OAI21X1 U607 ( .A(n1042), .B(n974), .C(n340), .Y(n847) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n340) );
  OAI21X1 U609 ( .A(n1043), .B(n974), .C(n341), .Y(n848) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n341) );
  OAI21X1 U611 ( .A(n1044), .B(n974), .C(n342), .Y(n849) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n342) );
  OAI21X1 U613 ( .A(n1045), .B(n974), .C(n343), .Y(n850) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n343) );
  OAI21X1 U615 ( .A(n1046), .B(n974), .C(n344), .Y(n851) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n344) );
  OAI21X1 U617 ( .A(n1047), .B(n974), .C(n345), .Y(n852) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n345) );
  OAI21X1 U619 ( .A(n1048), .B(n974), .C(n346), .Y(n853) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n346) );
  OAI21X1 U621 ( .A(n1049), .B(n974), .C(n347), .Y(n854) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n347) );
  NAND3X1 U623 ( .A(n967), .B(n1012), .C(n228), .Y(n339) );
  OAI21X1 U624 ( .A(n1034), .B(n8), .C(n349), .Y(n855) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n349) );
  OAI21X1 U626 ( .A(n1035), .B(n8), .C(n350), .Y(n856) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n350) );
  OAI21X1 U628 ( .A(n1036), .B(n8), .C(n351), .Y(n857) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n351) );
  OAI21X1 U630 ( .A(n1037), .B(n8), .C(n352), .Y(n858) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n352) );
  OAI21X1 U632 ( .A(n1038), .B(n8), .C(n353), .Y(n859) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n353) );
  OAI21X1 U634 ( .A(n1039), .B(n8), .C(n354), .Y(n860) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n354) );
  OAI21X1 U636 ( .A(n1040), .B(n8), .C(n355), .Y(n861) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n355) );
  OAI21X1 U638 ( .A(n1041), .B(n8), .C(n356), .Y(n862) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n356) );
  NOR2X1 U641 ( .A(n964), .B(\addr_1c<4> ), .Y(n59) );
  OAI21X1 U642 ( .A(n1042), .B(n972), .C(n359), .Y(n863) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n359) );
  OAI21X1 U644 ( .A(n1043), .B(n972), .C(n360), .Y(n864) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n360) );
  OAI21X1 U646 ( .A(n1044), .B(n972), .C(n361), .Y(n865) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n361) );
  OAI21X1 U648 ( .A(n1045), .B(n972), .C(n362), .Y(n866) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n362) );
  OAI21X1 U650 ( .A(n1046), .B(n972), .C(n363), .Y(n867) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n363) );
  OAI21X1 U652 ( .A(n1047), .B(n972), .C(n364), .Y(n868) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n364) );
  OAI21X1 U654 ( .A(n1048), .B(n972), .C(n365), .Y(n869) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n365) );
  OAI21X1 U656 ( .A(n1049), .B(n972), .C(n366), .Y(n870) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n366) );
  NAND3X1 U658 ( .A(n967), .B(n1013), .C(n248), .Y(n358) );
  NOR3X1 U661 ( .A(n370), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n369) );
  NOR3X1 U662 ( .A(n371), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n368) );
  AOI21X1 U663 ( .A(n473), .B(n373), .C(n963), .Y(n1050) );
  OAI21X1 U665 ( .A(rd), .B(n374), .C(wr), .Y(n373) );
  NAND3X1 U667 ( .A(n375), .B(n1029), .C(n376), .Y(n374) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n376) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n375) );
  AOI21X1 U670 ( .A(n460), .B(n378), .C(n1020), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n380), .C(n4), .Y(n378) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n91), .C(\mem<0><1> ), .D(n248), .Y(n383) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n71), .C(\mem<2><1> ), .D(n228), .Y(n382) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n91), .C(\mem<4><1> ), .D(n248), .Y(n385) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n71), .C(\mem<6><1> ), .D(n228), .Y(n384) );
  AOI22X1 U678 ( .A(n288), .B(n893), .C(n249), .D(n933), .Y(n377) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n91), .C(\mem<12><1> ), .D(n248), .Y(
        n389) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n71), .C(\mem<14><1> ), .D(n228), .Y(
        n388) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n91), .C(\mem<8><1> ), .D(n248), .Y(n391) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n71), .C(\mem<10><1> ), .D(n228), .Y(
        n390) );
  AOI21X1 U685 ( .A(n448), .B(n393), .C(n1020), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n940), .B(n395), .C(n950), .Y(n393) );
  AOI21X1 U687 ( .A(n397), .B(n398), .C(n971), .Y(n396) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n91), .C(\mem<0><0> ), .D(n248), .Y(n398) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n71), .C(\mem<2><0> ), .D(n228), .Y(n397) );
  AOI21X1 U690 ( .A(n399), .B(n400), .C(n970), .Y(n394) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n91), .C(\mem<4><0> ), .D(n248), .Y(n400) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n71), .C(\mem<6><0> ), .D(n228), .Y(n399) );
  AOI22X1 U693 ( .A(n288), .B(n891), .C(n249), .D(n931), .Y(n392) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n91), .C(\mem<12><0> ), .D(n248), .Y(
        n404) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n71), .C(\mem<14><0> ), .D(n228), .Y(
        n403) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n91), .C(\mem<8><0> ), .D(n248), .Y(n406) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n71), .C(\mem<10><0> ), .D(n228), .Y(
        n405) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n407) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n199), .C(\mem<19><7> ), .D(n179), .Y(
        n414) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n160), .C(\mem<23><7> ), .D(n140), .Y(
        n413) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n121), .C(\mem<27><7> ), .D(n101), .Y(
        n411) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n81), .C(\mem<31><7> ), .D(n60), .Y(n410) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n357), .C(\mem<3><7> ), .D(n338), .Y(n419) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n318), .C(\mem<7><7> ), .D(n299), .Y(n418) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n278), .C(\mem<11><7> ), .D(n259), .Y(
        n416) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n238), .C(\mem<15><7> ), .D(n218), .Y(
        n415) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n420) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n199), .C(\mem<19><6> ), .D(n179), .Y(
        n427) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n160), .C(\mem<23><6> ), .D(n140), .Y(
        n426) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n121), .C(\mem<27><6> ), .D(n101), .Y(
        n424) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n81), .C(\mem<31><6> ), .D(n60), .Y(n423) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n357), .C(\mem<3><6> ), .D(n338), .Y(n432) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n318), .C(\mem<7><6> ), .D(n299), .Y(n431) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n278), .C(\mem<11><6> ), .D(n259), .Y(
        n429) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n238), .C(\mem<15><6> ), .D(n218), .Y(
        n428) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n433) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n199), .C(\mem<19><5> ), .D(n179), .Y(
        n440) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n160), .C(\mem<23><5> ), .D(n140), .Y(
        n439) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n121), .C(\mem<27><5> ), .D(n101), .Y(
        n437) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n81), .C(\mem<31><5> ), .D(n60), .Y(n436) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n357), .C(\mem<3><5> ), .D(n338), .Y(n445) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n318), .C(\mem<7><5> ), .D(n299), .Y(n444) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n278), .C(\mem<11><5> ), .D(n259), .Y(
        n442) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n238), .C(\mem<15><5> ), .D(n218), .Y(
        n441) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n446) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n199), .C(\mem<19><4> ), .D(n179), .Y(
        n453) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n160), .C(\mem<23><4> ), .D(n140), .Y(
        n452) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n121), .C(\mem<27><4> ), .D(n101), .Y(
        n450) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n81), .C(\mem<31><4> ), .D(n60), .Y(n449) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n357), .C(\mem<3><4> ), .D(n338), .Y(n458) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n318), .C(\mem<7><4> ), .D(n299), .Y(n457) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n278), .C(\mem<11><4> ), .D(n259), .Y(
        n455) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n238), .C(\mem<15><4> ), .D(n218), .Y(
        n454) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n459) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n199), .C(\mem<19><3> ), .D(n179), .Y(
        n466) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n160), .C(\mem<23><3> ), .D(n140), .Y(
        n465) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n121), .C(\mem<27><3> ), .D(n101), .Y(
        n463) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n81), .C(\mem<31><3> ), .D(n60), .Y(n462) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n357), .C(\mem<3><3> ), .D(n338), .Y(n471) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n318), .C(\mem<7><3> ), .D(n299), .Y(n470) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n278), .C(\mem<11><3> ), .D(n259), .Y(
        n468) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n238), .C(\mem<15><3> ), .D(n218), .Y(
        n467) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n472) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n199), .C(\mem<19><2> ), .D(n179), .Y(
        n479) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n160), .C(\mem<23><2> ), .D(n140), .Y(
        n478) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n121), .C(\mem<27><2> ), .D(n101), .Y(
        n476) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n81), .C(\mem<31><2> ), .D(n60), .Y(n475) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n357), .C(\mem<3><2> ), .D(n338), .Y(n484) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n318), .C(\mem<7><2> ), .D(n299), .Y(n483) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n278), .C(\mem<11><2> ), .D(n259), .Y(
        n481) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n238), .C(\mem<15><2> ), .D(n218), .Y(
        n480) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n485) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n199), .C(\mem<19><1> ), .D(n179), .Y(
        n492) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n160), .C(\mem<23><1> ), .D(n140), .Y(
        n491) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n121), .C(\mem<27><1> ), .D(n101), .Y(
        n489) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n81), .C(\mem<31><1> ), .D(n60), .Y(n488) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n357), .C(\mem<3><1> ), .D(n338), .Y(n497) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n318), .C(\mem<7><1> ), .D(n299), .Y(n496) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n278), .C(\mem<11><1> ), .D(n259), .Y(
        n494) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n238), .C(\mem<15><1> ), .D(n218), .Y(
        n493) );
  AOI21X1 U777 ( .A(n447), .B(n499), .C(n1020), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n939), .B(n501), .C(n949), .Y(n499) );
  AOI21X1 U779 ( .A(n503), .B(n504), .C(n971), .Y(n502) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n91), .C(\mem<0><7> ), .D(n248), .Y(n504) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n71), .C(\mem<2><7> ), .D(n228), .Y(n503) );
  AOI21X1 U782 ( .A(n505), .B(n506), .C(n970), .Y(n500) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n91), .C(\mem<4><7> ), .D(n248), .Y(n506) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n71), .C(\mem<6><7> ), .D(n228), .Y(n505) );
  AOI22X1 U785 ( .A(n288), .B(n889), .C(n249), .D(n929), .Y(n498) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n91), .C(\mem<12><7> ), .D(n248), .Y(
        n510) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n71), .C(\mem<14><7> ), .D(n228), .Y(
        n509) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n91), .C(\mem<8><7> ), .D(n248), .Y(n512) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n71), .C(\mem<10><7> ), .D(n228), .Y(
        n511) );
  AOI21X1 U792 ( .A(n435), .B(n514), .C(n1020), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n938), .B(n516), .C(n948), .Y(n514) );
  AOI21X1 U794 ( .A(n518), .B(n519), .C(n971), .Y(n517) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n91), .C(\mem<0><6> ), .D(n248), .Y(n519) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n71), .C(\mem<2><6> ), .D(n228), .Y(n518) );
  AOI21X1 U797 ( .A(n520), .B(n521), .C(n970), .Y(n515) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n91), .C(\mem<4><6> ), .D(n248), .Y(n521) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n71), .C(\mem<6><6> ), .D(n228), .Y(n520) );
  AOI22X1 U800 ( .A(n288), .B(n887), .C(n249), .D(n927), .Y(n513) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n91), .C(\mem<12><6> ), .D(n248), .Y(
        n525) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n71), .C(\mem<14><6> ), .D(n228), .Y(
        n524) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n91), .C(\mem<8><6> ), .D(n248), .Y(n527) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n71), .C(\mem<10><6> ), .D(n228), .Y(
        n526) );
  AOI21X1 U807 ( .A(n434), .B(n529), .C(n1020), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n937), .B(n531), .C(n947), .Y(n529) );
  AOI21X1 U809 ( .A(n533), .B(n534), .C(n971), .Y(n532) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n91), .C(\mem<0><5> ), .D(n248), .Y(n534) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n71), .C(\mem<2><5> ), .D(n228), .Y(n533) );
  AOI21X1 U812 ( .A(n535), .B(n536), .C(n970), .Y(n530) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n91), .C(\mem<4><5> ), .D(n248), .Y(n536) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n71), .C(\mem<6><5> ), .D(n228), .Y(n535) );
  AOI22X1 U815 ( .A(n288), .B(n885), .C(n249), .D(n925), .Y(n528) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n91), .C(\mem<12><5> ), .D(n248), .Y(
        n540) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n71), .C(\mem<14><5> ), .D(n228), .Y(
        n539) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n91), .C(\mem<8><5> ), .D(n248), .Y(n542) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n71), .C(\mem<10><5> ), .D(n228), .Y(
        n541) );
  AOI21X1 U822 ( .A(n422), .B(n544), .C(n1020), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n936), .B(n546), .C(n946), .Y(n544) );
  AOI21X1 U824 ( .A(n548), .B(n549), .C(n971), .Y(n547) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n91), .C(\mem<0><4> ), .D(n248), .Y(n549) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n71), .C(\mem<2><4> ), .D(n228), .Y(n548) );
  AOI21X1 U827 ( .A(n550), .B(n551), .C(n970), .Y(n545) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n91), .C(\mem<4><4> ), .D(n248), .Y(n551) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n71), .C(\mem<6><4> ), .D(n228), .Y(n550) );
  AOI22X1 U830 ( .A(n288), .B(n883), .C(n249), .D(n923), .Y(n543) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n91), .C(\mem<12><4> ), .D(n248), .Y(
        n555) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n71), .C(\mem<14><4> ), .D(n228), .Y(
        n554) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n91), .C(\mem<8><4> ), .D(n248), .Y(n557) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n71), .C(\mem<10><4> ), .D(n228), .Y(
        n556) );
  AOI21X1 U837 ( .A(n421), .B(n559), .C(n1020), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n935), .B(n561), .C(n945), .Y(n559) );
  AOI21X1 U839 ( .A(n563), .B(n564), .C(n971), .Y(n562) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n91), .C(\mem<0><3> ), .D(n248), .Y(n564) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n71), .C(\mem<2><3> ), .D(n228), .Y(n563) );
  AOI21X1 U842 ( .A(n565), .B(n566), .C(n970), .Y(n560) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n91), .C(\mem<4><3> ), .D(n248), .Y(n566) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n71), .C(\mem<6><3> ), .D(n228), .Y(n565) );
  AOI22X1 U845 ( .A(n288), .B(n881), .C(n249), .D(n921), .Y(n558) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n91), .C(\mem<12><3> ), .D(n248), .Y(
        n570) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n71), .C(\mem<14><3> ), .D(n228), .Y(
        n569) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n91), .C(\mem<8><3> ), .D(n248), .Y(n572) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n71), .C(\mem<10><3> ), .D(n228), .Y(
        n571) );
  AOI21X1 U852 ( .A(n409), .B(n574), .C(n1020), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n934), .B(n576), .C(n944), .Y(n574) );
  AOI21X1 U854 ( .A(n578), .B(n579), .C(n971), .Y(n577) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n91), .C(\mem<0><2> ), .D(n248), .Y(n579) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n71), .C(\mem<2><2> ), .D(n228), .Y(n578) );
  AOI21X1 U857 ( .A(n580), .B(n581), .C(n970), .Y(n575) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n91), .C(\mem<4><2> ), .D(n248), .Y(n581) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n71), .C(\mem<6><2> ), .D(n228), .Y(n580) );
  AOI22X1 U860 ( .A(n288), .B(n879), .C(n249), .D(n919), .Y(n573) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n91), .C(\mem<12><2> ), .D(n248), .Y(
        n585) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n71), .C(\mem<14><2> ), .D(n228), .Y(
        n584) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n91), .C(\mem<8><2> ), .D(n248), .Y(n587) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n71), .C(\mem<10><2> ), .D(n228), .Y(
        n586) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n588) );
  NOR2X1 U868 ( .A(n1033), .B(\addr_1c<4> ), .Y(n589) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n590) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n199), .C(\mem<19><0> ), .D(n179), .Y(
        n597) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n160), .C(\mem<23><0> ), .D(n140), .Y(
        n596) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n121), .C(\mem<27><0> ), .D(n101), .Y(
        n594) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n81), .C(\mem<31><0> ), .D(n60), .Y(n593) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n357), .C(\mem<3><0> ), .D(n338), .Y(n604) );
  NAND2X1 U877 ( .A(n1031), .B(n1032), .Y(n367) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n318), .C(\mem<7><0> ), .D(n299), .Y(n603) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1032), .Y(n328) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n278), .C(\mem<11><0> ), .D(n259), .Y(
        n601) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n238), .C(\mem<15><0> ), .D(n218), .Y(
        n600) );
  dff_203 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1016) );
  dff_202 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1016) );
  dff_185 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1016)
         );
  dff_186 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1016)
         );
  dff_187 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1016)
         );
  dff_188 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1016)
         );
  dff_189 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1016)
         );
  dff_190 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1016)
         );
  dff_191 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1016)
         );
  dff_192 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1016)
         );
  dff_193 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1016)
         );
  dff_194 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1016)
         );
  dff_195 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1016) );
  dff_196 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1016) );
  dff_197 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1016) );
  dff_169 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1015) );
  dff_170 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1015) );
  dff_171 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1015) );
  dff_172 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1015) );
  dff_173 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1015) );
  dff_174 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1015) );
  dff_175 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1015) );
  dff_176 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1015) );
  dff_177 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1016) );
  dff_178 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1015) );
  dff_179 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1016) );
  dff_180 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1015) );
  dff_181 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1016) );
  dff_182 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1015) );
  dff_183 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1016) );
  dff_184 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1015) );
  dff_153 \reg2[0]  ( .q(\data_out<0> ), .d(n1028), .clk(clk), .rst(n1016) );
  dff_154 \reg2[1]  ( .q(\data_out<1> ), .d(n1027), .clk(clk), .rst(n1016) );
  dff_155 \reg2[2]  ( .q(\data_out<2> ), .d(n1026), .clk(clk), .rst(n1016) );
  dff_156 \reg2[3]  ( .q(\data_out<3> ), .d(n1025), .clk(clk), .rst(n1016) );
  dff_157 \reg2[4]  ( .q(\data_out<4> ), .d(n1024), .clk(clk), .rst(n1016) );
  dff_158 \reg2[5]  ( .q(\data_out<5> ), .d(n1023), .clk(clk), .rst(n1016) );
  dff_159 \reg2[6]  ( .q(\data_out<6> ), .d(n1022), .clk(clk), .rst(n1016) );
  dff_160 \reg2[7]  ( .q(\data_out<7> ), .d(n1021), .clk(clk), .rst(n1016) );
  dff_161 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1016) );
  dff_162 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1016) );
  dff_163 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1016) );
  dff_164 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1016) );
  dff_165 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1016) );
  dff_166 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1016) );
  dff_167 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1016) );
  dff_168 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1016) );
  dff_201 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1016) );
  dff_200 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1016) );
  dff_199 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1016) );
  dff_198 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1016) );
  INVX1 U2 ( .A(rd), .Y(n1019) );
  INVX1 U3 ( .A(rst), .Y(n1017) );
  OR2X1 U4 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n371) );
  AND2X1 U5 ( .A(\addr_1c<4> ), .B(n357), .Y(n49) );
  INVX1 U6 ( .A(n1017), .Y(n1015) );
  INVX1 U7 ( .A(\addr_1c<3> ), .Y(n1033) );
  INVX1 U8 ( .A(\addr_1c<2> ), .Y(n1032) );
  INVX1 U23 ( .A(\addr_1c<1> ), .Y(n1031) );
  OR2X1 U24 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n370) );
  AND2X1 U25 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n598) );
  AND2X1 U26 ( .A(\addr_1c<3> ), .B(n1030), .Y(n599) );
  AND2X1 U27 ( .A(n249), .B(n965), .Y(n70) );
  AND2X1 U28 ( .A(n288), .B(n965), .Y(n111) );
  AND2X1 U29 ( .A(\addr_1c<0> ), .B(n1033), .Y(n605) );
  AND2X1 U35 ( .A(n1030), .B(n1033), .Y(n606) );
  INVX1 U36 ( .A(\addr_1c<0> ), .Y(n1030) );
  INVX1 U37 ( .A(wr1), .Y(n1029) );
  AND2X1 U38 ( .A(\addr_1c<2> ), .B(n1031), .Y(n288) );
  AND2X1 U39 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n249) );
  AND2X1 U40 ( .A(n599), .B(n249), .Y(n81) );
  AND2X1 U41 ( .A(n288), .B(n598), .Y(n101) );
  AND2X1 U42 ( .A(n288), .B(n599), .Y(n121) );
  AND2X1 U43 ( .A(n941), .B(n598), .Y(n140) );
  AND2X1 U44 ( .A(n941), .B(n599), .Y(n160) );
  AND2X1 U46 ( .A(n598), .B(n951), .Y(n179) );
  AND2X1 U47 ( .A(n599), .B(n951), .Y(n199) );
  AND2X1 U48 ( .A(n605), .B(n249), .Y(n218) );
  AND2X1 U49 ( .A(n249), .B(n606), .Y(n238) );
  AND2X1 U50 ( .A(n605), .B(n288), .Y(n259) );
  AND2X1 U51 ( .A(n288), .B(n606), .Y(n278) );
  AND2X1 U52 ( .A(n605), .B(n941), .Y(n299) );
  AND2X1 U53 ( .A(n941), .B(n606), .Y(n318) );
  OR2X1 U54 ( .A(n970), .B(n964), .Y(n968) );
  AND2X1 U55 ( .A(n605), .B(n951), .Y(n338) );
  OR2X1 U56 ( .A(n964), .B(n971), .Y(n966) );
  AND2X1 U57 ( .A(n49), .B(\mem<32><0> ), .Y(n395) );
  AND2X1 U58 ( .A(n49), .B(\mem<32><1> ), .Y(n380) );
  AND2X1 U59 ( .A(n49), .B(\mem<32><2> ), .Y(n576) );
  AND2X1 U60 ( .A(n49), .B(\mem<32><3> ), .Y(n561) );
  AND2X1 U61 ( .A(n49), .B(\mem<32><4> ), .Y(n546) );
  AND2X1 U62 ( .A(n49), .B(\mem<32><5> ), .Y(n531) );
  AND2X1 U63 ( .A(n49), .B(\mem<32><6> ), .Y(n516) );
  AND2X1 U64 ( .A(n49), .B(\mem<32><7> ), .Y(n501) );
  INVX1 U65 ( .A(rd1), .Y(n1020) );
  INVX1 U66 ( .A(n1017), .Y(n1016) );
  BUFX2 U67 ( .A(n961), .Y(n1010) );
  BUFX2 U68 ( .A(n961), .Y(n1009) );
  BUFX2 U69 ( .A(n960), .Y(n1007) );
  BUFX2 U70 ( .A(n960), .Y(n1006) );
  BUFX2 U71 ( .A(n959), .Y(n1004) );
  BUFX2 U72 ( .A(n959), .Y(n1003) );
  BUFX2 U73 ( .A(n958), .Y(n1001) );
  BUFX2 U74 ( .A(n958), .Y(n1000) );
  BUFX2 U75 ( .A(n957), .Y(n990) );
  BUFX2 U76 ( .A(n957), .Y(n989) );
  BUFX2 U77 ( .A(n956), .Y(n987) );
  BUFX2 U78 ( .A(n956), .Y(n986) );
  BUFX2 U79 ( .A(n955), .Y(n984) );
  BUFX2 U80 ( .A(n955), .Y(n983) );
  BUFX2 U81 ( .A(n954), .Y(n981) );
  BUFX2 U82 ( .A(n954), .Y(n980) );
  INVX1 U83 ( .A(\data_in_1c<0> ), .Y(n1034) );
  INVX1 U84 ( .A(\data_in_1c<1> ), .Y(n1035) );
  INVX1 U85 ( .A(\data_in_1c<2> ), .Y(n1036) );
  INVX1 U86 ( .A(\data_in_1c<3> ), .Y(n1037) );
  INVX1 U87 ( .A(\data_in_1c<4> ), .Y(n1038) );
  INVX1 U88 ( .A(\data_in_1c<5> ), .Y(n1039) );
  INVX1 U89 ( .A(\data_in_1c<6> ), .Y(n1040) );
  INVX1 U90 ( .A(\data_in_1c<7> ), .Y(n1041) );
  INVX1 U91 ( .A(\data_in_1c<8> ), .Y(n1042) );
  INVX1 U92 ( .A(\data_in_1c<9> ), .Y(n1043) );
  INVX1 U93 ( .A(\data_in_1c<10> ), .Y(n1044) );
  INVX1 U129 ( .A(\data_in_1c<11> ), .Y(n1045) );
  INVX1 U589 ( .A(\data_in_1c<12> ), .Y(n1046) );
  INVX1 U640 ( .A(\data_in_1c<13> ), .Y(n1047) );
  INVX1 U659 ( .A(\data_in_1c<14> ), .Y(n1048) );
  INVX1 U660 ( .A(\data_in_1c<15> ), .Y(n1049) );
  INVX1 U664 ( .A(wr), .Y(n1018) );
  INVX1 U666 ( .A(n590), .Y(n1028) );
  INVX1 U672 ( .A(n485), .Y(n1027) );
  INVX1 U675 ( .A(n472), .Y(n1026) );
  INVX1 U679 ( .A(n459), .Y(n1025) );
  INVX1 U682 ( .A(n446), .Y(n1024) );
  INVX1 U694 ( .A(n433), .Y(n1023) );
  INVX1 U697 ( .A(n420), .Y(n1022) );
  INVX1 U701 ( .A(n407), .Y(n1021) );
  INVX1 U706 ( .A(n48), .Y(n1014) );
  AND2X1 U712 ( .A(wr1), .B(n1017), .Y(n48) );
  INVX1 U717 ( .A(n1014), .Y(n1012) );
  INVX1 U723 ( .A(n1014), .Y(n1013) );
  AND2X1 U728 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U734 ( .A(n1), .Y(n2) );
  AND2X1 U739 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U745 ( .A(n3), .Y(n4) );
  AND2X1 U750 ( .A(n60), .B(n189), .Y(n5) );
  INVX1 U756 ( .A(n5), .Y(n6) );
  AND2X1 U761 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U767 ( .A(n7), .Y(n8) );
  OR2X1 U772 ( .A(n487), .B(n10), .Y(n9) );
  OR2X1 U786 ( .A(n474), .B(n486), .Y(n10) );
  OR2X1 U789 ( .A(n522), .B(n12), .Y(n11) );
  OR2X1 U801 ( .A(n507), .B(n508), .Y(n12) );
  OR2X1 U804 ( .A(n538), .B(n14), .Y(n13) );
  OR2X1 U816 ( .A(n523), .B(n537), .Y(n14) );
  OR2X1 U819 ( .A(n567), .B(n16), .Y(n15) );
  OR2X1 U831 ( .A(n552), .B(n553), .Y(n16) );
  OR2X1 U834 ( .A(n583), .B(n18), .Y(n17) );
  OR2X1 U846 ( .A(n568), .B(n582), .Y(n18) );
  OR2X1 U849 ( .A(n871), .B(n20), .Y(n19) );
  OR2X1 U861 ( .A(n591), .B(n592), .Y(n20) );
  OR2X1 U864 ( .A(n874), .B(n22), .Y(n21) );
  OR2X1 U870 ( .A(n872), .B(n873), .Y(n22) );
  OR2X1 U875 ( .A(n877), .B(n24), .Y(n23) );
  OR2X1 U882 ( .A(n875), .B(n876), .Y(n24) );
  OR2X1 U883 ( .A(n896), .B(n26), .Y(n25) );
  OR2X1 U884 ( .A(n894), .B(n895), .Y(n26) );
  OR2X1 U885 ( .A(n899), .B(n28), .Y(n27) );
  OR2X1 U886 ( .A(n897), .B(n898), .Y(n28) );
  OR2X1 U887 ( .A(n902), .B(n30), .Y(n29) );
  OR2X1 U888 ( .A(n900), .B(n901), .Y(n30) );
  OR2X1 U889 ( .A(n905), .B(n32), .Y(n31) );
  OR2X1 U890 ( .A(n903), .B(n904), .Y(n32) );
  OR2X1 U891 ( .A(n908), .B(n34), .Y(n33) );
  OR2X1 U892 ( .A(n906), .B(n907), .Y(n34) );
  OR2X1 U893 ( .A(n911), .B(n36), .Y(n35) );
  OR2X1 U894 ( .A(n909), .B(n910), .Y(n36) );
  OR2X1 U895 ( .A(n914), .B(n38), .Y(n37) );
  OR2X1 U896 ( .A(n912), .B(n913), .Y(n38) );
  OR2X1 U897 ( .A(n917), .B(n150), .Y(n50) );
  OR2X1 U898 ( .A(n915), .B(n916), .Y(n150) );
  AND2X1 U899 ( .A(n973), .B(n48), .Y(n189) );
  AND2X1 U900 ( .A(n48), .B(n357), .Y(n289) );
  AND2X1 U901 ( .A(n941), .B(n943), .Y(n348) );
  INVX1 U902 ( .A(n348), .Y(n372) );
  AND2X1 U903 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U904 ( .A(n379), .Y(n381) );
  AND2X1 U905 ( .A(n941), .B(n942), .Y(n386) );
  INVX1 U906 ( .A(n386), .Y(n387) );
  AND2X1 U907 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U908 ( .A(n401), .Y(n402) );
  BUFX2 U909 ( .A(n1050), .Y(err) );
  BUFX2 U910 ( .A(n573), .Y(n409) );
  BUFX2 U911 ( .A(n558), .Y(n421) );
  BUFX2 U912 ( .A(n543), .Y(n422) );
  BUFX2 U913 ( .A(n528), .Y(n434) );
  BUFX2 U914 ( .A(n513), .Y(n435) );
  BUFX2 U915 ( .A(n498), .Y(n447) );
  BUFX2 U916 ( .A(n392), .Y(n448) );
  BUFX2 U917 ( .A(n377), .Y(n460) );
  AND2X2 U918 ( .A(rd), .B(n374), .Y(n461) );
  INVX1 U919 ( .A(n461), .Y(n473) );
  INVX1 U920 ( .A(n602), .Y(n474) );
  INVX1 U921 ( .A(n601), .Y(n486) );
  INVX1 U922 ( .A(n600), .Y(n487) );
  INVX1 U923 ( .A(n495), .Y(n507) );
  INVX1 U924 ( .A(n494), .Y(n508) );
  INVX1 U925 ( .A(n493), .Y(n522) );
  INVX1 U926 ( .A(n482), .Y(n523) );
  INVX1 U927 ( .A(n481), .Y(n537) );
  INVX1 U928 ( .A(n480), .Y(n538) );
  INVX1 U929 ( .A(n469), .Y(n552) );
  INVX1 U930 ( .A(n468), .Y(n553) );
  INVX1 U931 ( .A(n467), .Y(n567) );
  INVX1 U932 ( .A(n456), .Y(n568) );
  INVX1 U933 ( .A(n455), .Y(n582) );
  INVX1 U934 ( .A(n454), .Y(n583) );
  INVX1 U935 ( .A(n443), .Y(n591) );
  INVX1 U936 ( .A(n442), .Y(n592) );
  INVX1 U937 ( .A(n441), .Y(n871) );
  INVX1 U938 ( .A(n430), .Y(n872) );
  INVX1 U939 ( .A(n429), .Y(n873) );
  INVX1 U940 ( .A(n428), .Y(n874) );
  INVX1 U941 ( .A(n417), .Y(n875) );
  INVX1 U942 ( .A(n416), .Y(n876) );
  INVX1 U943 ( .A(n415), .Y(n877) );
  AND2X2 U944 ( .A(n586), .B(n587), .Y(n878) );
  INVX1 U945 ( .A(n878), .Y(n879) );
  AND2X2 U946 ( .A(n571), .B(n572), .Y(n880) );
  INVX1 U947 ( .A(n880), .Y(n881) );
  AND2X2 U948 ( .A(n556), .B(n557), .Y(n882) );
  INVX1 U949 ( .A(n882), .Y(n883) );
  AND2X2 U950 ( .A(n541), .B(n542), .Y(n884) );
  INVX1 U951 ( .A(n884), .Y(n885) );
  AND2X2 U952 ( .A(n526), .B(n527), .Y(n886) );
  INVX1 U953 ( .A(n886), .Y(n887) );
  AND2X2 U954 ( .A(n511), .B(n512), .Y(n888) );
  INVX1 U955 ( .A(n888), .Y(n889) );
  AND2X2 U956 ( .A(n405), .B(n406), .Y(n890) );
  INVX1 U957 ( .A(n890), .Y(n891) );
  AND2X2 U958 ( .A(n390), .B(n391), .Y(n892) );
  INVX1 U959 ( .A(n892), .Y(n893) );
  INVX1 U960 ( .A(n595), .Y(n894) );
  INVX1 U961 ( .A(n594), .Y(n895) );
  INVX1 U962 ( .A(n593), .Y(n896) );
  INVX1 U963 ( .A(n490), .Y(n897) );
  INVX1 U964 ( .A(n489), .Y(n898) );
  INVX1 U965 ( .A(n488), .Y(n899) );
  INVX1 U966 ( .A(n477), .Y(n900) );
  INVX1 U967 ( .A(n476), .Y(n901) );
  INVX1 U968 ( .A(n475), .Y(n902) );
  INVX1 U969 ( .A(n464), .Y(n903) );
  INVX1 U970 ( .A(n463), .Y(n904) );
  INVX1 U971 ( .A(n462), .Y(n905) );
  INVX1 U972 ( .A(n451), .Y(n906) );
  INVX1 U973 ( .A(n450), .Y(n907) );
  INVX1 U974 ( .A(n449), .Y(n908) );
  INVX1 U975 ( .A(n438), .Y(n909) );
  INVX1 U976 ( .A(n437), .Y(n910) );
  INVX1 U977 ( .A(n436), .Y(n911) );
  INVX1 U978 ( .A(n425), .Y(n912) );
  INVX1 U979 ( .A(n424), .Y(n913) );
  INVX1 U980 ( .A(n423), .Y(n914) );
  INVX1 U981 ( .A(n412), .Y(n915) );
  INVX1 U982 ( .A(n411), .Y(n916) );
  INVX1 U983 ( .A(n410), .Y(n917) );
  AND2X2 U984 ( .A(n584), .B(n585), .Y(n918) );
  INVX1 U985 ( .A(n918), .Y(n919) );
  AND2X2 U986 ( .A(n569), .B(n570), .Y(n920) );
  INVX1 U987 ( .A(n920), .Y(n921) );
  AND2X2 U988 ( .A(n554), .B(n555), .Y(n922) );
  INVX1 U989 ( .A(n922), .Y(n923) );
  AND2X2 U990 ( .A(n539), .B(n540), .Y(n924) );
  INVX1 U991 ( .A(n924), .Y(n925) );
  AND2X2 U992 ( .A(n524), .B(n525), .Y(n926) );
  INVX1 U993 ( .A(n926), .Y(n927) );
  AND2X2 U994 ( .A(n509), .B(n510), .Y(n928) );
  INVX1 U995 ( .A(n928), .Y(n929) );
  AND2X2 U996 ( .A(n403), .B(n404), .Y(n930) );
  INVX1 U997 ( .A(n930), .Y(n931) );
  AND2X2 U998 ( .A(n388), .B(n389), .Y(n932) );
  INVX1 U999 ( .A(n932), .Y(n933) );
  BUFX2 U1000 ( .A(n575), .Y(n934) );
  BUFX2 U1001 ( .A(n560), .Y(n935) );
  BUFX2 U1002 ( .A(n545), .Y(n936) );
  BUFX2 U1003 ( .A(n530), .Y(n937) );
  BUFX2 U1004 ( .A(n515), .Y(n938) );
  BUFX2 U1005 ( .A(n500), .Y(n939) );
  BUFX2 U1006 ( .A(n394), .Y(n940) );
  INVX1 U1007 ( .A(n970), .Y(n941) );
  INVX1 U1008 ( .A(n385), .Y(n942) );
  INVX1 U1009 ( .A(n384), .Y(n943) );
  BUFX2 U1010 ( .A(n328), .Y(n970) );
  BUFX2 U1011 ( .A(n577), .Y(n944) );
  BUFX2 U1012 ( .A(n562), .Y(n945) );
  BUFX2 U1013 ( .A(n547), .Y(n946) );
  BUFX2 U1014 ( .A(n532), .Y(n947) );
  BUFX2 U1015 ( .A(n517), .Y(n948) );
  BUFX2 U1016 ( .A(n502), .Y(n949) );
  BUFX2 U1017 ( .A(n396), .Y(n950) );
  INVX1 U1018 ( .A(n971), .Y(n951) );
  INVX1 U1019 ( .A(n383), .Y(n952) );
  INVX1 U1020 ( .A(n382), .Y(n953) );
  BUFX2 U1021 ( .A(n367), .Y(n971) );
  BUFX2 U1022 ( .A(n358), .Y(n972) );
  BUFX2 U1023 ( .A(n339), .Y(n974) );
  BUFX2 U1024 ( .A(n329), .Y(n975) );
  BUFX2 U1025 ( .A(n319), .Y(n976) );
  BUFX2 U1026 ( .A(n309), .Y(n977) );
  BUFX2 U1027 ( .A(n300), .Y(n978) );
  BUFX2 U1028 ( .A(n290), .Y(n979) );
  BUFX2 U1029 ( .A(n269), .Y(n982) );
  BUFX2 U1030 ( .A(n250), .Y(n985) );
  BUFX2 U1031 ( .A(n229), .Y(n988) );
  BUFX2 U1032 ( .A(n209), .Y(n991) );
  BUFX2 U1033 ( .A(n200), .Y(n992) );
  BUFX2 U1034 ( .A(n190), .Y(n993) );
  BUFX2 U1035 ( .A(n180), .Y(n994) );
  BUFX2 U1036 ( .A(n170), .Y(n995) );
  BUFX2 U1037 ( .A(n161), .Y(n996) );
  BUFX2 U1038 ( .A(n151), .Y(n997) );
  BUFX2 U1039 ( .A(n141), .Y(n998) );
  BUFX2 U1040 ( .A(n131), .Y(n999) );
  BUFX2 U1041 ( .A(n112), .Y(n1002) );
  BUFX2 U1042 ( .A(n92), .Y(n1005) );
  BUFX2 U1043 ( .A(n72), .Y(n1008) );
  BUFX2 U1044 ( .A(n59), .Y(n973) );
  AND2X1 U1045 ( .A(n249), .B(n598), .Y(n60) );
  BUFX2 U1046 ( .A(n39), .Y(n1011) );
  BUFX2 U1047 ( .A(n279), .Y(n954) );
  BUFX2 U1048 ( .A(n260), .Y(n955) );
  BUFX2 U1049 ( .A(n239), .Y(n956) );
  BUFX2 U1050 ( .A(n219), .Y(n957) );
  BUFX2 U1051 ( .A(n122), .Y(n958) );
  BUFX2 U1052 ( .A(n102), .Y(n959) );
  BUFX2 U1053 ( .A(n82), .Y(n960) );
  BUFX2 U1054 ( .A(n61), .Y(n961) );
  AND2X1 U1055 ( .A(enable), .B(n1017), .Y(n962) );
  INVX1 U1056 ( .A(n962), .Y(n963) );
  INVX1 U1057 ( .A(n965), .Y(n964) );
  AND2X1 U1058 ( .A(n368), .B(n369), .Y(n965) );
  INVX1 U1059 ( .A(n966), .Y(n967) );
  INVX1 U1060 ( .A(n968), .Y(n969) );
  AND2X1 U1061 ( .A(n951), .B(n606), .Y(n357) );
endmodule


module final_memory_2 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1842, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1050), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1051), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1052), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1053), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1054), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1055), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1056), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1057), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1058), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1059), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1060), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1061), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1062), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1063), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1064), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1065), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1066), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1067), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1068), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1069), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1070), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1071), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1072), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1073), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1074), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1075), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1076), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1077), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1078), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1079), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1080), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1081), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1082), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1083), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1084), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1085), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1086), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1087), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1088), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1089), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1090), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1091), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1092), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1093), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1094), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1095), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1096), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1097), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1098), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1099), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1100), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1101), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1102), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1103), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1104), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1105), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1106), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1107), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1108), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1109), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1110), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1111), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1112), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1113), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1114), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1115), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1116), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1117), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1118), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1119), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1120), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1121), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1122), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1123), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1124), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1125), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1126), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1127), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1128), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1129), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1130), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1131), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1132), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1133), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1134), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1135), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1136), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1137), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1138), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1139), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1140), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1141), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1142), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1143), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1144), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1145), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1146), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1147), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1148), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1149), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1150), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1151), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1152), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1153), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1154), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1155), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1156), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1157), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1158), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1159), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1160), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1161), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1162), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1163), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1164), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1165), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1166), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1167), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1168), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1169), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1170), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1171), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1172), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1173), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1174), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1175), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1176), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1177), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1178), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1179), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1180), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1181), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1182), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1183), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1184), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1185), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1186), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1187), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1188), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1189), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1190), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1191), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1192), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1193), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1194), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1195), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1196), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1197), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1198), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1199), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1200), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1201), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1202), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1203), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1204), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1205), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1206), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1207), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1208), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1209), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1210), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1211), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1212), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1213), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1214), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1215), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1216), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1217), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1218), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1219), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1220), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1221), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1222), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1223), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1224), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1225), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1226), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1227), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1228), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1229), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1230), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1231), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1232), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1233), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1234), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1235), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1236), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1237), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1238), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1239), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1240), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1241), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1242), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1243), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1244), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1245), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1246), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1247), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1248), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1249), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1250), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1251), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1252), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1253), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1254), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1255), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1256), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1257), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1258), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1259), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1260), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1261), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1262), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1263), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1264), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1265), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1266), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1267), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1268), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1269), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1270), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1271), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1272), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1273), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1274), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1275), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1276), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1277), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1278), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1279), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1280), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1281), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1282), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1283), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1284), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1285), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1286), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1287), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1288), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1289), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1290), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1291), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1292), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1293), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1294), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1295), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1296), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1297), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1298), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1299), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1300), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1301), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1302), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1303), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1304), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1305), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1306), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1307), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1308), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1309), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1310), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1311), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1312), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1313), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1481), .B(n1480), .Y(n1482) );
  AND2X2 U10 ( .A(n1476), .B(n1475), .Y(n1477) );
  AND2X2 U11 ( .A(n1470), .B(n1469), .Y(n1471) );
  AND2X2 U12 ( .A(n1465), .B(n1464), .Y(n1466) );
  AND2X2 U13 ( .A(n1459), .B(n1458), .Y(n1460) );
  AND2X2 U14 ( .A(n1454), .B(n1453), .Y(n1455) );
  AND2X2 U15 ( .A(n1448), .B(n1447), .Y(n1449) );
  AND2X2 U16 ( .A(n1443), .B(n1442), .Y(n1444) );
  AND2X2 U17 ( .A(n1437), .B(n1436), .Y(n1438) );
  AND2X2 U18 ( .A(n1432), .B(n1431), .Y(n1433) );
  AND2X2 U19 ( .A(n1426), .B(n1425), .Y(n1427) );
  AND2X2 U20 ( .A(n1421), .B(n1420), .Y(n1422) );
  AND2X2 U21 ( .A(n1415), .B(n1414), .Y(n1416) );
  AND2X2 U22 ( .A(n1410), .B(n1409), .Y(n1411) );
  AND2X2 U30 ( .A(n1330), .B(n1030), .Y(n1635) );
  AND2X2 U31 ( .A(n1329), .B(n1030), .Y(n1790) );
  AND2X2 U32 ( .A(n1330), .B(\addr_1c<0> ), .Y(n1655) );
  AND2X2 U33 ( .A(n1329), .B(\addr_1c<0> ), .Y(n1810) );
  AND2X2 U34 ( .A(n1324), .B(n1323), .Y(n1325) );
  AND2X2 U45 ( .A(n1317), .B(n1316), .Y(n1318) );
  NOR3X1 U94 ( .A(n1026), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1027), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1042), .C(n1840), .Y(n1313) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1840) );
  OAI21X1 U98 ( .A(n1011), .B(n1043), .C(n1839), .Y(n1312) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1839) );
  OAI21X1 U100 ( .A(n1011), .B(n1044), .C(n1838), .Y(n1311) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1838) );
  OAI21X1 U102 ( .A(n1011), .B(n1045), .C(n1837), .Y(n1310) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1837) );
  OAI21X1 U104 ( .A(n1011), .B(n1046), .C(n1836), .Y(n1309) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1836) );
  OAI21X1 U106 ( .A(n1011), .B(n1047), .C(n1835), .Y(n1308) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1835) );
  OAI21X1 U108 ( .A(n1011), .B(n1048), .C(n1834), .Y(n1307) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1834) );
  OAI21X1 U110 ( .A(n1011), .B(n1049), .C(n1833), .Y(n1306) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1833) );
  NAND3X1 U112 ( .A(n1012), .B(n1831), .C(n965), .Y(n1841) );
  OAI21X1 U113 ( .A(n6), .B(n1034), .C(n1830), .Y(n1305) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1830) );
  OAI21X1 U115 ( .A(n6), .B(n1035), .C(n1829), .Y(n1304) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1829) );
  OAI21X1 U117 ( .A(n6), .B(n1036), .C(n1828), .Y(n1303) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1828) );
  OAI21X1 U119 ( .A(n6), .B(n1037), .C(n1827), .Y(n1302) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1827) );
  OAI21X1 U121 ( .A(n6), .B(n1038), .C(n1826), .Y(n1301) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1826) );
  OAI21X1 U123 ( .A(n6), .B(n1039), .C(n1825), .Y(n1300) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1825) );
  OAI21X1 U125 ( .A(n6), .B(n1040), .C(n1824), .Y(n1299) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1824) );
  OAI21X1 U127 ( .A(n6), .B(n1041), .C(n1823), .Y(n1298) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1823) );
  OAI21X1 U130 ( .A(n1042), .B(n1010), .C(n1819), .Y(n1297) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1819) );
  OAI21X1 U132 ( .A(n1043), .B(n1009), .C(n1818), .Y(n1296) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1818) );
  OAI21X1 U134 ( .A(n1044), .B(n1009), .C(n1817), .Y(n1295) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1817) );
  OAI21X1 U136 ( .A(n1045), .B(n1009), .C(n1816), .Y(n1294) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1816) );
  OAI21X1 U138 ( .A(n1046), .B(n1009), .C(n1815), .Y(n1293) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1815) );
  OAI21X1 U140 ( .A(n1047), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1814) );
  OAI21X1 U142 ( .A(n1048), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1813) );
  OAI21X1 U144 ( .A(n1049), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1812) );
  NAND3X1 U146 ( .A(n1811), .B(n1832), .C(n1810), .Y(n1820) );
  OAI21X1 U147 ( .A(n1034), .B(n1008), .C(n1808), .Y(n1289) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1808) );
  OAI21X1 U149 ( .A(n1035), .B(n1008), .C(n1807), .Y(n1288) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1807) );
  OAI21X1 U151 ( .A(n1036), .B(n1008), .C(n1806), .Y(n1287) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1806) );
  OAI21X1 U153 ( .A(n1037), .B(n1008), .C(n1805), .Y(n1286) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1805) );
  OAI21X1 U155 ( .A(n1038), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1804) );
  OAI21X1 U157 ( .A(n1039), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1803) );
  OAI21X1 U159 ( .A(n1040), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1802) );
  OAI21X1 U161 ( .A(n1041), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1801) );
  NAND3X1 U163 ( .A(n973), .B(n1013), .C(n1800), .Y(n1809) );
  OAI21X1 U164 ( .A(n1042), .B(n1007), .C(n1798), .Y(n1281) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1798) );
  OAI21X1 U166 ( .A(n1043), .B(n1006), .C(n1797), .Y(n1280) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1797) );
  OAI21X1 U168 ( .A(n1044), .B(n1006), .C(n1796), .Y(n1279) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1796) );
  OAI21X1 U170 ( .A(n1045), .B(n1006), .C(n1795), .Y(n1278) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1795) );
  OAI21X1 U172 ( .A(n1046), .B(n1006), .C(n1794), .Y(n1277) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1794) );
  OAI21X1 U174 ( .A(n1047), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1793) );
  OAI21X1 U176 ( .A(n1048), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1792) );
  OAI21X1 U178 ( .A(n1049), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1791) );
  NAND3X1 U180 ( .A(n1811), .B(n1832), .C(n1790), .Y(n1799) );
  OAI21X1 U181 ( .A(n1034), .B(n1005), .C(n1788), .Y(n1273) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1788) );
  OAI21X1 U183 ( .A(n1035), .B(n1005), .C(n1787), .Y(n1272) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1787) );
  OAI21X1 U185 ( .A(n1036), .B(n1005), .C(n1786), .Y(n1271) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1786) );
  OAI21X1 U187 ( .A(n1037), .B(n1005), .C(n1785), .Y(n1270) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1785) );
  OAI21X1 U189 ( .A(n1038), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1784) );
  OAI21X1 U191 ( .A(n1039), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1783) );
  OAI21X1 U193 ( .A(n1040), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1782) );
  OAI21X1 U195 ( .A(n1041), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1781) );
  NAND3X1 U197 ( .A(n973), .B(n1012), .C(n1780), .Y(n1789) );
  OAI21X1 U198 ( .A(n1042), .B(n1004), .C(n1778), .Y(n1265) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1778) );
  OAI21X1 U200 ( .A(n1043), .B(n1003), .C(n1777), .Y(n1264) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1777) );
  OAI21X1 U202 ( .A(n1044), .B(n1003), .C(n1776), .Y(n1263) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1776) );
  OAI21X1 U204 ( .A(n1045), .B(n1003), .C(n1775), .Y(n1262) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1775) );
  OAI21X1 U206 ( .A(n1046), .B(n1003), .C(n1774), .Y(n1261) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1774) );
  OAI21X1 U208 ( .A(n1047), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1773) );
  OAI21X1 U210 ( .A(n1048), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1772) );
  OAI21X1 U212 ( .A(n1049), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1771) );
  NAND3X1 U214 ( .A(n1810), .B(n1013), .C(n1770), .Y(n1779) );
  OAI21X1 U215 ( .A(n1034), .B(n1002), .C(n1768), .Y(n1257) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1768) );
  OAI21X1 U217 ( .A(n1035), .B(n1002), .C(n1767), .Y(n1256) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1767) );
  OAI21X1 U219 ( .A(n1036), .B(n1002), .C(n1766), .Y(n1255) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1766) );
  OAI21X1 U221 ( .A(n1037), .B(n1002), .C(n1765), .Y(n1254) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1765) );
  OAI21X1 U223 ( .A(n1038), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1764) );
  OAI21X1 U225 ( .A(n1039), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1763) );
  OAI21X1 U227 ( .A(n1040), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1762) );
  OAI21X1 U229 ( .A(n1041), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1761) );
  NAND3X1 U231 ( .A(n973), .B(n1013), .C(n1760), .Y(n1769) );
  OAI21X1 U232 ( .A(n1042), .B(n1001), .C(n1758), .Y(n1249) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1758) );
  OAI21X1 U234 ( .A(n1043), .B(n1000), .C(n1757), .Y(n1248) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1757) );
  OAI21X1 U236 ( .A(n1044), .B(n1000), .C(n1756), .Y(n1247) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1756) );
  OAI21X1 U238 ( .A(n1045), .B(n1000), .C(n1755), .Y(n1246) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1755) );
  OAI21X1 U240 ( .A(n1046), .B(n1000), .C(n1754), .Y(n1245) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1754) );
  OAI21X1 U242 ( .A(n1047), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1753) );
  OAI21X1 U244 ( .A(n1048), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1752) );
  OAI21X1 U246 ( .A(n1049), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1751) );
  NAND3X1 U248 ( .A(n1790), .B(n1013), .C(n1770), .Y(n1759) );
  OAI21X1 U249 ( .A(n1034), .B(n999), .C(n1749), .Y(n1241) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1749) );
  OAI21X1 U251 ( .A(n1035), .B(n999), .C(n1748), .Y(n1240) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1748) );
  OAI21X1 U253 ( .A(n1036), .B(n999), .C(n1747), .Y(n1239) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1747) );
  OAI21X1 U255 ( .A(n1037), .B(n999), .C(n1746), .Y(n1238) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1746) );
  OAI21X1 U257 ( .A(n1038), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1745) );
  OAI21X1 U259 ( .A(n1039), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1744) );
  OAI21X1 U261 ( .A(n1040), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1743) );
  OAI21X1 U263 ( .A(n1041), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1742) );
  NAND3X1 U265 ( .A(n973), .B(n1013), .C(n1741), .Y(n1750) );
  OAI21X1 U266 ( .A(n1042), .B(n998), .C(n1739), .Y(n1233) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1739) );
  OAI21X1 U268 ( .A(n1043), .B(n998), .C(n1738), .Y(n1232) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1738) );
  OAI21X1 U270 ( .A(n1044), .B(n998), .C(n1737), .Y(n1231) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1737) );
  OAI21X1 U272 ( .A(n1045), .B(n998), .C(n1736), .Y(n1230) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1736) );
  OAI21X1 U274 ( .A(n1046), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1735) );
  OAI21X1 U276 ( .A(n1047), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1734) );
  OAI21X1 U278 ( .A(n1048), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1733) );
  OAI21X1 U280 ( .A(n1049), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1732) );
  NAND3X1 U282 ( .A(n1810), .B(n1013), .C(n969), .Y(n1740) );
  OAI21X1 U283 ( .A(n1034), .B(n997), .C(n1730), .Y(n1225) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1730) );
  OAI21X1 U285 ( .A(n1035), .B(n997), .C(n1729), .Y(n1224) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1729) );
  OAI21X1 U287 ( .A(n1036), .B(n997), .C(n1728), .Y(n1223) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1728) );
  OAI21X1 U289 ( .A(n1037), .B(n997), .C(n1727), .Y(n1222) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1727) );
  OAI21X1 U291 ( .A(n1038), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1726) );
  OAI21X1 U293 ( .A(n1039), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1725) );
  OAI21X1 U295 ( .A(n1040), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1724) );
  OAI21X1 U297 ( .A(n1041), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1723) );
  NAND3X1 U299 ( .A(n973), .B(n1013), .C(n1722), .Y(n1731) );
  OAI21X1 U300 ( .A(n1042), .B(n996), .C(n1720), .Y(n1217) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1720) );
  OAI21X1 U302 ( .A(n1043), .B(n996), .C(n1719), .Y(n1216) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1719) );
  OAI21X1 U304 ( .A(n1044), .B(n996), .C(n1718), .Y(n1215) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1718) );
  OAI21X1 U306 ( .A(n1045), .B(n996), .C(n1717), .Y(n1214) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1717) );
  OAI21X1 U308 ( .A(n1046), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1716) );
  OAI21X1 U310 ( .A(n1047), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1715) );
  OAI21X1 U312 ( .A(n1048), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1714) );
  OAI21X1 U314 ( .A(n1049), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1713) );
  NAND3X1 U316 ( .A(n1790), .B(n1013), .C(n969), .Y(n1721) );
  OAI21X1 U317 ( .A(n1034), .B(n995), .C(n1711), .Y(n1209) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1711) );
  OAI21X1 U319 ( .A(n1035), .B(n995), .C(n1710), .Y(n1208) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1710) );
  OAI21X1 U321 ( .A(n1036), .B(n995), .C(n1709), .Y(n1207) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1709) );
  OAI21X1 U323 ( .A(n1037), .B(n995), .C(n1708), .Y(n1206) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1708) );
  OAI21X1 U325 ( .A(n1038), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1707) );
  OAI21X1 U327 ( .A(n1039), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1706) );
  OAI21X1 U329 ( .A(n1040), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1705) );
  OAI21X1 U331 ( .A(n1041), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1704) );
  NAND3X1 U333 ( .A(n973), .B(n1013), .C(n1703), .Y(n1712) );
  OAI21X1 U334 ( .A(n1042), .B(n994), .C(n1701), .Y(n1201) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1701) );
  OAI21X1 U336 ( .A(n1043), .B(n994), .C(n1700), .Y(n1200) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1700) );
  OAI21X1 U338 ( .A(n1044), .B(n994), .C(n1699), .Y(n1199) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1699) );
  OAI21X1 U340 ( .A(n1045), .B(n994), .C(n1698), .Y(n1198) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1698) );
  OAI21X1 U342 ( .A(n1046), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1697) );
  OAI21X1 U344 ( .A(n1047), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1696) );
  OAI21X1 U346 ( .A(n1048), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1695) );
  OAI21X1 U348 ( .A(n1049), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1694) );
  NAND3X1 U350 ( .A(n1810), .B(n1013), .C(n967), .Y(n1702) );
  OAI21X1 U351 ( .A(n1034), .B(n993), .C(n1692), .Y(n1193) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1692) );
  OAI21X1 U353 ( .A(n1035), .B(n993), .C(n1691), .Y(n1192) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1691) );
  OAI21X1 U355 ( .A(n1036), .B(n993), .C(n1690), .Y(n1191) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1690) );
  OAI21X1 U357 ( .A(n1037), .B(n993), .C(n1689), .Y(n1190) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1689) );
  OAI21X1 U359 ( .A(n1038), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1688) );
  OAI21X1 U361 ( .A(n1039), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1687) );
  OAI21X1 U363 ( .A(n1040), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1686) );
  OAI21X1 U365 ( .A(n1041), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1685) );
  NAND3X1 U367 ( .A(n973), .B(n1013), .C(n1684), .Y(n1693) );
  OAI21X1 U368 ( .A(n1042), .B(n992), .C(n1682), .Y(n1185) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1682) );
  OAI21X1 U370 ( .A(n1043), .B(n992), .C(n1681), .Y(n1184) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1681) );
  OAI21X1 U372 ( .A(n1044), .B(n992), .C(n1680), .Y(n1183) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1680) );
  OAI21X1 U374 ( .A(n1045), .B(n992), .C(n1679), .Y(n1182) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1679) );
  OAI21X1 U376 ( .A(n1046), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1678) );
  OAI21X1 U378 ( .A(n1047), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1677) );
  OAI21X1 U380 ( .A(n1048), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1676) );
  OAI21X1 U382 ( .A(n1049), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1675) );
  NAND3X1 U384 ( .A(n1790), .B(n1013), .C(n967), .Y(n1683) );
  OAI21X1 U385 ( .A(n1034), .B(n991), .C(n1673), .Y(n1177) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1673) );
  OAI21X1 U387 ( .A(n1035), .B(n991), .C(n1672), .Y(n1176) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1672) );
  OAI21X1 U389 ( .A(n1036), .B(n991), .C(n1671), .Y(n1175) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1671) );
  OAI21X1 U391 ( .A(n1037), .B(n991), .C(n1670), .Y(n1174) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1670) );
  OAI21X1 U393 ( .A(n1038), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1669) );
  OAI21X1 U395 ( .A(n1039), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1668) );
  OAI21X1 U397 ( .A(n1040), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1667) );
  OAI21X1 U399 ( .A(n1041), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1666) );
  NAND3X1 U401 ( .A(n973), .B(n1013), .C(n1665), .Y(n1674) );
  OAI21X1 U402 ( .A(n1042), .B(n990), .C(n1663), .Y(n1169) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1663) );
  OAI21X1 U404 ( .A(n1043), .B(n989), .C(n1662), .Y(n1168) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1662) );
  OAI21X1 U406 ( .A(n1044), .B(n989), .C(n1661), .Y(n1167) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1661) );
  OAI21X1 U408 ( .A(n1045), .B(n989), .C(n1660), .Y(n1166) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1660) );
  OAI21X1 U410 ( .A(n1046), .B(n989), .C(n1659), .Y(n1165) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1659) );
  OAI21X1 U412 ( .A(n1047), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1658) );
  OAI21X1 U414 ( .A(n1048), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1657) );
  OAI21X1 U416 ( .A(n1049), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1656) );
  NAND3X1 U418 ( .A(n1811), .B(n1012), .C(n1655), .Y(n1664) );
  OAI21X1 U419 ( .A(n1034), .B(n988), .C(n1653), .Y(n1161) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1653) );
  OAI21X1 U421 ( .A(n1035), .B(n988), .C(n1652), .Y(n1160) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1652) );
  OAI21X1 U423 ( .A(n1036), .B(n988), .C(n1651), .Y(n1159) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1651) );
  OAI21X1 U425 ( .A(n1037), .B(n988), .C(n1650), .Y(n1158) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1650) );
  OAI21X1 U427 ( .A(n1038), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1649) );
  OAI21X1 U429 ( .A(n1039), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1648) );
  OAI21X1 U431 ( .A(n1040), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1647) );
  OAI21X1 U433 ( .A(n1041), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1646) );
  NAND3X1 U435 ( .A(n973), .B(n1012), .C(n1645), .Y(n1654) );
  OAI21X1 U436 ( .A(n1042), .B(n987), .C(n1643), .Y(n1153) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1643) );
  OAI21X1 U438 ( .A(n1043), .B(n986), .C(n1642), .Y(n1152) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1642) );
  OAI21X1 U440 ( .A(n1044), .B(n986), .C(n1641), .Y(n1151) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1641) );
  OAI21X1 U442 ( .A(n1045), .B(n986), .C(n1640), .Y(n1150) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1640) );
  OAI21X1 U444 ( .A(n1046), .B(n986), .C(n1639), .Y(n1149) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1639) );
  OAI21X1 U446 ( .A(n1047), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1638) );
  OAI21X1 U448 ( .A(n1048), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1637) );
  OAI21X1 U450 ( .A(n1049), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1636) );
  NAND3X1 U452 ( .A(n1811), .B(n1012), .C(n1635), .Y(n1644) );
  OAI21X1 U453 ( .A(n1034), .B(n985), .C(n1632), .Y(n1145) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1632) );
  OAI21X1 U455 ( .A(n1035), .B(n985), .C(n1631), .Y(n1144) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1631) );
  OAI21X1 U457 ( .A(n1036), .B(n985), .C(n1630), .Y(n1143) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1630) );
  OAI21X1 U459 ( .A(n1037), .B(n985), .C(n1629), .Y(n1142) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1629) );
  OAI21X1 U461 ( .A(n1038), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1628) );
  OAI21X1 U463 ( .A(n1039), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1627) );
  OAI21X1 U465 ( .A(n1040), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1626) );
  OAI21X1 U467 ( .A(n1041), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1625) );
  NAND3X1 U469 ( .A(n973), .B(n1012), .C(n1624), .Y(n1633) );
  OAI21X1 U470 ( .A(n1042), .B(n984), .C(n1622), .Y(n1137) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1622) );
  OAI21X1 U472 ( .A(n1043), .B(n983), .C(n1621), .Y(n1136) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1621) );
  OAI21X1 U474 ( .A(n1044), .B(n983), .C(n1620), .Y(n1135) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1620) );
  OAI21X1 U476 ( .A(n1045), .B(n983), .C(n1619), .Y(n1134) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1619) );
  OAI21X1 U478 ( .A(n1046), .B(n983), .C(n1618), .Y(n1133) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1618) );
  OAI21X1 U480 ( .A(n1047), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1617) );
  OAI21X1 U482 ( .A(n1048), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1616) );
  OAI21X1 U484 ( .A(n1049), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1615) );
  NAND3X1 U486 ( .A(n1770), .B(n1012), .C(n1655), .Y(n1623) );
  OAI21X1 U487 ( .A(n1034), .B(n982), .C(n1613), .Y(n1129) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1613) );
  OAI21X1 U489 ( .A(n1035), .B(n982), .C(n1612), .Y(n1128) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1612) );
  OAI21X1 U491 ( .A(n1036), .B(n982), .C(n1611), .Y(n1127) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1611) );
  OAI21X1 U493 ( .A(n1037), .B(n982), .C(n1610), .Y(n1126) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1610) );
  OAI21X1 U495 ( .A(n1038), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1609) );
  OAI21X1 U497 ( .A(n1039), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1608) );
  OAI21X1 U499 ( .A(n1040), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1607) );
  OAI21X1 U501 ( .A(n1041), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1606) );
  NAND3X1 U503 ( .A(n973), .B(n1012), .C(n1605), .Y(n1614) );
  OAI21X1 U504 ( .A(n1042), .B(n981), .C(n1603), .Y(n1121) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1603) );
  OAI21X1 U506 ( .A(n1043), .B(n980), .C(n1602), .Y(n1120) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1602) );
  OAI21X1 U508 ( .A(n1044), .B(n980), .C(n1601), .Y(n1119) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1601) );
  OAI21X1 U510 ( .A(n1045), .B(n980), .C(n1600), .Y(n1118) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1600) );
  OAI21X1 U512 ( .A(n1046), .B(n980), .C(n1599), .Y(n1117) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1599) );
  OAI21X1 U514 ( .A(n1047), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1598) );
  OAI21X1 U516 ( .A(n1048), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1597) );
  OAI21X1 U518 ( .A(n1049), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1596) );
  NAND3X1 U520 ( .A(n1770), .B(n1012), .C(n1635), .Y(n1604) );
  OAI21X1 U521 ( .A(n1034), .B(n979), .C(n1593), .Y(n1113) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1593) );
  OAI21X1 U523 ( .A(n1035), .B(n979), .C(n1592), .Y(n1112) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1592) );
  OAI21X1 U525 ( .A(n1036), .B(n979), .C(n1591), .Y(n1111) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1591) );
  OAI21X1 U527 ( .A(n1037), .B(n979), .C(n1590), .Y(n1110) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1590) );
  OAI21X1 U529 ( .A(n1038), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1589) );
  OAI21X1 U531 ( .A(n1039), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1588) );
  OAI21X1 U533 ( .A(n1040), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1587) );
  OAI21X1 U535 ( .A(n1041), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1586) );
  NAND3X1 U537 ( .A(n973), .B(n1012), .C(n1585), .Y(n1594) );
  OAI21X1 U538 ( .A(n1042), .B(n978), .C(n1583), .Y(n1105) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1583) );
  OAI21X1 U540 ( .A(n1043), .B(n978), .C(n1582), .Y(n1104) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1582) );
  OAI21X1 U542 ( .A(n1044), .B(n978), .C(n1581), .Y(n1103) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1581) );
  OAI21X1 U544 ( .A(n1045), .B(n978), .C(n1580), .Y(n1102) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1580) );
  OAI21X1 U546 ( .A(n1046), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1579) );
  OAI21X1 U548 ( .A(n1047), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1578) );
  OAI21X1 U550 ( .A(n1048), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1577) );
  OAI21X1 U552 ( .A(n1049), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1576) );
  NAND3X1 U554 ( .A(n969), .B(n1012), .C(n1655), .Y(n1584) );
  OAI21X1 U555 ( .A(n1034), .B(n977), .C(n1574), .Y(n1097) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1574) );
  OAI21X1 U557 ( .A(n1035), .B(n977), .C(n1573), .Y(n1096) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1573) );
  OAI21X1 U559 ( .A(n1036), .B(n977), .C(n1572), .Y(n1095) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1572) );
  OAI21X1 U561 ( .A(n1037), .B(n977), .C(n1571), .Y(n1094) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1571) );
  OAI21X1 U563 ( .A(n1038), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1570) );
  OAI21X1 U565 ( .A(n1039), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1569) );
  OAI21X1 U567 ( .A(n1040), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1568) );
  OAI21X1 U569 ( .A(n1041), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1567) );
  NAND3X1 U571 ( .A(n973), .B(n1012), .C(n1566), .Y(n1575) );
  OAI21X1 U572 ( .A(n1042), .B(n976), .C(n1564), .Y(n1089) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1564) );
  OAI21X1 U574 ( .A(n1043), .B(n976), .C(n1563), .Y(n1088) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1563) );
  OAI21X1 U576 ( .A(n1044), .B(n976), .C(n1562), .Y(n1087) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1562) );
  OAI21X1 U578 ( .A(n1045), .B(n976), .C(n1561), .Y(n1086) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1561) );
  OAI21X1 U580 ( .A(n1046), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1560) );
  OAI21X1 U582 ( .A(n1047), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1559) );
  OAI21X1 U584 ( .A(n1048), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1558) );
  OAI21X1 U586 ( .A(n1049), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1557) );
  NAND3X1 U588 ( .A(n969), .B(n1012), .C(n1635), .Y(n1565) );
  OAI21X1 U590 ( .A(n1034), .B(n975), .C(n1554), .Y(n1081) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1554) );
  OAI21X1 U592 ( .A(n1035), .B(n975), .C(n1553), .Y(n1080) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1553) );
  OAI21X1 U594 ( .A(n1036), .B(n975), .C(n1552), .Y(n1079) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1552) );
  OAI21X1 U596 ( .A(n1037), .B(n975), .C(n1551), .Y(n1078) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1551) );
  OAI21X1 U598 ( .A(n1038), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1550) );
  OAI21X1 U600 ( .A(n1039), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1549) );
  OAI21X1 U602 ( .A(n1040), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1548) );
  OAI21X1 U604 ( .A(n1041), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1547) );
  NAND3X1 U606 ( .A(n973), .B(n1012), .C(n1546), .Y(n1555) );
  OAI21X1 U607 ( .A(n1042), .B(n974), .C(n1544), .Y(n1073) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1544) );
  OAI21X1 U609 ( .A(n1043), .B(n974), .C(n1543), .Y(n1072) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1543) );
  OAI21X1 U611 ( .A(n1044), .B(n974), .C(n1542), .Y(n1071) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1542) );
  OAI21X1 U613 ( .A(n1045), .B(n974), .C(n1541), .Y(n1070) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1541) );
  OAI21X1 U615 ( .A(n1046), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1540) );
  OAI21X1 U617 ( .A(n1047), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1539) );
  OAI21X1 U619 ( .A(n1048), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1538) );
  OAI21X1 U621 ( .A(n1049), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1537) );
  NAND3X1 U623 ( .A(n967), .B(n1012), .C(n1655), .Y(n1545) );
  OAI21X1 U624 ( .A(n1034), .B(n8), .C(n1536), .Y(n1065) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1536) );
  OAI21X1 U626 ( .A(n1035), .B(n8), .C(n1535), .Y(n1064) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1535) );
  OAI21X1 U628 ( .A(n1036), .B(n8), .C(n1534), .Y(n1063) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1534) );
  OAI21X1 U630 ( .A(n1037), .B(n8), .C(n1533), .Y(n1062) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1533) );
  OAI21X1 U632 ( .A(n1038), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1532) );
  OAI21X1 U634 ( .A(n1039), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1531) );
  OAI21X1 U636 ( .A(n1040), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1530) );
  OAI21X1 U638 ( .A(n1041), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1529) );
  NOR2X1 U641 ( .A(n964), .B(\addr_1c<4> ), .Y(n1822) );
  OAI21X1 U642 ( .A(n1042), .B(n972), .C(n1526), .Y(n1057) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1526) );
  OAI21X1 U644 ( .A(n1043), .B(n972), .C(n1525), .Y(n1056) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1525) );
  OAI21X1 U646 ( .A(n1044), .B(n972), .C(n1524), .Y(n1055) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1524) );
  OAI21X1 U648 ( .A(n1045), .B(n972), .C(n1523), .Y(n1054) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1523) );
  OAI21X1 U650 ( .A(n1046), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1522) );
  OAI21X1 U652 ( .A(n1047), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1521) );
  OAI21X1 U654 ( .A(n1048), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1520) );
  OAI21X1 U656 ( .A(n1049), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1519) );
  NAND3X1 U658 ( .A(n967), .B(n1013), .C(n1635), .Y(n1527) );
  NOR3X1 U661 ( .A(n1515), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1516) );
  NOR3X1 U662 ( .A(n1514), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1517) );
  AOI21X1 U663 ( .A(n461), .B(n1513), .C(n963), .Y(n1842) );
  OAI21X1 U665 ( .A(rd), .B(n1512), .C(wr), .Y(n1513) );
  NAND3X1 U667 ( .A(n1511), .B(n1029), .C(n1510), .Y(n1512) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1510) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1511) );
  AOI21X1 U670 ( .A(n448), .B(n1508), .C(n1028), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1507), .C(n4), .Y(n1508) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1790), .C(\mem<0><1> ), .D(n1635), .Y(
        n1505) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1810), .C(\mem<2><1> ), .D(n1655), .Y(
        n1506) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1790), .C(\mem<4><1> ), .D(n1635), .Y(
        n1503) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1810), .C(\mem<6><1> ), .D(n1655), .Y(
        n1504) );
  AOI22X1 U678 ( .A(n1595), .B(n892), .C(n1634), .D(n932), .Y(n1509) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1790), .C(\mem<12><1> ), .D(n1635), .Y(
        n1501) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1810), .C(\mem<14><1> ), .D(n1655), .Y(
        n1502) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1790), .C(\mem<8><1> ), .D(n1635), .Y(
        n1499) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1810), .C(\mem<10><1> ), .D(n1655), .Y(
        n1500) );
  AOI21X1 U685 ( .A(n447), .B(n1497), .C(n1028), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1495), .C(n950), .Y(n1497) );
  AOI21X1 U687 ( .A(n1493), .B(n1492), .C(n971), .Y(n1494) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1790), .C(\mem<0><0> ), .D(n1635), .Y(
        n1492) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1810), .C(\mem<2><0> ), .D(n1655), .Y(
        n1493) );
  AOI21X1 U690 ( .A(n1491), .B(n1490), .C(n970), .Y(n1496) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1790), .C(\mem<4><0> ), .D(n1635), .Y(
        n1490) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1810), .C(\mem<6><0> ), .D(n1655), .Y(
        n1491) );
  AOI22X1 U693 ( .A(n1595), .B(n890), .C(n1634), .D(n930), .Y(n1498) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1790), .C(\mem<12><0> ), .D(n1635), .Y(
        n1488) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1810), .C(\mem<14><0> ), .D(n1655), .Y(
        n1489) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1790), .C(\mem<8><0> ), .D(n1635), .Y(
        n1486) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1810), .C(\mem<10><0> ), .D(n1655), .Y(
        n1487) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1485) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1684), .C(\mem<19><7> ), .D(n1703), .Y(
        n1480) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1722), .C(\mem<23><7> ), .D(n1741), .Y(
        n1481) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1760), .C(\mem<27><7> ), .D(n1780), .Y(
        n1483) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1800), .C(\mem<31><7> ), .D(n1821), .Y(
        n1484) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1528), .C(\mem<3><7> ), .D(n1546), .Y(
        n1475) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1566), .C(\mem<7><7> ), .D(n1585), .Y(
        n1476) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1605), .C(\mem<11><7> ), .D(n1624), .Y(
        n1478) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1645), .C(\mem<15><7> ), .D(n1665), .Y(
        n1479) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1474) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1684), .C(\mem<19><6> ), .D(n1703), .Y(
        n1469) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1722), .C(\mem<23><6> ), .D(n1741), .Y(
        n1470) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1760), .C(\mem<27><6> ), .D(n1780), .Y(
        n1472) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1800), .C(\mem<31><6> ), .D(n1821), .Y(
        n1473) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1528), .C(\mem<3><6> ), .D(n1546), .Y(
        n1464) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1566), .C(\mem<7><6> ), .D(n1585), .Y(
        n1465) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1605), .C(\mem<11><6> ), .D(n1624), .Y(
        n1467) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1645), .C(\mem<15><6> ), .D(n1665), .Y(
        n1468) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1463) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1684), .C(\mem<19><5> ), .D(n1703), .Y(
        n1458) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1722), .C(\mem<23><5> ), .D(n1741), .Y(
        n1459) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1760), .C(\mem<27><5> ), .D(n1780), .Y(
        n1461) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1800), .C(\mem<31><5> ), .D(n1821), .Y(
        n1462) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1528), .C(\mem<3><5> ), .D(n1546), .Y(
        n1453) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1566), .C(\mem<7><5> ), .D(n1585), .Y(
        n1454) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1605), .C(\mem<11><5> ), .D(n1624), .Y(
        n1456) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1645), .C(\mem<15><5> ), .D(n1665), .Y(
        n1457) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1452) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1684), .C(\mem<19><4> ), .D(n1703), .Y(
        n1447) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1722), .C(\mem<23><4> ), .D(n1741), .Y(
        n1448) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1760), .C(\mem<27><4> ), .D(n1780), .Y(
        n1450) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1800), .C(\mem<31><4> ), .D(n1821), .Y(
        n1451) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1528), .C(\mem<3><4> ), .D(n1546), .Y(
        n1442) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1566), .C(\mem<7><4> ), .D(n1585), .Y(
        n1443) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1605), .C(\mem<11><4> ), .D(n1624), .Y(
        n1445) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1645), .C(\mem<15><4> ), .D(n1665), .Y(
        n1446) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1441) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1684), .C(\mem<19><3> ), .D(n1703), .Y(
        n1436) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1722), .C(\mem<23><3> ), .D(n1741), .Y(
        n1437) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1760), .C(\mem<27><3> ), .D(n1780), .Y(
        n1439) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1800), .C(\mem<31><3> ), .D(n1821), .Y(
        n1440) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1528), .C(\mem<3><3> ), .D(n1546), .Y(
        n1431) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1566), .C(\mem<7><3> ), .D(n1585), .Y(
        n1432) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1605), .C(\mem<11><3> ), .D(n1624), .Y(
        n1434) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1645), .C(\mem<15><3> ), .D(n1665), .Y(
        n1435) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1430) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1684), .C(\mem<19><2> ), .D(n1703), .Y(
        n1425) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1722), .C(\mem<23><2> ), .D(n1741), .Y(
        n1426) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1760), .C(\mem<27><2> ), .D(n1780), .Y(
        n1428) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1800), .C(\mem<31><2> ), .D(n1821), .Y(
        n1429) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1528), .C(\mem<3><2> ), .D(n1546), .Y(
        n1420) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1566), .C(\mem<7><2> ), .D(n1585), .Y(
        n1421) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1605), .C(\mem<11><2> ), .D(n1624), .Y(
        n1423) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1645), .C(\mem<15><2> ), .D(n1665), .Y(
        n1424) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1419) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1684), .C(\mem<19><1> ), .D(n1703), .Y(
        n1414) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1722), .C(\mem<23><1> ), .D(n1741), .Y(
        n1415) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1760), .C(\mem<27><1> ), .D(n1780), .Y(
        n1417) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1800), .C(\mem<31><1> ), .D(n1821), .Y(
        n1418) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1528), .C(\mem<3><1> ), .D(n1546), .Y(
        n1409) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1566), .C(\mem<7><1> ), .D(n1585), .Y(
        n1410) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1605), .C(\mem<11><1> ), .D(n1624), .Y(
        n1412) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1645), .C(\mem<15><1> ), .D(n1665), .Y(
        n1413) );
  AOI21X1 U777 ( .A(n435), .B(n1407), .C(n1028), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1405), .C(n949), .Y(n1407) );
  AOI21X1 U779 ( .A(n1403), .B(n1402), .C(n971), .Y(n1404) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1790), .C(\mem<0><7> ), .D(n1635), .Y(
        n1402) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1810), .C(\mem<2><7> ), .D(n1655), .Y(
        n1403) );
  AOI21X1 U782 ( .A(n1401), .B(n1400), .C(n970), .Y(n1406) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1790), .C(\mem<4><7> ), .D(n1635), .Y(
        n1400) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1810), .C(\mem<6><7> ), .D(n1655), .Y(
        n1401) );
  AOI22X1 U785 ( .A(n1595), .B(n888), .C(n1634), .D(n928), .Y(n1408) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1790), .C(\mem<12><7> ), .D(n1635), .Y(
        n1398) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1810), .C(\mem<14><7> ), .D(n1655), .Y(
        n1399) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1790), .C(\mem<8><7> ), .D(n1635), .Y(
        n1396) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1810), .C(\mem<10><7> ), .D(n1655), .Y(
        n1397) );
  AOI21X1 U792 ( .A(n434), .B(n1394), .C(n1028), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1392), .C(n948), .Y(n1394) );
  AOI21X1 U794 ( .A(n1390), .B(n1389), .C(n971), .Y(n1391) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1790), .C(\mem<0><6> ), .D(n1635), .Y(
        n1389) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1810), .C(\mem<2><6> ), .D(n1655), .Y(
        n1390) );
  AOI21X1 U797 ( .A(n1388), .B(n1387), .C(n970), .Y(n1393) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1790), .C(\mem<4><6> ), .D(n1635), .Y(
        n1387) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1810), .C(\mem<6><6> ), .D(n1655), .Y(
        n1388) );
  AOI22X1 U800 ( .A(n1595), .B(n886), .C(n1634), .D(n926), .Y(n1395) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1790), .C(\mem<12><6> ), .D(n1635), .Y(
        n1385) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1810), .C(\mem<14><6> ), .D(n1655), .Y(
        n1386) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1790), .C(\mem<8><6> ), .D(n1635), .Y(
        n1383) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1810), .C(\mem<10><6> ), .D(n1655), .Y(
        n1384) );
  AOI21X1 U807 ( .A(n422), .B(n1381), .C(n1028), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1379), .C(n947), .Y(n1381) );
  AOI21X1 U809 ( .A(n1377), .B(n1376), .C(n971), .Y(n1378) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1790), .C(\mem<0><5> ), .D(n1635), .Y(
        n1376) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1810), .C(\mem<2><5> ), .D(n1655), .Y(
        n1377) );
  AOI21X1 U812 ( .A(n1375), .B(n1374), .C(n970), .Y(n1380) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1790), .C(\mem<4><5> ), .D(n1635), .Y(
        n1374) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1810), .C(\mem<6><5> ), .D(n1655), .Y(
        n1375) );
  AOI22X1 U815 ( .A(n1595), .B(n884), .C(n1634), .D(n924), .Y(n1382) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1790), .C(\mem<12><5> ), .D(n1635), .Y(
        n1372) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1810), .C(\mem<14><5> ), .D(n1655), .Y(
        n1373) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1790), .C(\mem<8><5> ), .D(n1635), .Y(
        n1370) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1810), .C(\mem<10><5> ), .D(n1655), .Y(
        n1371) );
  AOI21X1 U822 ( .A(n421), .B(n1368), .C(n1028), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1366), .C(n946), .Y(n1368) );
  AOI21X1 U824 ( .A(n1364), .B(n1363), .C(n971), .Y(n1365) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1790), .C(\mem<0><4> ), .D(n1635), .Y(
        n1363) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1810), .C(\mem<2><4> ), .D(n1655), .Y(
        n1364) );
  AOI21X1 U827 ( .A(n1362), .B(n1361), .C(n970), .Y(n1367) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1790), .C(\mem<4><4> ), .D(n1635), .Y(
        n1361) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1810), .C(\mem<6><4> ), .D(n1655), .Y(
        n1362) );
  AOI22X1 U830 ( .A(n1595), .B(n882), .C(n1634), .D(n922), .Y(n1369) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1790), .C(\mem<12><4> ), .D(n1635), .Y(
        n1359) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1810), .C(\mem<14><4> ), .D(n1655), .Y(
        n1360) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1790), .C(\mem<8><4> ), .D(n1635), .Y(
        n1357) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1810), .C(\mem<10><4> ), .D(n1655), .Y(
        n1358) );
  AOI21X1 U837 ( .A(n409), .B(n1355), .C(n1028), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1353), .C(n945), .Y(n1355) );
  AOI21X1 U839 ( .A(n1351), .B(n1350), .C(n971), .Y(n1352) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1790), .C(\mem<0><3> ), .D(n1635), .Y(
        n1350) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1810), .C(\mem<2><3> ), .D(n1655), .Y(
        n1351) );
  AOI21X1 U842 ( .A(n1349), .B(n1348), .C(n970), .Y(n1354) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1790), .C(\mem<4><3> ), .D(n1635), .Y(
        n1348) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1810), .C(\mem<6><3> ), .D(n1655), .Y(
        n1349) );
  AOI22X1 U845 ( .A(n1595), .B(n880), .C(n1634), .D(n920), .Y(n1356) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1790), .C(\mem<12><3> ), .D(n1635), .Y(
        n1346) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1810), .C(\mem<14><3> ), .D(n1655), .Y(
        n1347) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1790), .C(\mem<8><3> ), .D(n1635), .Y(
        n1344) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1810), .C(\mem<10><3> ), .D(n1655), .Y(
        n1345) );
  AOI21X1 U852 ( .A(n408), .B(n1342), .C(n1028), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1340), .C(n944), .Y(n1342) );
  AOI21X1 U854 ( .A(n1338), .B(n1337), .C(n971), .Y(n1339) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1790), .C(\mem<0><2> ), .D(n1635), .Y(
        n1337) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1810), .C(\mem<2><2> ), .D(n1655), .Y(
        n1338) );
  AOI21X1 U857 ( .A(n1336), .B(n1335), .C(n970), .Y(n1341) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1790), .C(\mem<4><2> ), .D(n1635), .Y(
        n1335) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1810), .C(\mem<6><2> ), .D(n1655), .Y(
        n1336) );
  AOI22X1 U860 ( .A(n1595), .B(n878), .C(n1634), .D(n918), .Y(n1343) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1790), .C(\mem<12><2> ), .D(n1635), .Y(
        n1333) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1810), .C(\mem<14><2> ), .D(n1655), .Y(
        n1334) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1790), .C(\mem<8><2> ), .D(n1635), .Y(
        n1331) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1810), .C(\mem<10><2> ), .D(n1655), .Y(
        n1332) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1330) );
  NOR2X1 U868 ( .A(n1033), .B(\addr_1c<4> ), .Y(n1329) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1328) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1684), .C(\mem<19><0> ), .D(n1703), .Y(
        n1323) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1722), .C(\mem<23><0> ), .D(n1741), .Y(
        n1324) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1760), .C(\mem<27><0> ), .D(n1780), .Y(
        n1326) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1800), .C(\mem<31><0> ), .D(n1821), .Y(
        n1327) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1528), .C(\mem<3><0> ), .D(n1546), .Y(
        n1316) );
  NAND2X1 U877 ( .A(n1031), .B(n1032), .Y(n1518) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1566), .C(\mem<7><0> ), .D(n1585), .Y(
        n1317) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1032), .Y(n1556) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1605), .C(\mem<11><0> ), .D(n1624), .Y(
        n1319) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1645), .C(\mem<15><0> ), .D(n1665), .Y(
        n1320) );
  dff_152 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1016) );
  dff_151 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1016) );
  dff_150 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1016)
         );
  dff_149 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1016)
         );
  dff_148 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1016)
         );
  dff_147 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1016)
         );
  dff_146 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1016)
         );
  dff_145 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1016)
         );
  dff_144 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1016)
         );
  dff_143 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1016)
         );
  dff_142 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1016)
         );
  dff_141 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1016)
         );
  dff_140 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(
        n1016) );
  dff_139 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(
        n1016) );
  dff_138 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(
        n1016) );
  dff_137 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1015) );
  dff_136 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1015) );
  dff_135 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1015) );
  dff_134 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1015) );
  dff_133 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1015) );
  dff_132 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1015) );
  dff_131 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1015) );
  dff_130 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1015) );
  dff_129 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1016) );
  dff_128 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1015) );
  dff_127 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1016) );
  dff_126 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1015) );
  dff_125 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1016) );
  dff_124 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1015) );
  dff_123 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1016) );
  dff_122 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1015) );
  dff_121 \reg2[0]  ( .q(\data_out<0> ), .d(n1025), .clk(clk), .rst(n1016) );
  dff_120 \reg2[1]  ( .q(\data_out<1> ), .d(n1024), .clk(clk), .rst(n1016) );
  dff_119 \reg2[2]  ( .q(\data_out<2> ), .d(n1023), .clk(clk), .rst(n1016) );
  dff_118 \reg2[3]  ( .q(\data_out<3> ), .d(n1022), .clk(clk), .rst(n1016) );
  dff_117 \reg2[4]  ( .q(\data_out<4> ), .d(n1021), .clk(clk), .rst(n1016) );
  dff_116 \reg2[5]  ( .q(\data_out<5> ), .d(n1020), .clk(clk), .rst(n1016) );
  dff_115 \reg2[6]  ( .q(\data_out<6> ), .d(n1019), .clk(clk), .rst(n1016) );
  dff_114 \reg2[7]  ( .q(\data_out<7> ), .d(n1018), .clk(clk), .rst(n1016) );
  dff_113 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), 
        .rst(n1016) );
  dff_112 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), 
        .rst(n1016) );
  dff_111 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1016) );
  dff_110 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1016) );
  dff_109 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1016) );
  dff_108 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1016) );
  dff_107 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1016) );
  dff_106 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1016) );
  dff_105 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1016) );
  dff_104 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1016) );
  dff_103 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1016) );
  dff_102 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1016) );
  INVX1 U2 ( .A(rd), .Y(n1027) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1514) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n1528), .Y(n1831) );
  INVX1 U5 ( .A(rst), .Y(n1017) );
  INVX1 U6 ( .A(n1017), .Y(n1015) );
  INVX1 U7 ( .A(\addr_1c<3> ), .Y(n1033) );
  INVX1 U8 ( .A(\addr_1c<2> ), .Y(n1032) );
  OR2X1 U23 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1515) );
  AND2X1 U24 ( .A(n1634), .B(n965), .Y(n1811) );
  AND2X1 U25 ( .A(n1595), .B(n965), .Y(n1770) );
  INVX1 U26 ( .A(\addr_1c<0> ), .Y(n1030) );
  AND2X1 U27 ( .A(n1030), .B(n1033), .Y(n1314) );
  AND2X1 U28 ( .A(\addr_1c<0> ), .B(n1033), .Y(n1315) );
  AND2X1 U29 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1322) );
  AND2X1 U35 ( .A(\addr_1c<3> ), .B(n1030), .Y(n1321) );
  INVX1 U36 ( .A(\addr_1c<1> ), .Y(n1031) );
  INVX1 U37 ( .A(wr1), .Y(n1029) );
  AND2X1 U38 ( .A(n1595), .B(n1322), .Y(n1780) );
  AND2X1 U39 ( .A(n1595), .B(n1321), .Y(n1760) );
  AND2X1 U40 ( .A(n940), .B(n1322), .Y(n1741) );
  AND2X1 U41 ( .A(n940), .B(n1321), .Y(n1722) );
  AND2X1 U42 ( .A(n1322), .B(n951), .Y(n1703) );
  AND2X1 U43 ( .A(n1321), .B(n951), .Y(n1684) );
  AND2X1 U44 ( .A(n1315), .B(n1595), .Y(n1624) );
  AND2X1 U46 ( .A(n1595), .B(n1314), .Y(n1605) );
  AND2X1 U47 ( .A(n1315), .B(n940), .Y(n1585) );
  AND2X1 U48 ( .A(n940), .B(n1314), .Y(n1566) );
  OR2X1 U49 ( .A(n970), .B(n964), .Y(n968) );
  AND2X1 U50 ( .A(n1315), .B(n951), .Y(n1546) );
  OR2X1 U51 ( .A(n964), .B(n971), .Y(n966) );
  AND2X1 U52 ( .A(n1634), .B(n1314), .Y(n1645) );
  AND2X1 U53 ( .A(n1315), .B(n1634), .Y(n1665) );
  AND2X1 U54 ( .A(n1321), .B(n1634), .Y(n1800) );
  AND2X1 U55 ( .A(\addr_1c<2> ), .B(n1031), .Y(n1595) );
  AND2X1 U56 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1634) );
  BUFX2 U57 ( .A(n961), .Y(n1010) );
  BUFX2 U58 ( .A(n961), .Y(n1009) );
  BUFX2 U59 ( .A(n960), .Y(n1007) );
  BUFX2 U60 ( .A(n960), .Y(n1006) );
  BUFX2 U61 ( .A(n959), .Y(n1004) );
  BUFX2 U62 ( .A(n959), .Y(n1003) );
  BUFX2 U63 ( .A(n958), .Y(n1001) );
  BUFX2 U64 ( .A(n958), .Y(n1000) );
  BUFX2 U65 ( .A(n957), .Y(n990) );
  BUFX2 U66 ( .A(n957), .Y(n989) );
  BUFX2 U67 ( .A(n956), .Y(n987) );
  BUFX2 U68 ( .A(n956), .Y(n986) );
  BUFX2 U69 ( .A(n955), .Y(n984) );
  BUFX2 U70 ( .A(n955), .Y(n983) );
  BUFX2 U71 ( .A(n954), .Y(n981) );
  BUFX2 U72 ( .A(n954), .Y(n980) );
  INVX1 U73 ( .A(\data_in_1c<0> ), .Y(n1034) );
  INVX1 U74 ( .A(\data_in_1c<1> ), .Y(n1035) );
  INVX1 U75 ( .A(\data_in_1c<2> ), .Y(n1036) );
  INVX1 U76 ( .A(\data_in_1c<3> ), .Y(n1037) );
  INVX1 U77 ( .A(\data_in_1c<4> ), .Y(n1038) );
  INVX1 U78 ( .A(\data_in_1c<5> ), .Y(n1039) );
  INVX1 U79 ( .A(\data_in_1c<6> ), .Y(n1040) );
  INVX1 U80 ( .A(\data_in_1c<7> ), .Y(n1041) );
  INVX1 U81 ( .A(\data_in_1c<8> ), .Y(n1042) );
  INVX1 U82 ( .A(\data_in_1c<9> ), .Y(n1043) );
  INVX1 U83 ( .A(\data_in_1c<10> ), .Y(n1044) );
  INVX1 U84 ( .A(\data_in_1c<11> ), .Y(n1045) );
  INVX1 U85 ( .A(\data_in_1c<12> ), .Y(n1046) );
  INVX1 U86 ( .A(\data_in_1c<13> ), .Y(n1047) );
  INVX1 U87 ( .A(\data_in_1c<14> ), .Y(n1048) );
  INVX1 U88 ( .A(\data_in_1c<15> ), .Y(n1049) );
  AND2X1 U89 ( .A(n1831), .B(\mem<32><0> ), .Y(n1495) );
  AND2X1 U90 ( .A(n1831), .B(\mem<32><1> ), .Y(n1507) );
  AND2X1 U91 ( .A(n1831), .B(\mem<32><2> ), .Y(n1340) );
  AND2X1 U92 ( .A(n1831), .B(\mem<32><3> ), .Y(n1353) );
  AND2X1 U93 ( .A(n1831), .B(\mem<32><4> ), .Y(n1366) );
  AND2X1 U129 ( .A(n1831), .B(\mem<32><5> ), .Y(n1379) );
  AND2X1 U589 ( .A(n1831), .B(\mem<32><6> ), .Y(n1392) );
  AND2X1 U640 ( .A(n1831), .B(\mem<32><7> ), .Y(n1405) );
  INVX1 U659 ( .A(rd1), .Y(n1028) );
  INVX1 U660 ( .A(n1017), .Y(n1016) );
  INVX1 U664 ( .A(wr), .Y(n1026) );
  INVX1 U666 ( .A(n1328), .Y(n1025) );
  INVX1 U672 ( .A(n1419), .Y(n1024) );
  INVX1 U675 ( .A(n1430), .Y(n1023) );
  INVX1 U679 ( .A(n1441), .Y(n1022) );
  INVX1 U682 ( .A(n1452), .Y(n1021) );
  INVX1 U694 ( .A(n1463), .Y(n1020) );
  INVX1 U697 ( .A(n1474), .Y(n1019) );
  INVX1 U701 ( .A(n1485), .Y(n1018) );
  INVX1 U706 ( .A(n1832), .Y(n1014) );
  AND2X1 U712 ( .A(wr1), .B(n1017), .Y(n1832) );
  INVX1 U717 ( .A(n1014), .Y(n1012) );
  INVX1 U723 ( .A(n1014), .Y(n1013) );
  AND2X1 U728 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U734 ( .A(n1), .Y(n2) );
  AND2X1 U739 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U745 ( .A(n3), .Y(n4) );
  AND2X1 U750 ( .A(n1821), .B(n189), .Y(n5) );
  INVX1 U756 ( .A(n5), .Y(n6) );
  AND2X1 U761 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U767 ( .A(n7), .Y(n8) );
  OR2X1 U772 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U786 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U789 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U801 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U804 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U816 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U819 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U831 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U834 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U846 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U849 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U861 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U864 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U870 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U875 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U882 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U883 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U884 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U885 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U886 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U887 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U888 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U889 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U890 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U891 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U892 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U893 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U894 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U895 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U896 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U897 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U898 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U899 ( .A(n973), .B(n1832), .Y(n189) );
  AND2X1 U900 ( .A(n1832), .B(n1528), .Y(n289) );
  AND2X1 U901 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U902 ( .A(n348), .Y(n372) );
  AND2X1 U903 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U904 ( .A(n379), .Y(n381) );
  AND2X1 U905 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U906 ( .A(n386), .Y(n387) );
  AND2X1 U907 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U908 ( .A(n401), .Y(n402) );
  BUFX2 U909 ( .A(n1343), .Y(n408) );
  BUFX2 U910 ( .A(n1356), .Y(n409) );
  BUFX2 U911 ( .A(n1369), .Y(n421) );
  BUFX2 U912 ( .A(n1382), .Y(n422) );
  BUFX2 U913 ( .A(n1395), .Y(n434) );
  BUFX2 U914 ( .A(n1408), .Y(n435) );
  BUFX2 U915 ( .A(n1498), .Y(n447) );
  BUFX2 U916 ( .A(n1509), .Y(n448) );
  AND2X2 U917 ( .A(rd), .B(n1512), .Y(n460) );
  INVX1 U918 ( .A(n460), .Y(n461) );
  INVX1 U919 ( .A(n1318), .Y(n473) );
  INVX1 U920 ( .A(n1319), .Y(n474) );
  INVX1 U921 ( .A(n1320), .Y(n486) );
  INVX1 U922 ( .A(n1411), .Y(n487) );
  INVX1 U923 ( .A(n1412), .Y(n507) );
  INVX1 U924 ( .A(n1413), .Y(n508) );
  INVX1 U925 ( .A(n1422), .Y(n522) );
  INVX1 U926 ( .A(n1423), .Y(n523) );
  INVX1 U927 ( .A(n1424), .Y(n537) );
  INVX1 U928 ( .A(n1433), .Y(n538) );
  INVX1 U929 ( .A(n1434), .Y(n552) );
  INVX1 U930 ( .A(n1435), .Y(n553) );
  INVX1 U931 ( .A(n1444), .Y(n567) );
  INVX1 U932 ( .A(n1445), .Y(n568) );
  INVX1 U933 ( .A(n1446), .Y(n582) );
  INVX1 U934 ( .A(n1455), .Y(n583) );
  INVX1 U935 ( .A(n1456), .Y(n591) );
  INVX1 U936 ( .A(n1457), .Y(n592) );
  INVX1 U937 ( .A(n1466), .Y(n871) );
  INVX1 U938 ( .A(n1467), .Y(n872) );
  INVX1 U939 ( .A(n1468), .Y(n873) );
  INVX1 U940 ( .A(n1477), .Y(n874) );
  INVX1 U941 ( .A(n1478), .Y(n875) );
  INVX1 U942 ( .A(n1479), .Y(n876) );
  AND2X2 U943 ( .A(n1332), .B(n1331), .Y(n877) );
  INVX1 U944 ( .A(n877), .Y(n878) );
  AND2X2 U945 ( .A(n1345), .B(n1344), .Y(n879) );
  INVX1 U946 ( .A(n879), .Y(n880) );
  AND2X2 U947 ( .A(n1358), .B(n1357), .Y(n881) );
  INVX1 U948 ( .A(n881), .Y(n882) );
  AND2X2 U949 ( .A(n1371), .B(n1370), .Y(n883) );
  INVX1 U950 ( .A(n883), .Y(n884) );
  AND2X2 U951 ( .A(n1384), .B(n1383), .Y(n885) );
  INVX1 U952 ( .A(n885), .Y(n886) );
  AND2X2 U953 ( .A(n1397), .B(n1396), .Y(n887) );
  INVX1 U954 ( .A(n887), .Y(n888) );
  AND2X2 U955 ( .A(n1487), .B(n1486), .Y(n889) );
  INVX1 U956 ( .A(n889), .Y(n890) );
  AND2X2 U957 ( .A(n1500), .B(n1499), .Y(n891) );
  INVX1 U958 ( .A(n891), .Y(n892) );
  INVX1 U959 ( .A(n1325), .Y(n893) );
  INVX1 U960 ( .A(n1326), .Y(n894) );
  INVX1 U961 ( .A(n1327), .Y(n895) );
  INVX1 U962 ( .A(n1416), .Y(n896) );
  INVX1 U963 ( .A(n1417), .Y(n897) );
  INVX1 U964 ( .A(n1418), .Y(n898) );
  INVX1 U965 ( .A(n1427), .Y(n899) );
  INVX1 U966 ( .A(n1428), .Y(n900) );
  INVX1 U967 ( .A(n1429), .Y(n901) );
  INVX1 U968 ( .A(n1438), .Y(n902) );
  INVX1 U969 ( .A(n1439), .Y(n903) );
  INVX1 U970 ( .A(n1440), .Y(n904) );
  INVX1 U971 ( .A(n1449), .Y(n905) );
  INVX1 U972 ( .A(n1450), .Y(n906) );
  INVX1 U973 ( .A(n1451), .Y(n907) );
  INVX1 U974 ( .A(n1460), .Y(n908) );
  INVX1 U975 ( .A(n1461), .Y(n909) );
  INVX1 U976 ( .A(n1462), .Y(n910) );
  INVX1 U977 ( .A(n1471), .Y(n911) );
  INVX1 U978 ( .A(n1472), .Y(n912) );
  INVX1 U979 ( .A(n1473), .Y(n913) );
  INVX1 U980 ( .A(n1482), .Y(n914) );
  INVX1 U981 ( .A(n1483), .Y(n915) );
  INVX1 U982 ( .A(n1484), .Y(n916) );
  AND2X2 U983 ( .A(n1334), .B(n1333), .Y(n917) );
  INVX1 U984 ( .A(n917), .Y(n918) );
  AND2X2 U985 ( .A(n1347), .B(n1346), .Y(n919) );
  INVX1 U986 ( .A(n919), .Y(n920) );
  AND2X2 U987 ( .A(n1360), .B(n1359), .Y(n921) );
  INVX1 U988 ( .A(n921), .Y(n922) );
  AND2X2 U989 ( .A(n1373), .B(n1372), .Y(n923) );
  INVX1 U990 ( .A(n923), .Y(n924) );
  AND2X2 U991 ( .A(n1386), .B(n1385), .Y(n925) );
  INVX1 U992 ( .A(n925), .Y(n926) );
  AND2X2 U993 ( .A(n1399), .B(n1398), .Y(n927) );
  INVX1 U994 ( .A(n927), .Y(n928) );
  AND2X2 U995 ( .A(n1489), .B(n1488), .Y(n929) );
  INVX1 U996 ( .A(n929), .Y(n930) );
  AND2X2 U997 ( .A(n1502), .B(n1501), .Y(n931) );
  INVX1 U998 ( .A(n931), .Y(n932) );
  BUFX2 U999 ( .A(n1341), .Y(n933) );
  BUFX2 U1000 ( .A(n1354), .Y(n934) );
  BUFX2 U1001 ( .A(n1367), .Y(n935) );
  BUFX2 U1002 ( .A(n1380), .Y(n936) );
  BUFX2 U1003 ( .A(n1393), .Y(n937) );
  BUFX2 U1004 ( .A(n1406), .Y(n938) );
  BUFX2 U1005 ( .A(n1496), .Y(n939) );
  INVX1 U1006 ( .A(n970), .Y(n940) );
  INVX1 U1007 ( .A(n1503), .Y(n941) );
  INVX1 U1008 ( .A(n1504), .Y(n942) );
  BUFX2 U1009 ( .A(n1556), .Y(n970) );
  BUFX2 U1010 ( .A(n1842), .Y(err) );
  BUFX2 U1011 ( .A(n1339), .Y(n944) );
  BUFX2 U1012 ( .A(n1352), .Y(n945) );
  BUFX2 U1013 ( .A(n1365), .Y(n946) );
  BUFX2 U1014 ( .A(n1378), .Y(n947) );
  BUFX2 U1015 ( .A(n1391), .Y(n948) );
  BUFX2 U1016 ( .A(n1404), .Y(n949) );
  BUFX2 U1017 ( .A(n1494), .Y(n950) );
  INVX1 U1018 ( .A(n971), .Y(n951) );
  INVX1 U1019 ( .A(n1505), .Y(n952) );
  INVX1 U1020 ( .A(n1506), .Y(n953) );
  BUFX2 U1021 ( .A(n1518), .Y(n971) );
  BUFX2 U1022 ( .A(n1527), .Y(n972) );
  BUFX2 U1023 ( .A(n1545), .Y(n974) );
  BUFX2 U1024 ( .A(n1555), .Y(n975) );
  BUFX2 U1025 ( .A(n1565), .Y(n976) );
  BUFX2 U1026 ( .A(n1575), .Y(n977) );
  BUFX2 U1027 ( .A(n1584), .Y(n978) );
  BUFX2 U1028 ( .A(n1594), .Y(n979) );
  BUFX2 U1029 ( .A(n1614), .Y(n982) );
  BUFX2 U1030 ( .A(n1633), .Y(n985) );
  BUFX2 U1031 ( .A(n1654), .Y(n988) );
  BUFX2 U1032 ( .A(n1674), .Y(n991) );
  BUFX2 U1033 ( .A(n1683), .Y(n992) );
  BUFX2 U1034 ( .A(n1693), .Y(n993) );
  BUFX2 U1035 ( .A(n1702), .Y(n994) );
  BUFX2 U1036 ( .A(n1712), .Y(n995) );
  BUFX2 U1037 ( .A(n1721), .Y(n996) );
  BUFX2 U1038 ( .A(n1731), .Y(n997) );
  BUFX2 U1039 ( .A(n1740), .Y(n998) );
  BUFX2 U1040 ( .A(n1750), .Y(n999) );
  BUFX2 U1041 ( .A(n1769), .Y(n1002) );
  BUFX2 U1042 ( .A(n1789), .Y(n1005) );
  BUFX2 U1043 ( .A(n1809), .Y(n1008) );
  BUFX2 U1044 ( .A(n1822), .Y(n973) );
  AND2X1 U1045 ( .A(n1634), .B(n1322), .Y(n1821) );
  BUFX2 U1046 ( .A(n1841), .Y(n1011) );
  BUFX2 U1047 ( .A(n1604), .Y(n954) );
  BUFX2 U1048 ( .A(n1623), .Y(n955) );
  BUFX2 U1049 ( .A(n1644), .Y(n956) );
  BUFX2 U1050 ( .A(n1664), .Y(n957) );
  BUFX2 U1051 ( .A(n1759), .Y(n958) );
  BUFX2 U1052 ( .A(n1779), .Y(n959) );
  BUFX2 U1053 ( .A(n1799), .Y(n960) );
  BUFX2 U1054 ( .A(n1820), .Y(n961) );
  AND2X1 U1055 ( .A(enable), .B(n1017), .Y(n962) );
  INVX1 U1056 ( .A(n962), .Y(n963) );
  INVX1 U1057 ( .A(n965), .Y(n964) );
  AND2X1 U1058 ( .A(n1517), .B(n1516), .Y(n965) );
  INVX1 U1059 ( .A(n966), .Y(n967) );
  INVX1 U1060 ( .A(n968), .Y(n969) );
  AND2X1 U1061 ( .A(n951), .B(n1314), .Y(n1528) );
endmodule


module final_memory_1 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1842, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1050), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1051), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1052), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1053), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1054), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1055), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1056), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1057), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1058), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1059), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1060), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1061), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1062), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1063), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1064), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1065), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1066), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1067), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1068), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1069), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1070), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1071), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1072), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1073), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1074), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1075), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1076), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1077), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1078), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1079), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1080), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1081), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1082), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1083), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1084), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1085), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1086), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1087), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1088), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1089), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1090), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1091), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1092), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1093), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1094), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1095), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1096), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1097), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1098), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1099), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1100), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1101), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1102), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1103), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1104), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1105), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1106), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1107), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1108), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1109), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1110), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1111), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1112), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1113), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1114), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1115), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1116), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1117), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1118), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1119), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1120), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1121), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1122), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1123), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1124), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1125), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1126), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1127), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1128), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1129), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1130), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1131), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1132), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1133), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1134), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1135), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1136), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1137), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1138), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1139), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1140), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1141), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1142), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1143), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1144), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1145), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1146), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1147), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1148), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1149), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1150), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1151), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1152), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1153), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1154), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1155), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1156), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1157), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1158), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1159), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1160), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1161), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1162), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1163), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1164), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1165), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1166), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1167), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1168), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1169), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1170), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1171), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1172), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1173), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1174), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1175), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1176), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1177), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1178), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1179), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1180), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1181), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1182), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1183), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1184), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1185), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1186), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1187), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1188), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1189), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1190), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1191), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1192), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1193), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1194), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1195), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1196), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1197), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1198), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1199), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1200), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1201), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1202), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1203), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1204), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1205), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1206), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1207), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1208), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1209), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1210), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1211), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1212), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1213), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1214), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1215), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1216), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1217), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1218), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1219), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1220), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1221), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1222), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1223), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1224), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1225), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1226), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1227), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1228), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1229), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1230), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1231), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1232), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1233), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1234), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1235), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1236), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1237), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1238), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1239), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1240), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1241), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1242), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1243), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1244), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1245), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1246), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1247), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1248), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1249), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1250), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1251), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1252), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1253), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1254), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1255), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1256), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1257), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1258), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1259), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1260), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1261), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1262), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1263), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1264), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1265), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1266), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1267), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1268), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1269), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1270), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1271), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1272), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1273), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1274), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1275), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1276), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1277), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1278), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1279), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1280), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1281), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1282), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1283), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1284), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1285), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1286), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1287), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1288), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1289), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1290), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1291), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1292), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1293), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1294), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1295), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1296), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1297), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1298), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1299), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1300), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1301), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1302), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1303), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1304), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1305), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1306), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1307), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1308), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1309), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1310), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1311), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1312), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1313), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1481), .B(n1480), .Y(n1482) );
  AND2X2 U10 ( .A(n1476), .B(n1475), .Y(n1477) );
  AND2X2 U11 ( .A(n1470), .B(n1469), .Y(n1471) );
  AND2X2 U12 ( .A(n1465), .B(n1464), .Y(n1466) );
  AND2X2 U13 ( .A(n1459), .B(n1458), .Y(n1460) );
  AND2X2 U14 ( .A(n1454), .B(n1453), .Y(n1455) );
  AND2X2 U15 ( .A(n1448), .B(n1447), .Y(n1449) );
  AND2X2 U16 ( .A(n1443), .B(n1442), .Y(n1444) );
  AND2X2 U17 ( .A(n1437), .B(n1436), .Y(n1438) );
  AND2X2 U18 ( .A(n1432), .B(n1431), .Y(n1433) );
  AND2X2 U19 ( .A(n1426), .B(n1425), .Y(n1427) );
  AND2X2 U20 ( .A(n1421), .B(n1420), .Y(n1422) );
  AND2X2 U21 ( .A(n1415), .B(n1414), .Y(n1416) );
  AND2X2 U22 ( .A(n1410), .B(n1409), .Y(n1411) );
  AND2X2 U30 ( .A(n1330), .B(n1030), .Y(n1635) );
  AND2X2 U31 ( .A(n1329), .B(n1030), .Y(n1790) );
  AND2X2 U32 ( .A(n1330), .B(\addr_1c<0> ), .Y(n1655) );
  AND2X2 U33 ( .A(n1329), .B(\addr_1c<0> ), .Y(n1810) );
  AND2X2 U34 ( .A(n1324), .B(n1323), .Y(n1325) );
  AND2X2 U45 ( .A(n1317), .B(n1316), .Y(n1318) );
  NOR3X1 U94 ( .A(n1026), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1027), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1042), .C(n1840), .Y(n1313) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1840) );
  OAI21X1 U98 ( .A(n1011), .B(n1043), .C(n1839), .Y(n1312) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1839) );
  OAI21X1 U100 ( .A(n1011), .B(n1044), .C(n1838), .Y(n1311) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1838) );
  OAI21X1 U102 ( .A(n1011), .B(n1045), .C(n1837), .Y(n1310) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1837) );
  OAI21X1 U104 ( .A(n1011), .B(n1046), .C(n1836), .Y(n1309) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1836) );
  OAI21X1 U106 ( .A(n1011), .B(n1047), .C(n1835), .Y(n1308) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1835) );
  OAI21X1 U108 ( .A(n1011), .B(n1048), .C(n1834), .Y(n1307) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1834) );
  OAI21X1 U110 ( .A(n1011), .B(n1049), .C(n1833), .Y(n1306) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1833) );
  NAND3X1 U112 ( .A(n1012), .B(n1831), .C(n965), .Y(n1841) );
  OAI21X1 U113 ( .A(n6), .B(n1034), .C(n1830), .Y(n1305) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1830) );
  OAI21X1 U115 ( .A(n6), .B(n1035), .C(n1829), .Y(n1304) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1829) );
  OAI21X1 U117 ( .A(n6), .B(n1036), .C(n1828), .Y(n1303) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1828) );
  OAI21X1 U119 ( .A(n6), .B(n1037), .C(n1827), .Y(n1302) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1827) );
  OAI21X1 U121 ( .A(n6), .B(n1038), .C(n1826), .Y(n1301) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1826) );
  OAI21X1 U123 ( .A(n6), .B(n1039), .C(n1825), .Y(n1300) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1825) );
  OAI21X1 U125 ( .A(n6), .B(n1040), .C(n1824), .Y(n1299) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1824) );
  OAI21X1 U127 ( .A(n6), .B(n1041), .C(n1823), .Y(n1298) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1823) );
  OAI21X1 U130 ( .A(n1042), .B(n1010), .C(n1819), .Y(n1297) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1819) );
  OAI21X1 U132 ( .A(n1043), .B(n1009), .C(n1818), .Y(n1296) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1818) );
  OAI21X1 U134 ( .A(n1044), .B(n1009), .C(n1817), .Y(n1295) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1817) );
  OAI21X1 U136 ( .A(n1045), .B(n1009), .C(n1816), .Y(n1294) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1816) );
  OAI21X1 U138 ( .A(n1046), .B(n1009), .C(n1815), .Y(n1293) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1815) );
  OAI21X1 U140 ( .A(n1047), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1814) );
  OAI21X1 U142 ( .A(n1048), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1813) );
  OAI21X1 U144 ( .A(n1049), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1812) );
  NAND3X1 U146 ( .A(n1811), .B(n1832), .C(n1810), .Y(n1820) );
  OAI21X1 U147 ( .A(n1034), .B(n1008), .C(n1808), .Y(n1289) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1808) );
  OAI21X1 U149 ( .A(n1035), .B(n1008), .C(n1807), .Y(n1288) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1807) );
  OAI21X1 U151 ( .A(n1036), .B(n1008), .C(n1806), .Y(n1287) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1806) );
  OAI21X1 U153 ( .A(n1037), .B(n1008), .C(n1805), .Y(n1286) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1805) );
  OAI21X1 U155 ( .A(n1038), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1804) );
  OAI21X1 U157 ( .A(n1039), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1803) );
  OAI21X1 U159 ( .A(n1040), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1802) );
  OAI21X1 U161 ( .A(n1041), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1801) );
  NAND3X1 U163 ( .A(n973), .B(n1013), .C(n1800), .Y(n1809) );
  OAI21X1 U164 ( .A(n1042), .B(n1007), .C(n1798), .Y(n1281) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1798) );
  OAI21X1 U166 ( .A(n1043), .B(n1006), .C(n1797), .Y(n1280) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1797) );
  OAI21X1 U168 ( .A(n1044), .B(n1006), .C(n1796), .Y(n1279) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1796) );
  OAI21X1 U170 ( .A(n1045), .B(n1006), .C(n1795), .Y(n1278) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1795) );
  OAI21X1 U172 ( .A(n1046), .B(n1006), .C(n1794), .Y(n1277) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1794) );
  OAI21X1 U174 ( .A(n1047), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1793) );
  OAI21X1 U176 ( .A(n1048), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1792) );
  OAI21X1 U178 ( .A(n1049), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1791) );
  NAND3X1 U180 ( .A(n1811), .B(n1832), .C(n1790), .Y(n1799) );
  OAI21X1 U181 ( .A(n1034), .B(n1005), .C(n1788), .Y(n1273) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1788) );
  OAI21X1 U183 ( .A(n1035), .B(n1005), .C(n1787), .Y(n1272) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1787) );
  OAI21X1 U185 ( .A(n1036), .B(n1005), .C(n1786), .Y(n1271) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1786) );
  OAI21X1 U187 ( .A(n1037), .B(n1005), .C(n1785), .Y(n1270) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1785) );
  OAI21X1 U189 ( .A(n1038), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1784) );
  OAI21X1 U191 ( .A(n1039), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1783) );
  OAI21X1 U193 ( .A(n1040), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1782) );
  OAI21X1 U195 ( .A(n1041), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1781) );
  NAND3X1 U197 ( .A(n973), .B(n1012), .C(n1780), .Y(n1789) );
  OAI21X1 U198 ( .A(n1042), .B(n1004), .C(n1778), .Y(n1265) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1778) );
  OAI21X1 U200 ( .A(n1043), .B(n1003), .C(n1777), .Y(n1264) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1777) );
  OAI21X1 U202 ( .A(n1044), .B(n1003), .C(n1776), .Y(n1263) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1776) );
  OAI21X1 U204 ( .A(n1045), .B(n1003), .C(n1775), .Y(n1262) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1775) );
  OAI21X1 U206 ( .A(n1046), .B(n1003), .C(n1774), .Y(n1261) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1774) );
  OAI21X1 U208 ( .A(n1047), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1773) );
  OAI21X1 U210 ( .A(n1048), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1772) );
  OAI21X1 U212 ( .A(n1049), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1771) );
  NAND3X1 U214 ( .A(n1810), .B(n1013), .C(n1770), .Y(n1779) );
  OAI21X1 U215 ( .A(n1034), .B(n1002), .C(n1768), .Y(n1257) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1768) );
  OAI21X1 U217 ( .A(n1035), .B(n1002), .C(n1767), .Y(n1256) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1767) );
  OAI21X1 U219 ( .A(n1036), .B(n1002), .C(n1766), .Y(n1255) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1766) );
  OAI21X1 U221 ( .A(n1037), .B(n1002), .C(n1765), .Y(n1254) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1765) );
  OAI21X1 U223 ( .A(n1038), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1764) );
  OAI21X1 U225 ( .A(n1039), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1763) );
  OAI21X1 U227 ( .A(n1040), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1762) );
  OAI21X1 U229 ( .A(n1041), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1761) );
  NAND3X1 U231 ( .A(n973), .B(n1013), .C(n1760), .Y(n1769) );
  OAI21X1 U232 ( .A(n1042), .B(n1001), .C(n1758), .Y(n1249) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1758) );
  OAI21X1 U234 ( .A(n1043), .B(n1000), .C(n1757), .Y(n1248) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1757) );
  OAI21X1 U236 ( .A(n1044), .B(n1000), .C(n1756), .Y(n1247) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1756) );
  OAI21X1 U238 ( .A(n1045), .B(n1000), .C(n1755), .Y(n1246) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1755) );
  OAI21X1 U240 ( .A(n1046), .B(n1000), .C(n1754), .Y(n1245) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1754) );
  OAI21X1 U242 ( .A(n1047), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1753) );
  OAI21X1 U244 ( .A(n1048), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1752) );
  OAI21X1 U246 ( .A(n1049), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1751) );
  NAND3X1 U248 ( .A(n1790), .B(n1013), .C(n1770), .Y(n1759) );
  OAI21X1 U249 ( .A(n1034), .B(n999), .C(n1749), .Y(n1241) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1749) );
  OAI21X1 U251 ( .A(n1035), .B(n999), .C(n1748), .Y(n1240) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1748) );
  OAI21X1 U253 ( .A(n1036), .B(n999), .C(n1747), .Y(n1239) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1747) );
  OAI21X1 U255 ( .A(n1037), .B(n999), .C(n1746), .Y(n1238) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1746) );
  OAI21X1 U257 ( .A(n1038), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1745) );
  OAI21X1 U259 ( .A(n1039), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1744) );
  OAI21X1 U261 ( .A(n1040), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1743) );
  OAI21X1 U263 ( .A(n1041), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1742) );
  NAND3X1 U265 ( .A(n973), .B(n1013), .C(n1741), .Y(n1750) );
  OAI21X1 U266 ( .A(n1042), .B(n998), .C(n1739), .Y(n1233) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1739) );
  OAI21X1 U268 ( .A(n1043), .B(n998), .C(n1738), .Y(n1232) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1738) );
  OAI21X1 U270 ( .A(n1044), .B(n998), .C(n1737), .Y(n1231) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1737) );
  OAI21X1 U272 ( .A(n1045), .B(n998), .C(n1736), .Y(n1230) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1736) );
  OAI21X1 U274 ( .A(n1046), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1735) );
  OAI21X1 U276 ( .A(n1047), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1734) );
  OAI21X1 U278 ( .A(n1048), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1733) );
  OAI21X1 U280 ( .A(n1049), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1732) );
  NAND3X1 U282 ( .A(n1810), .B(n1013), .C(n969), .Y(n1740) );
  OAI21X1 U283 ( .A(n1034), .B(n997), .C(n1730), .Y(n1225) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1730) );
  OAI21X1 U285 ( .A(n1035), .B(n997), .C(n1729), .Y(n1224) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1729) );
  OAI21X1 U287 ( .A(n1036), .B(n997), .C(n1728), .Y(n1223) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1728) );
  OAI21X1 U289 ( .A(n1037), .B(n997), .C(n1727), .Y(n1222) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1727) );
  OAI21X1 U291 ( .A(n1038), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1726) );
  OAI21X1 U293 ( .A(n1039), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1725) );
  OAI21X1 U295 ( .A(n1040), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1724) );
  OAI21X1 U297 ( .A(n1041), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1723) );
  NAND3X1 U299 ( .A(n973), .B(n1013), .C(n1722), .Y(n1731) );
  OAI21X1 U300 ( .A(n1042), .B(n996), .C(n1720), .Y(n1217) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1720) );
  OAI21X1 U302 ( .A(n1043), .B(n996), .C(n1719), .Y(n1216) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1719) );
  OAI21X1 U304 ( .A(n1044), .B(n996), .C(n1718), .Y(n1215) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1718) );
  OAI21X1 U306 ( .A(n1045), .B(n996), .C(n1717), .Y(n1214) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1717) );
  OAI21X1 U308 ( .A(n1046), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1716) );
  OAI21X1 U310 ( .A(n1047), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1715) );
  OAI21X1 U312 ( .A(n1048), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1714) );
  OAI21X1 U314 ( .A(n1049), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1713) );
  NAND3X1 U316 ( .A(n1790), .B(n1013), .C(n969), .Y(n1721) );
  OAI21X1 U317 ( .A(n1034), .B(n995), .C(n1711), .Y(n1209) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1711) );
  OAI21X1 U319 ( .A(n1035), .B(n995), .C(n1710), .Y(n1208) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1710) );
  OAI21X1 U321 ( .A(n1036), .B(n995), .C(n1709), .Y(n1207) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1709) );
  OAI21X1 U323 ( .A(n1037), .B(n995), .C(n1708), .Y(n1206) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1708) );
  OAI21X1 U325 ( .A(n1038), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1707) );
  OAI21X1 U327 ( .A(n1039), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1706) );
  OAI21X1 U329 ( .A(n1040), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1705) );
  OAI21X1 U331 ( .A(n1041), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1704) );
  NAND3X1 U333 ( .A(n973), .B(n1013), .C(n1703), .Y(n1712) );
  OAI21X1 U334 ( .A(n1042), .B(n994), .C(n1701), .Y(n1201) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1701) );
  OAI21X1 U336 ( .A(n1043), .B(n994), .C(n1700), .Y(n1200) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1700) );
  OAI21X1 U338 ( .A(n1044), .B(n994), .C(n1699), .Y(n1199) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1699) );
  OAI21X1 U340 ( .A(n1045), .B(n994), .C(n1698), .Y(n1198) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1698) );
  OAI21X1 U342 ( .A(n1046), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1697) );
  OAI21X1 U344 ( .A(n1047), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1696) );
  OAI21X1 U346 ( .A(n1048), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1695) );
  OAI21X1 U348 ( .A(n1049), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1694) );
  NAND3X1 U350 ( .A(n1810), .B(n1013), .C(n967), .Y(n1702) );
  OAI21X1 U351 ( .A(n1034), .B(n993), .C(n1692), .Y(n1193) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1692) );
  OAI21X1 U353 ( .A(n1035), .B(n993), .C(n1691), .Y(n1192) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1691) );
  OAI21X1 U355 ( .A(n1036), .B(n993), .C(n1690), .Y(n1191) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1690) );
  OAI21X1 U357 ( .A(n1037), .B(n993), .C(n1689), .Y(n1190) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1689) );
  OAI21X1 U359 ( .A(n1038), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1688) );
  OAI21X1 U361 ( .A(n1039), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1687) );
  OAI21X1 U363 ( .A(n1040), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1686) );
  OAI21X1 U365 ( .A(n1041), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1685) );
  NAND3X1 U367 ( .A(n973), .B(n1013), .C(n1684), .Y(n1693) );
  OAI21X1 U368 ( .A(n1042), .B(n992), .C(n1682), .Y(n1185) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1682) );
  OAI21X1 U370 ( .A(n1043), .B(n992), .C(n1681), .Y(n1184) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1681) );
  OAI21X1 U372 ( .A(n1044), .B(n992), .C(n1680), .Y(n1183) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1680) );
  OAI21X1 U374 ( .A(n1045), .B(n992), .C(n1679), .Y(n1182) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1679) );
  OAI21X1 U376 ( .A(n1046), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1678) );
  OAI21X1 U378 ( .A(n1047), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1677) );
  OAI21X1 U380 ( .A(n1048), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1676) );
  OAI21X1 U382 ( .A(n1049), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1675) );
  NAND3X1 U384 ( .A(n1790), .B(n1013), .C(n967), .Y(n1683) );
  OAI21X1 U385 ( .A(n1034), .B(n991), .C(n1673), .Y(n1177) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1673) );
  OAI21X1 U387 ( .A(n1035), .B(n991), .C(n1672), .Y(n1176) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1672) );
  OAI21X1 U389 ( .A(n1036), .B(n991), .C(n1671), .Y(n1175) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1671) );
  OAI21X1 U391 ( .A(n1037), .B(n991), .C(n1670), .Y(n1174) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1670) );
  OAI21X1 U393 ( .A(n1038), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1669) );
  OAI21X1 U395 ( .A(n1039), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1668) );
  OAI21X1 U397 ( .A(n1040), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1667) );
  OAI21X1 U399 ( .A(n1041), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1666) );
  NAND3X1 U401 ( .A(n973), .B(n1013), .C(n1665), .Y(n1674) );
  OAI21X1 U402 ( .A(n1042), .B(n990), .C(n1663), .Y(n1169) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1663) );
  OAI21X1 U404 ( .A(n1043), .B(n989), .C(n1662), .Y(n1168) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1662) );
  OAI21X1 U406 ( .A(n1044), .B(n989), .C(n1661), .Y(n1167) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1661) );
  OAI21X1 U408 ( .A(n1045), .B(n989), .C(n1660), .Y(n1166) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1660) );
  OAI21X1 U410 ( .A(n1046), .B(n989), .C(n1659), .Y(n1165) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1659) );
  OAI21X1 U412 ( .A(n1047), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1658) );
  OAI21X1 U414 ( .A(n1048), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1657) );
  OAI21X1 U416 ( .A(n1049), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1656) );
  NAND3X1 U418 ( .A(n1811), .B(n1012), .C(n1655), .Y(n1664) );
  OAI21X1 U419 ( .A(n1034), .B(n988), .C(n1653), .Y(n1161) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1653) );
  OAI21X1 U421 ( .A(n1035), .B(n988), .C(n1652), .Y(n1160) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1652) );
  OAI21X1 U423 ( .A(n1036), .B(n988), .C(n1651), .Y(n1159) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1651) );
  OAI21X1 U425 ( .A(n1037), .B(n988), .C(n1650), .Y(n1158) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1650) );
  OAI21X1 U427 ( .A(n1038), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1649) );
  OAI21X1 U429 ( .A(n1039), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1648) );
  OAI21X1 U431 ( .A(n1040), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1647) );
  OAI21X1 U433 ( .A(n1041), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1646) );
  NAND3X1 U435 ( .A(n973), .B(n1012), .C(n1645), .Y(n1654) );
  OAI21X1 U436 ( .A(n1042), .B(n987), .C(n1643), .Y(n1153) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1643) );
  OAI21X1 U438 ( .A(n1043), .B(n986), .C(n1642), .Y(n1152) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1642) );
  OAI21X1 U440 ( .A(n1044), .B(n986), .C(n1641), .Y(n1151) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1641) );
  OAI21X1 U442 ( .A(n1045), .B(n986), .C(n1640), .Y(n1150) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1640) );
  OAI21X1 U444 ( .A(n1046), .B(n986), .C(n1639), .Y(n1149) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1639) );
  OAI21X1 U446 ( .A(n1047), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1638) );
  OAI21X1 U448 ( .A(n1048), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1637) );
  OAI21X1 U450 ( .A(n1049), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1636) );
  NAND3X1 U452 ( .A(n1811), .B(n1012), .C(n1635), .Y(n1644) );
  OAI21X1 U453 ( .A(n1034), .B(n985), .C(n1632), .Y(n1145) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1632) );
  OAI21X1 U455 ( .A(n1035), .B(n985), .C(n1631), .Y(n1144) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1631) );
  OAI21X1 U457 ( .A(n1036), .B(n985), .C(n1630), .Y(n1143) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1630) );
  OAI21X1 U459 ( .A(n1037), .B(n985), .C(n1629), .Y(n1142) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1629) );
  OAI21X1 U461 ( .A(n1038), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1628) );
  OAI21X1 U463 ( .A(n1039), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1627) );
  OAI21X1 U465 ( .A(n1040), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1626) );
  OAI21X1 U467 ( .A(n1041), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1625) );
  NAND3X1 U469 ( .A(n973), .B(n1012), .C(n1624), .Y(n1633) );
  OAI21X1 U470 ( .A(n1042), .B(n984), .C(n1622), .Y(n1137) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1622) );
  OAI21X1 U472 ( .A(n1043), .B(n983), .C(n1621), .Y(n1136) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1621) );
  OAI21X1 U474 ( .A(n1044), .B(n983), .C(n1620), .Y(n1135) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1620) );
  OAI21X1 U476 ( .A(n1045), .B(n983), .C(n1619), .Y(n1134) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1619) );
  OAI21X1 U478 ( .A(n1046), .B(n983), .C(n1618), .Y(n1133) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1618) );
  OAI21X1 U480 ( .A(n1047), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1617) );
  OAI21X1 U482 ( .A(n1048), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1616) );
  OAI21X1 U484 ( .A(n1049), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1615) );
  NAND3X1 U486 ( .A(n1770), .B(n1012), .C(n1655), .Y(n1623) );
  OAI21X1 U487 ( .A(n1034), .B(n982), .C(n1613), .Y(n1129) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1613) );
  OAI21X1 U489 ( .A(n1035), .B(n982), .C(n1612), .Y(n1128) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1612) );
  OAI21X1 U491 ( .A(n1036), .B(n982), .C(n1611), .Y(n1127) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1611) );
  OAI21X1 U493 ( .A(n1037), .B(n982), .C(n1610), .Y(n1126) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1610) );
  OAI21X1 U495 ( .A(n1038), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1609) );
  OAI21X1 U497 ( .A(n1039), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1608) );
  OAI21X1 U499 ( .A(n1040), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1607) );
  OAI21X1 U501 ( .A(n1041), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1606) );
  NAND3X1 U503 ( .A(n973), .B(n1012), .C(n1605), .Y(n1614) );
  OAI21X1 U504 ( .A(n1042), .B(n981), .C(n1603), .Y(n1121) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1603) );
  OAI21X1 U506 ( .A(n1043), .B(n980), .C(n1602), .Y(n1120) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1602) );
  OAI21X1 U508 ( .A(n1044), .B(n980), .C(n1601), .Y(n1119) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1601) );
  OAI21X1 U510 ( .A(n1045), .B(n980), .C(n1600), .Y(n1118) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1600) );
  OAI21X1 U512 ( .A(n1046), .B(n980), .C(n1599), .Y(n1117) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1599) );
  OAI21X1 U514 ( .A(n1047), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1598) );
  OAI21X1 U516 ( .A(n1048), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1597) );
  OAI21X1 U518 ( .A(n1049), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1596) );
  NAND3X1 U520 ( .A(n1770), .B(n1012), .C(n1635), .Y(n1604) );
  OAI21X1 U521 ( .A(n1034), .B(n979), .C(n1593), .Y(n1113) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1593) );
  OAI21X1 U523 ( .A(n1035), .B(n979), .C(n1592), .Y(n1112) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1592) );
  OAI21X1 U525 ( .A(n1036), .B(n979), .C(n1591), .Y(n1111) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1591) );
  OAI21X1 U527 ( .A(n1037), .B(n979), .C(n1590), .Y(n1110) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1590) );
  OAI21X1 U529 ( .A(n1038), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1589) );
  OAI21X1 U531 ( .A(n1039), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1588) );
  OAI21X1 U533 ( .A(n1040), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1587) );
  OAI21X1 U535 ( .A(n1041), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1586) );
  NAND3X1 U537 ( .A(n973), .B(n1012), .C(n1585), .Y(n1594) );
  OAI21X1 U538 ( .A(n1042), .B(n978), .C(n1583), .Y(n1105) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1583) );
  OAI21X1 U540 ( .A(n1043), .B(n978), .C(n1582), .Y(n1104) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1582) );
  OAI21X1 U542 ( .A(n1044), .B(n978), .C(n1581), .Y(n1103) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1581) );
  OAI21X1 U544 ( .A(n1045), .B(n978), .C(n1580), .Y(n1102) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1580) );
  OAI21X1 U546 ( .A(n1046), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1579) );
  OAI21X1 U548 ( .A(n1047), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1578) );
  OAI21X1 U550 ( .A(n1048), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1577) );
  OAI21X1 U552 ( .A(n1049), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1576) );
  NAND3X1 U554 ( .A(n969), .B(n1012), .C(n1655), .Y(n1584) );
  OAI21X1 U555 ( .A(n1034), .B(n977), .C(n1574), .Y(n1097) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1574) );
  OAI21X1 U557 ( .A(n1035), .B(n977), .C(n1573), .Y(n1096) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1573) );
  OAI21X1 U559 ( .A(n1036), .B(n977), .C(n1572), .Y(n1095) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1572) );
  OAI21X1 U561 ( .A(n1037), .B(n977), .C(n1571), .Y(n1094) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1571) );
  OAI21X1 U563 ( .A(n1038), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1570) );
  OAI21X1 U565 ( .A(n1039), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1569) );
  OAI21X1 U567 ( .A(n1040), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1568) );
  OAI21X1 U569 ( .A(n1041), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1567) );
  NAND3X1 U571 ( .A(n973), .B(n1012), .C(n1566), .Y(n1575) );
  OAI21X1 U572 ( .A(n1042), .B(n976), .C(n1564), .Y(n1089) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1564) );
  OAI21X1 U574 ( .A(n1043), .B(n976), .C(n1563), .Y(n1088) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1563) );
  OAI21X1 U576 ( .A(n1044), .B(n976), .C(n1562), .Y(n1087) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1562) );
  OAI21X1 U578 ( .A(n1045), .B(n976), .C(n1561), .Y(n1086) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1561) );
  OAI21X1 U580 ( .A(n1046), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1560) );
  OAI21X1 U582 ( .A(n1047), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1559) );
  OAI21X1 U584 ( .A(n1048), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1558) );
  OAI21X1 U586 ( .A(n1049), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1557) );
  NAND3X1 U588 ( .A(n969), .B(n1012), .C(n1635), .Y(n1565) );
  OAI21X1 U590 ( .A(n1034), .B(n975), .C(n1554), .Y(n1081) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1554) );
  OAI21X1 U592 ( .A(n1035), .B(n975), .C(n1553), .Y(n1080) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1553) );
  OAI21X1 U594 ( .A(n1036), .B(n975), .C(n1552), .Y(n1079) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1552) );
  OAI21X1 U596 ( .A(n1037), .B(n975), .C(n1551), .Y(n1078) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1551) );
  OAI21X1 U598 ( .A(n1038), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1550) );
  OAI21X1 U600 ( .A(n1039), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1549) );
  OAI21X1 U602 ( .A(n1040), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1548) );
  OAI21X1 U604 ( .A(n1041), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1547) );
  NAND3X1 U606 ( .A(n973), .B(n1012), .C(n1546), .Y(n1555) );
  OAI21X1 U607 ( .A(n1042), .B(n974), .C(n1544), .Y(n1073) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1544) );
  OAI21X1 U609 ( .A(n1043), .B(n974), .C(n1543), .Y(n1072) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1543) );
  OAI21X1 U611 ( .A(n1044), .B(n974), .C(n1542), .Y(n1071) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1542) );
  OAI21X1 U613 ( .A(n1045), .B(n974), .C(n1541), .Y(n1070) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1541) );
  OAI21X1 U615 ( .A(n1046), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1540) );
  OAI21X1 U617 ( .A(n1047), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1539) );
  OAI21X1 U619 ( .A(n1048), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1538) );
  OAI21X1 U621 ( .A(n1049), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1537) );
  NAND3X1 U623 ( .A(n967), .B(n1012), .C(n1655), .Y(n1545) );
  OAI21X1 U624 ( .A(n1034), .B(n8), .C(n1536), .Y(n1065) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1536) );
  OAI21X1 U626 ( .A(n1035), .B(n8), .C(n1535), .Y(n1064) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1535) );
  OAI21X1 U628 ( .A(n1036), .B(n8), .C(n1534), .Y(n1063) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1534) );
  OAI21X1 U630 ( .A(n1037), .B(n8), .C(n1533), .Y(n1062) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1533) );
  OAI21X1 U632 ( .A(n1038), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1532) );
  OAI21X1 U634 ( .A(n1039), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1531) );
  OAI21X1 U636 ( .A(n1040), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1530) );
  OAI21X1 U638 ( .A(n1041), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1529) );
  NOR2X1 U641 ( .A(n964), .B(\addr_1c<4> ), .Y(n1822) );
  OAI21X1 U642 ( .A(n1042), .B(n972), .C(n1526), .Y(n1057) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1526) );
  OAI21X1 U644 ( .A(n1043), .B(n972), .C(n1525), .Y(n1056) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1525) );
  OAI21X1 U646 ( .A(n1044), .B(n972), .C(n1524), .Y(n1055) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1524) );
  OAI21X1 U648 ( .A(n1045), .B(n972), .C(n1523), .Y(n1054) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1523) );
  OAI21X1 U650 ( .A(n1046), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1522) );
  OAI21X1 U652 ( .A(n1047), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1521) );
  OAI21X1 U654 ( .A(n1048), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1520) );
  OAI21X1 U656 ( .A(n1049), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1519) );
  NAND3X1 U658 ( .A(n967), .B(n1013), .C(n1635), .Y(n1527) );
  NOR3X1 U661 ( .A(n1515), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1516) );
  NOR3X1 U662 ( .A(n1514), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1517) );
  AOI21X1 U663 ( .A(n461), .B(n1513), .C(n963), .Y(n1842) );
  OAI21X1 U665 ( .A(rd), .B(n1512), .C(wr), .Y(n1513) );
  NAND3X1 U667 ( .A(n1511), .B(n1029), .C(n1510), .Y(n1512) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1510) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1511) );
  AOI21X1 U670 ( .A(n448), .B(n1508), .C(n1028), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1507), .C(n4), .Y(n1508) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1790), .C(\mem<0><1> ), .D(n1635), .Y(
        n1505) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1810), .C(\mem<2><1> ), .D(n1655), .Y(
        n1506) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1790), .C(\mem<4><1> ), .D(n1635), .Y(
        n1503) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1810), .C(\mem<6><1> ), .D(n1655), .Y(
        n1504) );
  AOI22X1 U678 ( .A(n1595), .B(n892), .C(n1634), .D(n932), .Y(n1509) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1790), .C(\mem<12><1> ), .D(n1635), .Y(
        n1501) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1810), .C(\mem<14><1> ), .D(n1655), .Y(
        n1502) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1790), .C(\mem<8><1> ), .D(n1635), .Y(
        n1499) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1810), .C(\mem<10><1> ), .D(n1655), .Y(
        n1500) );
  AOI21X1 U685 ( .A(n447), .B(n1497), .C(n1028), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1495), .C(n949), .Y(n1497) );
  AOI21X1 U687 ( .A(n1493), .B(n1492), .C(n971), .Y(n1494) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1790), .C(\mem<0><0> ), .D(n1635), .Y(
        n1492) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1810), .C(\mem<2><0> ), .D(n1655), .Y(
        n1493) );
  AOI21X1 U690 ( .A(n1491), .B(n1490), .C(n970), .Y(n1496) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1790), .C(\mem<4><0> ), .D(n1635), .Y(
        n1490) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1810), .C(\mem<6><0> ), .D(n1655), .Y(
        n1491) );
  AOI22X1 U693 ( .A(n1595), .B(n890), .C(n1634), .D(n930), .Y(n1498) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1790), .C(\mem<12><0> ), .D(n1635), .Y(
        n1488) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1810), .C(\mem<14><0> ), .D(n1655), .Y(
        n1489) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1790), .C(\mem<8><0> ), .D(n1635), .Y(
        n1486) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1810), .C(\mem<10><0> ), .D(n1655), .Y(
        n1487) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1485) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1684), .C(\mem<19><7> ), .D(n1703), .Y(
        n1480) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1722), .C(\mem<23><7> ), .D(n1741), .Y(
        n1481) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1760), .C(\mem<27><7> ), .D(n1780), .Y(
        n1483) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1800), .C(\mem<31><7> ), .D(n1821), .Y(
        n1484) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1528), .C(\mem<3><7> ), .D(n1546), .Y(
        n1475) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1566), .C(\mem<7><7> ), .D(n1585), .Y(
        n1476) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1605), .C(\mem<11><7> ), .D(n1624), .Y(
        n1478) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1645), .C(\mem<15><7> ), .D(n1665), .Y(
        n1479) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1474) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1684), .C(\mem<19><6> ), .D(n1703), .Y(
        n1469) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1722), .C(\mem<23><6> ), .D(n1741), .Y(
        n1470) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1760), .C(\mem<27><6> ), .D(n1780), .Y(
        n1472) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1800), .C(\mem<31><6> ), .D(n1821), .Y(
        n1473) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1528), .C(\mem<3><6> ), .D(n1546), .Y(
        n1464) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1566), .C(\mem<7><6> ), .D(n1585), .Y(
        n1465) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1605), .C(\mem<11><6> ), .D(n1624), .Y(
        n1467) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1645), .C(\mem<15><6> ), .D(n1665), .Y(
        n1468) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1463) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1684), .C(\mem<19><5> ), .D(n1703), .Y(
        n1458) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1722), .C(\mem<23><5> ), .D(n1741), .Y(
        n1459) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1760), .C(\mem<27><5> ), .D(n1780), .Y(
        n1461) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1800), .C(\mem<31><5> ), .D(n1821), .Y(
        n1462) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1528), .C(\mem<3><5> ), .D(n1546), .Y(
        n1453) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1566), .C(\mem<7><5> ), .D(n1585), .Y(
        n1454) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1605), .C(\mem<11><5> ), .D(n1624), .Y(
        n1456) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1645), .C(\mem<15><5> ), .D(n1665), .Y(
        n1457) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1452) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1684), .C(\mem<19><4> ), .D(n1703), .Y(
        n1447) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1722), .C(\mem<23><4> ), .D(n1741), .Y(
        n1448) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1760), .C(\mem<27><4> ), .D(n1780), .Y(
        n1450) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1800), .C(\mem<31><4> ), .D(n1821), .Y(
        n1451) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1528), .C(\mem<3><4> ), .D(n1546), .Y(
        n1442) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1566), .C(\mem<7><4> ), .D(n1585), .Y(
        n1443) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1605), .C(\mem<11><4> ), .D(n1624), .Y(
        n1445) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1645), .C(\mem<15><4> ), .D(n1665), .Y(
        n1446) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1441) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1684), .C(\mem<19><3> ), .D(n1703), .Y(
        n1436) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1722), .C(\mem<23><3> ), .D(n1741), .Y(
        n1437) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1760), .C(\mem<27><3> ), .D(n1780), .Y(
        n1439) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1800), .C(\mem<31><3> ), .D(n1821), .Y(
        n1440) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1528), .C(\mem<3><3> ), .D(n1546), .Y(
        n1431) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1566), .C(\mem<7><3> ), .D(n1585), .Y(
        n1432) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1605), .C(\mem<11><3> ), .D(n1624), .Y(
        n1434) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1645), .C(\mem<15><3> ), .D(n1665), .Y(
        n1435) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1430) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1684), .C(\mem<19><2> ), .D(n1703), .Y(
        n1425) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1722), .C(\mem<23><2> ), .D(n1741), .Y(
        n1426) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1760), .C(\mem<27><2> ), .D(n1780), .Y(
        n1428) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1800), .C(\mem<31><2> ), .D(n1821), .Y(
        n1429) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1528), .C(\mem<3><2> ), .D(n1546), .Y(
        n1420) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1566), .C(\mem<7><2> ), .D(n1585), .Y(
        n1421) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1605), .C(\mem<11><2> ), .D(n1624), .Y(
        n1423) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1645), .C(\mem<15><2> ), .D(n1665), .Y(
        n1424) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1419) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1684), .C(\mem<19><1> ), .D(n1703), .Y(
        n1414) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1722), .C(\mem<23><1> ), .D(n1741), .Y(
        n1415) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1760), .C(\mem<27><1> ), .D(n1780), .Y(
        n1417) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1800), .C(\mem<31><1> ), .D(n1821), .Y(
        n1418) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1528), .C(\mem<3><1> ), .D(n1546), .Y(
        n1409) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1566), .C(\mem<7><1> ), .D(n1585), .Y(
        n1410) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1605), .C(\mem<11><1> ), .D(n1624), .Y(
        n1412) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1645), .C(\mem<15><1> ), .D(n1665), .Y(
        n1413) );
  AOI21X1 U777 ( .A(n435), .B(n1407), .C(n1028), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1405), .C(n948), .Y(n1407) );
  AOI21X1 U779 ( .A(n1403), .B(n1402), .C(n971), .Y(n1404) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1790), .C(\mem<0><7> ), .D(n1635), .Y(
        n1402) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1810), .C(\mem<2><7> ), .D(n1655), .Y(
        n1403) );
  AOI21X1 U782 ( .A(n1401), .B(n1400), .C(n970), .Y(n1406) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1790), .C(\mem<4><7> ), .D(n1635), .Y(
        n1400) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1810), .C(\mem<6><7> ), .D(n1655), .Y(
        n1401) );
  AOI22X1 U785 ( .A(n1595), .B(n888), .C(n1634), .D(n928), .Y(n1408) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1790), .C(\mem<12><7> ), .D(n1635), .Y(
        n1398) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1810), .C(\mem<14><7> ), .D(n1655), .Y(
        n1399) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1790), .C(\mem<8><7> ), .D(n1635), .Y(
        n1396) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1810), .C(\mem<10><7> ), .D(n1655), .Y(
        n1397) );
  AOI21X1 U792 ( .A(n434), .B(n1394), .C(n1028), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1392), .C(n947), .Y(n1394) );
  AOI21X1 U794 ( .A(n1390), .B(n1389), .C(n971), .Y(n1391) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1790), .C(\mem<0><6> ), .D(n1635), .Y(
        n1389) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1810), .C(\mem<2><6> ), .D(n1655), .Y(
        n1390) );
  AOI21X1 U797 ( .A(n1388), .B(n1387), .C(n970), .Y(n1393) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1790), .C(\mem<4><6> ), .D(n1635), .Y(
        n1387) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1810), .C(\mem<6><6> ), .D(n1655), .Y(
        n1388) );
  AOI22X1 U800 ( .A(n1595), .B(n886), .C(n1634), .D(n926), .Y(n1395) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1790), .C(\mem<12><6> ), .D(n1635), .Y(
        n1385) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1810), .C(\mem<14><6> ), .D(n1655), .Y(
        n1386) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1790), .C(\mem<8><6> ), .D(n1635), .Y(
        n1383) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1810), .C(\mem<10><6> ), .D(n1655), .Y(
        n1384) );
  AOI21X1 U807 ( .A(n422), .B(n1381), .C(n1028), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1379), .C(n946), .Y(n1381) );
  AOI21X1 U809 ( .A(n1377), .B(n1376), .C(n971), .Y(n1378) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1790), .C(\mem<0><5> ), .D(n1635), .Y(
        n1376) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1810), .C(\mem<2><5> ), .D(n1655), .Y(
        n1377) );
  AOI21X1 U812 ( .A(n1375), .B(n1374), .C(n970), .Y(n1380) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1790), .C(\mem<4><5> ), .D(n1635), .Y(
        n1374) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1810), .C(\mem<6><5> ), .D(n1655), .Y(
        n1375) );
  AOI22X1 U815 ( .A(n1595), .B(n884), .C(n1634), .D(n924), .Y(n1382) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1790), .C(\mem<12><5> ), .D(n1635), .Y(
        n1372) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1810), .C(\mem<14><5> ), .D(n1655), .Y(
        n1373) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1790), .C(\mem<8><5> ), .D(n1635), .Y(
        n1370) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1810), .C(\mem<10><5> ), .D(n1655), .Y(
        n1371) );
  AOI21X1 U822 ( .A(n421), .B(n1368), .C(n1028), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1366), .C(n945), .Y(n1368) );
  AOI21X1 U824 ( .A(n1364), .B(n1363), .C(n971), .Y(n1365) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1790), .C(\mem<0><4> ), .D(n1635), .Y(
        n1363) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1810), .C(\mem<2><4> ), .D(n1655), .Y(
        n1364) );
  AOI21X1 U827 ( .A(n1362), .B(n1361), .C(n970), .Y(n1367) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1790), .C(\mem<4><4> ), .D(n1635), .Y(
        n1361) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1810), .C(\mem<6><4> ), .D(n1655), .Y(
        n1362) );
  AOI22X1 U830 ( .A(n1595), .B(n882), .C(n1634), .D(n922), .Y(n1369) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1790), .C(\mem<12><4> ), .D(n1635), .Y(
        n1359) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1810), .C(\mem<14><4> ), .D(n1655), .Y(
        n1360) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1790), .C(\mem<8><4> ), .D(n1635), .Y(
        n1357) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1810), .C(\mem<10><4> ), .D(n1655), .Y(
        n1358) );
  AOI21X1 U837 ( .A(n409), .B(n1355), .C(n1028), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1353), .C(n944), .Y(n1355) );
  AOI21X1 U839 ( .A(n1351), .B(n1350), .C(n971), .Y(n1352) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1790), .C(\mem<0><3> ), .D(n1635), .Y(
        n1350) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1810), .C(\mem<2><3> ), .D(n1655), .Y(
        n1351) );
  AOI21X1 U842 ( .A(n1349), .B(n1348), .C(n970), .Y(n1354) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1790), .C(\mem<4><3> ), .D(n1635), .Y(
        n1348) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1810), .C(\mem<6><3> ), .D(n1655), .Y(
        n1349) );
  AOI22X1 U845 ( .A(n1595), .B(n880), .C(n1634), .D(n920), .Y(n1356) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1790), .C(\mem<12><3> ), .D(n1635), .Y(
        n1346) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1810), .C(\mem<14><3> ), .D(n1655), .Y(
        n1347) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1790), .C(\mem<8><3> ), .D(n1635), .Y(
        n1344) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1810), .C(\mem<10><3> ), .D(n1655), .Y(
        n1345) );
  AOI21X1 U852 ( .A(n408), .B(n1342), .C(n1028), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1340), .C(n943), .Y(n1342) );
  AOI21X1 U854 ( .A(n1338), .B(n1337), .C(n971), .Y(n1339) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1790), .C(\mem<0><2> ), .D(n1635), .Y(
        n1337) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1810), .C(\mem<2><2> ), .D(n1655), .Y(
        n1338) );
  AOI21X1 U857 ( .A(n1336), .B(n1335), .C(n970), .Y(n1341) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1790), .C(\mem<4><2> ), .D(n1635), .Y(
        n1335) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1810), .C(\mem<6><2> ), .D(n1655), .Y(
        n1336) );
  AOI22X1 U860 ( .A(n1595), .B(n878), .C(n1634), .D(n918), .Y(n1343) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1790), .C(\mem<12><2> ), .D(n1635), .Y(
        n1333) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1810), .C(\mem<14><2> ), .D(n1655), .Y(
        n1334) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1790), .C(\mem<8><2> ), .D(n1635), .Y(
        n1331) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1810), .C(\mem<10><2> ), .D(n1655), .Y(
        n1332) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1330) );
  NOR2X1 U868 ( .A(n1033), .B(\addr_1c<4> ), .Y(n1329) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1328) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1684), .C(\mem<19><0> ), .D(n1703), .Y(
        n1323) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1722), .C(\mem<23><0> ), .D(n1741), .Y(
        n1324) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1760), .C(\mem<27><0> ), .D(n1780), .Y(
        n1326) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1800), .C(\mem<31><0> ), .D(n1821), .Y(
        n1327) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1528), .C(\mem<3><0> ), .D(n1546), .Y(
        n1316) );
  NAND2X1 U877 ( .A(n1031), .B(n1032), .Y(n1518) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1566), .C(\mem<7><0> ), .D(n1585), .Y(
        n1317) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1032), .Y(n1556) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1605), .C(\mem<11><0> ), .D(n1624), .Y(
        n1319) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1645), .C(\mem<15><0> ), .D(n1665), .Y(
        n1320) );
  dff_101 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(n1016) );
  dff_100 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(n1016) );
  dff_99 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(n1016)
         );
  dff_98 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(n1016)
         );
  dff_97 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(n1016)
         );
  dff_96 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(n1016)
         );
  dff_95 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(n1016)
         );
  dff_94 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(n1016)
         );
  dff_93 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(n1016)
         );
  dff_92 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(n1016)
         );
  dff_91 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(n1016)
         );
  dff_90 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(n1016)
         );
  dff_89 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(n1016) );
  dff_88 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(n1016) );
  dff_87 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(n1016) );
  dff_86 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        n1015) );
  dff_85 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        n1015) );
  dff_84 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        n1015) );
  dff_83 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        n1015) );
  dff_82 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        n1015) );
  dff_81 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        n1015) );
  dff_80 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        n1015) );
  dff_79 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        n1015) );
  dff_78 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        n1016) );
  dff_77 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        n1015) );
  dff_76 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(n1016) );
  dff_75 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(n1015) );
  dff_74 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(n1016) );
  dff_73 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(n1015) );
  dff_72 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(n1016) );
  dff_71 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(n1015) );
  dff_70 \reg2[0]  ( .q(\data_out<0> ), .d(n1025), .clk(clk), .rst(n1016) );
  dff_69 \reg2[1]  ( .q(\data_out<1> ), .d(n1024), .clk(clk), .rst(n1016) );
  dff_68 \reg2[2]  ( .q(\data_out<2> ), .d(n1023), .clk(clk), .rst(n1016) );
  dff_67 \reg2[3]  ( .q(\data_out<3> ), .d(n1022), .clk(clk), .rst(n1016) );
  dff_66 \reg2[4]  ( .q(\data_out<4> ), .d(n1021), .clk(clk), .rst(n1016) );
  dff_65 \reg2[5]  ( .q(\data_out<5> ), .d(n1020), .clk(clk), .rst(n1016) );
  dff_64 \reg2[6]  ( .q(\data_out<6> ), .d(n1019), .clk(clk), .rst(n1016) );
  dff_63 \reg2[7]  ( .q(\data_out<7> ), .d(n1018), .clk(clk), .rst(n1016) );
  dff_62 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        n1016) );
  dff_61 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        n1016) );
  dff_60 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(n1016) );
  dff_59 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(n1016) );
  dff_58 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(n1016) );
  dff_57 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(n1016) );
  dff_56 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(n1016) );
  dff_55 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(n1016) );
  dff_54 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(n1016) );
  dff_53 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(n1016) );
  dff_52 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(n1016) );
  dff_51 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(n1016) );
  INVX1 U2 ( .A(rd), .Y(n1027) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1514) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n1528), .Y(n1831) );
  INVX1 U5 ( .A(rst), .Y(n1017) );
  INVX1 U6 ( .A(n1017), .Y(n1015) );
  INVX1 U7 ( .A(\addr_1c<3> ), .Y(n1033) );
  INVX1 U8 ( .A(\addr_1c<2> ), .Y(n1032) );
  OR2X1 U23 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1515) );
  AND2X1 U24 ( .A(n1634), .B(n965), .Y(n1811) );
  AND2X1 U25 ( .A(n1595), .B(n965), .Y(n1770) );
  INVX1 U26 ( .A(\addr_1c<0> ), .Y(n1030) );
  AND2X1 U27 ( .A(n1030), .B(n1033), .Y(n1314) );
  AND2X1 U28 ( .A(\addr_1c<0> ), .B(n1033), .Y(n1315) );
  AND2X1 U29 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1322) );
  AND2X1 U35 ( .A(\addr_1c<3> ), .B(n1030), .Y(n1321) );
  INVX1 U36 ( .A(\addr_1c<1> ), .Y(n1031) );
  INVX1 U37 ( .A(wr1), .Y(n1029) );
  AND2X1 U38 ( .A(n1595), .B(n1322), .Y(n1780) );
  AND2X1 U39 ( .A(n1595), .B(n1321), .Y(n1760) );
  AND2X1 U40 ( .A(n940), .B(n1322), .Y(n1741) );
  AND2X1 U41 ( .A(n940), .B(n1321), .Y(n1722) );
  AND2X1 U42 ( .A(n1322), .B(n950), .Y(n1703) );
  AND2X1 U43 ( .A(n1321), .B(n950), .Y(n1684) );
  AND2X1 U44 ( .A(n1315), .B(n1595), .Y(n1624) );
  AND2X1 U46 ( .A(n1595), .B(n1314), .Y(n1605) );
  AND2X1 U47 ( .A(n1315), .B(n940), .Y(n1585) );
  AND2X1 U48 ( .A(n940), .B(n1314), .Y(n1566) );
  OR2X1 U49 ( .A(n970), .B(n964), .Y(n968) );
  AND2X1 U50 ( .A(n1315), .B(n950), .Y(n1546) );
  OR2X1 U51 ( .A(n964), .B(n971), .Y(n966) );
  AND2X1 U52 ( .A(n1634), .B(n1314), .Y(n1645) );
  AND2X1 U53 ( .A(n1315), .B(n1634), .Y(n1665) );
  AND2X1 U54 ( .A(n1321), .B(n1634), .Y(n1800) );
  AND2X1 U55 ( .A(\addr_1c<2> ), .B(n1031), .Y(n1595) );
  AND2X1 U56 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1634) );
  BUFX2 U57 ( .A(n961), .Y(n1010) );
  BUFX2 U58 ( .A(n961), .Y(n1009) );
  BUFX2 U59 ( .A(n960), .Y(n1007) );
  BUFX2 U60 ( .A(n960), .Y(n1006) );
  BUFX2 U61 ( .A(n959), .Y(n1004) );
  BUFX2 U62 ( .A(n959), .Y(n1003) );
  BUFX2 U63 ( .A(n958), .Y(n1001) );
  BUFX2 U64 ( .A(n958), .Y(n1000) );
  BUFX2 U65 ( .A(n957), .Y(n990) );
  BUFX2 U66 ( .A(n957), .Y(n989) );
  BUFX2 U67 ( .A(n956), .Y(n987) );
  BUFX2 U68 ( .A(n956), .Y(n986) );
  BUFX2 U69 ( .A(n955), .Y(n984) );
  BUFX2 U70 ( .A(n955), .Y(n983) );
  BUFX2 U71 ( .A(n954), .Y(n981) );
  BUFX2 U72 ( .A(n954), .Y(n980) );
  INVX1 U73 ( .A(\data_in_1c<0> ), .Y(n1034) );
  INVX1 U74 ( .A(\data_in_1c<1> ), .Y(n1035) );
  INVX1 U75 ( .A(\data_in_1c<2> ), .Y(n1036) );
  INVX1 U76 ( .A(\data_in_1c<3> ), .Y(n1037) );
  INVX1 U77 ( .A(\data_in_1c<4> ), .Y(n1038) );
  INVX1 U78 ( .A(\data_in_1c<5> ), .Y(n1039) );
  INVX1 U79 ( .A(\data_in_1c<6> ), .Y(n1040) );
  INVX1 U80 ( .A(\data_in_1c<7> ), .Y(n1041) );
  INVX1 U81 ( .A(\data_in_1c<8> ), .Y(n1042) );
  INVX1 U82 ( .A(\data_in_1c<9> ), .Y(n1043) );
  INVX1 U83 ( .A(\data_in_1c<10> ), .Y(n1044) );
  INVX1 U84 ( .A(\data_in_1c<11> ), .Y(n1045) );
  INVX1 U85 ( .A(\data_in_1c<12> ), .Y(n1046) );
  INVX1 U86 ( .A(\data_in_1c<13> ), .Y(n1047) );
  INVX1 U87 ( .A(\data_in_1c<14> ), .Y(n1048) );
  INVX1 U88 ( .A(\data_in_1c<15> ), .Y(n1049) );
  AND2X1 U89 ( .A(n1831), .B(\mem<32><0> ), .Y(n1495) );
  AND2X1 U90 ( .A(n1831), .B(\mem<32><1> ), .Y(n1507) );
  AND2X1 U91 ( .A(n1831), .B(\mem<32><2> ), .Y(n1340) );
  AND2X1 U92 ( .A(n1831), .B(\mem<32><3> ), .Y(n1353) );
  AND2X1 U93 ( .A(n1831), .B(\mem<32><4> ), .Y(n1366) );
  AND2X1 U129 ( .A(n1831), .B(\mem<32><5> ), .Y(n1379) );
  AND2X1 U589 ( .A(n1831), .B(\mem<32><6> ), .Y(n1392) );
  AND2X1 U640 ( .A(n1831), .B(\mem<32><7> ), .Y(n1405) );
  INVX1 U659 ( .A(rd1), .Y(n1028) );
  INVX1 U660 ( .A(n1017), .Y(n1016) );
  INVX1 U664 ( .A(wr), .Y(n1026) );
  INVX1 U666 ( .A(n1328), .Y(n1025) );
  INVX1 U672 ( .A(n1419), .Y(n1024) );
  INVX1 U675 ( .A(n1430), .Y(n1023) );
  INVX1 U679 ( .A(n1441), .Y(n1022) );
  INVX1 U682 ( .A(n1452), .Y(n1021) );
  INVX1 U694 ( .A(n1463), .Y(n1020) );
  INVX1 U697 ( .A(n1474), .Y(n1019) );
  INVX1 U701 ( .A(n1485), .Y(n1018) );
  INVX1 U706 ( .A(n1832), .Y(n1014) );
  AND2X1 U712 ( .A(wr1), .B(n1017), .Y(n1832) );
  INVX1 U717 ( .A(n1014), .Y(n1012) );
  INVX1 U723 ( .A(n1014), .Y(n1013) );
  AND2X1 U728 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U734 ( .A(n1), .Y(n2) );
  AND2X1 U739 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U745 ( .A(n3), .Y(n4) );
  AND2X1 U750 ( .A(n1821), .B(n189), .Y(n5) );
  INVX1 U756 ( .A(n5), .Y(n6) );
  AND2X1 U761 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U767 ( .A(n7), .Y(n8) );
  OR2X1 U772 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U786 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U789 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U801 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U804 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U816 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U819 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U831 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U834 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U846 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U849 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U861 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U864 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U870 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U875 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U882 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U883 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U884 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U885 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U886 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U887 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U888 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U889 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U890 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U891 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U892 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U893 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U894 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U895 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U896 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U897 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U898 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U899 ( .A(n973), .B(n1832), .Y(n189) );
  AND2X1 U900 ( .A(n1832), .B(n1528), .Y(n289) );
  AND2X1 U901 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U902 ( .A(n348), .Y(n372) );
  AND2X1 U903 ( .A(n950), .B(n952), .Y(n379) );
  INVX1 U904 ( .A(n379), .Y(n381) );
  AND2X1 U905 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U906 ( .A(n386), .Y(n387) );
  AND2X1 U907 ( .A(n950), .B(n951), .Y(n401) );
  INVX1 U908 ( .A(n401), .Y(n402) );
  BUFX2 U909 ( .A(n1343), .Y(n408) );
  BUFX2 U910 ( .A(n1356), .Y(n409) );
  BUFX2 U911 ( .A(n1369), .Y(n421) );
  BUFX2 U912 ( .A(n1382), .Y(n422) );
  BUFX2 U913 ( .A(n1395), .Y(n434) );
  BUFX2 U914 ( .A(n1408), .Y(n435) );
  BUFX2 U915 ( .A(n1498), .Y(n447) );
  BUFX2 U916 ( .A(n1509), .Y(n448) );
  AND2X2 U917 ( .A(rd), .B(n1512), .Y(n460) );
  INVX1 U918 ( .A(n460), .Y(n461) );
  INVX1 U919 ( .A(n1318), .Y(n473) );
  INVX1 U920 ( .A(n1319), .Y(n474) );
  INVX1 U921 ( .A(n1320), .Y(n486) );
  INVX1 U922 ( .A(n1411), .Y(n487) );
  INVX1 U923 ( .A(n1412), .Y(n507) );
  INVX1 U924 ( .A(n1413), .Y(n508) );
  INVX1 U925 ( .A(n1422), .Y(n522) );
  INVX1 U926 ( .A(n1423), .Y(n523) );
  INVX1 U927 ( .A(n1424), .Y(n537) );
  INVX1 U928 ( .A(n1433), .Y(n538) );
  INVX1 U929 ( .A(n1434), .Y(n552) );
  INVX1 U930 ( .A(n1435), .Y(n553) );
  INVX1 U931 ( .A(n1444), .Y(n567) );
  INVX1 U932 ( .A(n1445), .Y(n568) );
  INVX1 U933 ( .A(n1446), .Y(n582) );
  INVX1 U934 ( .A(n1455), .Y(n583) );
  INVX1 U935 ( .A(n1456), .Y(n591) );
  INVX1 U936 ( .A(n1457), .Y(n592) );
  INVX1 U937 ( .A(n1466), .Y(n871) );
  INVX1 U938 ( .A(n1467), .Y(n872) );
  INVX1 U939 ( .A(n1468), .Y(n873) );
  INVX1 U940 ( .A(n1477), .Y(n874) );
  INVX1 U941 ( .A(n1478), .Y(n875) );
  INVX1 U942 ( .A(n1479), .Y(n876) );
  AND2X2 U943 ( .A(n1332), .B(n1331), .Y(n877) );
  INVX1 U944 ( .A(n877), .Y(n878) );
  AND2X2 U945 ( .A(n1345), .B(n1344), .Y(n879) );
  INVX1 U946 ( .A(n879), .Y(n880) );
  AND2X2 U947 ( .A(n1358), .B(n1357), .Y(n881) );
  INVX1 U948 ( .A(n881), .Y(n882) );
  AND2X2 U949 ( .A(n1371), .B(n1370), .Y(n883) );
  INVX1 U950 ( .A(n883), .Y(n884) );
  AND2X2 U951 ( .A(n1384), .B(n1383), .Y(n885) );
  INVX1 U952 ( .A(n885), .Y(n886) );
  AND2X2 U953 ( .A(n1397), .B(n1396), .Y(n887) );
  INVX1 U954 ( .A(n887), .Y(n888) );
  AND2X2 U955 ( .A(n1487), .B(n1486), .Y(n889) );
  INVX1 U956 ( .A(n889), .Y(n890) );
  AND2X2 U957 ( .A(n1500), .B(n1499), .Y(n891) );
  INVX1 U958 ( .A(n891), .Y(n892) );
  INVX1 U959 ( .A(n1325), .Y(n893) );
  INVX1 U960 ( .A(n1326), .Y(n894) );
  INVX1 U961 ( .A(n1327), .Y(n895) );
  INVX1 U962 ( .A(n1416), .Y(n896) );
  INVX1 U963 ( .A(n1417), .Y(n897) );
  INVX1 U964 ( .A(n1418), .Y(n898) );
  INVX1 U965 ( .A(n1427), .Y(n899) );
  INVX1 U966 ( .A(n1428), .Y(n900) );
  INVX1 U967 ( .A(n1429), .Y(n901) );
  INVX1 U968 ( .A(n1438), .Y(n902) );
  INVX1 U969 ( .A(n1439), .Y(n903) );
  INVX1 U970 ( .A(n1440), .Y(n904) );
  INVX1 U971 ( .A(n1449), .Y(n905) );
  INVX1 U972 ( .A(n1450), .Y(n906) );
  INVX1 U973 ( .A(n1451), .Y(n907) );
  INVX1 U974 ( .A(n1460), .Y(n908) );
  INVX1 U975 ( .A(n1461), .Y(n909) );
  INVX1 U976 ( .A(n1462), .Y(n910) );
  INVX1 U977 ( .A(n1471), .Y(n911) );
  INVX1 U978 ( .A(n1472), .Y(n912) );
  INVX1 U979 ( .A(n1473), .Y(n913) );
  INVX1 U980 ( .A(n1482), .Y(n914) );
  INVX1 U981 ( .A(n1483), .Y(n915) );
  INVX1 U982 ( .A(n1484), .Y(n916) );
  AND2X2 U983 ( .A(n1334), .B(n1333), .Y(n917) );
  INVX1 U984 ( .A(n917), .Y(n918) );
  AND2X2 U985 ( .A(n1347), .B(n1346), .Y(n919) );
  INVX1 U986 ( .A(n919), .Y(n920) );
  AND2X2 U987 ( .A(n1360), .B(n1359), .Y(n921) );
  INVX1 U988 ( .A(n921), .Y(n922) );
  AND2X2 U989 ( .A(n1373), .B(n1372), .Y(n923) );
  INVX1 U990 ( .A(n923), .Y(n924) );
  AND2X2 U991 ( .A(n1386), .B(n1385), .Y(n925) );
  INVX1 U992 ( .A(n925), .Y(n926) );
  AND2X2 U993 ( .A(n1399), .B(n1398), .Y(n927) );
  INVX1 U994 ( .A(n927), .Y(n928) );
  AND2X2 U995 ( .A(n1489), .B(n1488), .Y(n929) );
  INVX1 U996 ( .A(n929), .Y(n930) );
  AND2X2 U997 ( .A(n1502), .B(n1501), .Y(n931) );
  INVX1 U998 ( .A(n931), .Y(n932) );
  BUFX2 U999 ( .A(n1341), .Y(n933) );
  BUFX2 U1000 ( .A(n1354), .Y(n934) );
  BUFX2 U1001 ( .A(n1367), .Y(n935) );
  BUFX2 U1002 ( .A(n1380), .Y(n936) );
  BUFX2 U1003 ( .A(n1393), .Y(n937) );
  BUFX2 U1004 ( .A(n1406), .Y(n938) );
  BUFX2 U1005 ( .A(n1496), .Y(n939) );
  INVX1 U1006 ( .A(n970), .Y(n940) );
  INVX1 U1007 ( .A(n1503), .Y(n941) );
  INVX1 U1008 ( .A(n1504), .Y(n942) );
  BUFX2 U1009 ( .A(n1556), .Y(n970) );
  BUFX2 U1010 ( .A(n1339), .Y(n943) );
  BUFX2 U1011 ( .A(n1352), .Y(n944) );
  BUFX2 U1012 ( .A(n1365), .Y(n945) );
  BUFX2 U1013 ( .A(n1378), .Y(n946) );
  BUFX2 U1014 ( .A(n1391), .Y(n947) );
  BUFX2 U1015 ( .A(n1404), .Y(n948) );
  BUFX2 U1016 ( .A(n1494), .Y(n949) );
  INVX1 U1017 ( .A(n971), .Y(n950) );
  INVX1 U1018 ( .A(n1505), .Y(n951) );
  INVX1 U1019 ( .A(n1506), .Y(n952) );
  BUFX2 U1020 ( .A(n1518), .Y(n971) );
  BUFX2 U1021 ( .A(n1842), .Y(err) );
  BUFX2 U1022 ( .A(n1527), .Y(n972) );
  BUFX2 U1023 ( .A(n1545), .Y(n974) );
  BUFX2 U1024 ( .A(n1555), .Y(n975) );
  BUFX2 U1025 ( .A(n1565), .Y(n976) );
  BUFX2 U1026 ( .A(n1575), .Y(n977) );
  BUFX2 U1027 ( .A(n1584), .Y(n978) );
  BUFX2 U1028 ( .A(n1594), .Y(n979) );
  BUFX2 U1029 ( .A(n1614), .Y(n982) );
  BUFX2 U1030 ( .A(n1633), .Y(n985) );
  BUFX2 U1031 ( .A(n1654), .Y(n988) );
  BUFX2 U1032 ( .A(n1674), .Y(n991) );
  BUFX2 U1033 ( .A(n1683), .Y(n992) );
  BUFX2 U1034 ( .A(n1693), .Y(n993) );
  BUFX2 U1035 ( .A(n1702), .Y(n994) );
  BUFX2 U1036 ( .A(n1712), .Y(n995) );
  BUFX2 U1037 ( .A(n1721), .Y(n996) );
  BUFX2 U1038 ( .A(n1731), .Y(n997) );
  BUFX2 U1039 ( .A(n1740), .Y(n998) );
  BUFX2 U1040 ( .A(n1750), .Y(n999) );
  BUFX2 U1041 ( .A(n1769), .Y(n1002) );
  BUFX2 U1042 ( .A(n1789), .Y(n1005) );
  BUFX2 U1043 ( .A(n1809), .Y(n1008) );
  BUFX2 U1044 ( .A(n1822), .Y(n973) );
  AND2X1 U1045 ( .A(n1634), .B(n1322), .Y(n1821) );
  BUFX2 U1046 ( .A(n1841), .Y(n1011) );
  BUFX2 U1047 ( .A(n1604), .Y(n954) );
  BUFX2 U1048 ( .A(n1623), .Y(n955) );
  BUFX2 U1049 ( .A(n1644), .Y(n956) );
  BUFX2 U1050 ( .A(n1664), .Y(n957) );
  BUFX2 U1051 ( .A(n1759), .Y(n958) );
  BUFX2 U1052 ( .A(n1779), .Y(n959) );
  BUFX2 U1053 ( .A(n1799), .Y(n960) );
  BUFX2 U1054 ( .A(n1820), .Y(n961) );
  AND2X1 U1055 ( .A(enable), .B(n1017), .Y(n962) );
  INVX1 U1056 ( .A(n962), .Y(n963) );
  INVX1 U1057 ( .A(n965), .Y(n964) );
  AND2X1 U1058 ( .A(n1517), .B(n1516), .Y(n965) );
  INVX1 U1059 ( .A(n966), .Y(n967) );
  INVX1 U1060 ( .A(n968), .Y(n969) );
  AND2X1 U1061 ( .A(n950), .B(n1314), .Y(n1528) );
endmodule


module final_memory_0 ( .data_out({\data_out<15> , \data_out<14> , 
        \data_out<13> , \data_out<12> , \data_out<11> , \data_out<10> , 
        \data_out<9> , \data_out<8> , \data_out<7> , \data_out<6> , 
        \data_out<5> , \data_out<4> , \data_out<3> , \data_out<2> , 
        \data_out<1> , \data_out<0> }), err, .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<12> , \addr<11> , \addr<10> , \addr<9> , 
        \addr<8> , \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , 
        \addr<2> , \addr<1> , \addr<0> }), wr, rd, enable, create_dump, 
    .bank_id({\bank_id<1> , \bank_id<0> }), clk, rst );
  input \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , \addr<12> , \addr<11> ,
         \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> , \addr<5> ,
         \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> , wr, rd, enable,
         create_dump, \bank_id<1> , \bank_id<0> , clk, rst;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , err;
  wire   n1840, rd0, wr0, rd1, wr1, \addr_1c<12> , \addr_1c<11> ,
         \addr_1c<10> , \addr_1c<9> , \addr_1c<8> , \addr_1c<7> , \addr_1c<6> ,
         \addr_1c<5> , \addr_1c<4> , \addr_1c<3> , \addr_1c<2> , \addr_1c<1> ,
         \addr_1c<0> , \data_in_1c<15> , \data_in_1c<14> , \data_in_1c<13> ,
         \data_in_1c<12> , \data_in_1c<11> , \data_in_1c<10> , \data_in_1c<9> ,
         \data_in_1c<8> , \data_in_1c<7> , \data_in_1c<6> , \data_in_1c<5> ,
         \data_in_1c<4> , \data_in_1c<3> , \data_in_1c<2> , \data_in_1c<1> ,
         \data_in_1c<0> , \mem<0><7> , \mem<0><6> , \mem<0><5> , \mem<0><4> ,
         \mem<0><3> , \mem<0><2> , \mem<0><1> , \mem<0><0> , \mem<1><7> ,
         \mem<1><6> , \mem<1><5> , \mem<1><4> , \mem<1><3> , \mem<1><2> ,
         \mem<1><1> , \mem<1><0> , \mem<2><7> , \mem<2><6> , \mem<2><5> ,
         \mem<2><4> , \mem<2><3> , \mem<2><2> , \mem<2><1> , \mem<2><0> ,
         \mem<3><7> , \mem<3><6> , \mem<3><5> , \mem<3><4> , \mem<3><3> ,
         \mem<3><2> , \mem<3><1> , \mem<3><0> , \mem<4><7> , \mem<4><6> ,
         \mem<4><5> , \mem<4><4> , \mem<4><3> , \mem<4><2> , \mem<4><1> ,
         \mem<4><0> , \mem<5><7> , \mem<5><6> , \mem<5><5> , \mem<5><4> ,
         \mem<5><3> , \mem<5><2> , \mem<5><1> , \mem<5><0> , \mem<6><7> ,
         \mem<6><6> , \mem<6><5> , \mem<6><4> , \mem<6><3> , \mem<6><2> ,
         \mem<6><1> , \mem<6><0> , \mem<7><7> , \mem<7><6> , \mem<7><5> ,
         \mem<7><4> , \mem<7><3> , \mem<7><2> , \mem<7><1> , \mem<7><0> ,
         \mem<8><7> , \mem<8><6> , \mem<8><5> , \mem<8><4> , \mem<8><3> ,
         \mem<8><2> , \mem<8><1> , \mem<8><0> , \mem<9><7> , \mem<9><6> ,
         \mem<9><5> , \mem<9><4> , \mem<9><3> , \mem<9><2> , \mem<9><1> ,
         \mem<9><0> , \mem<10><7> , \mem<10><6> , \mem<10><5> , \mem<10><4> ,
         \mem<10><3> , \mem<10><2> , \mem<10><1> , \mem<10><0> , \mem<11><7> ,
         \mem<11><6> , \mem<11><5> , \mem<11><4> , \mem<11><3> , \mem<11><2> ,
         \mem<11><1> , \mem<11><0> , \mem<12><7> , \mem<12><6> , \mem<12><5> ,
         \mem<12><4> , \mem<12><3> , \mem<12><2> , \mem<12><1> , \mem<12><0> ,
         \mem<13><7> , \mem<13><6> , \mem<13><5> , \mem<13><4> , \mem<13><3> ,
         \mem<13><2> , \mem<13><1> , \mem<13><0> , \mem<14><7> , \mem<14><6> ,
         \mem<14><5> , \mem<14><4> , \mem<14><3> , \mem<14><2> , \mem<14><1> ,
         \mem<14><0> , \mem<15><7> , \mem<15><6> , \mem<15><5> , \mem<15><4> ,
         \mem<15><3> , \mem<15><2> , \mem<15><1> , \mem<15><0> , \mem<16><7> ,
         \mem<16><6> , \mem<16><5> , \mem<16><4> , \mem<16><3> , \mem<16><2> ,
         \mem<16><1> , \mem<16><0> , \mem<17><7> , \mem<17><6> , \mem<17><5> ,
         \mem<17><4> , \mem<17><3> , \mem<17><2> , \mem<17><1> , \mem<17><0> ,
         \mem<18><7> , \mem<18><6> , \mem<18><5> , \mem<18><4> , \mem<18><3> ,
         \mem<18><2> , \mem<18><1> , \mem<18><0> , \mem<19><7> , \mem<19><6> ,
         \mem<19><5> , \mem<19><4> , \mem<19><3> , \mem<19><2> , \mem<19><1> ,
         \mem<19><0> , \mem<20><7> , \mem<20><6> , \mem<20><5> , \mem<20><4> ,
         \mem<20><3> , \mem<20><2> , \mem<20><1> , \mem<20><0> , \mem<21><7> ,
         \mem<21><6> , \mem<21><5> , \mem<21><4> , \mem<21><3> , \mem<21><2> ,
         \mem<21><1> , \mem<21><0> , \mem<22><7> , \mem<22><6> , \mem<22><5> ,
         \mem<22><4> , \mem<22><3> , \mem<22><2> , \mem<22><1> , \mem<22><0> ,
         \mem<23><7> , \mem<23><6> , \mem<23><5> , \mem<23><4> , \mem<23><3> ,
         \mem<23><2> , \mem<23><1> , \mem<23><0> , \mem<24><7> , \mem<24><6> ,
         \mem<24><5> , \mem<24><4> , \mem<24><3> , \mem<24><2> , \mem<24><1> ,
         \mem<24><0> , \mem<25><7> , \mem<25><6> , \mem<25><5> , \mem<25><4> ,
         \mem<25><3> , \mem<25><2> , \mem<25><1> , \mem<25><0> , \mem<26><7> ,
         \mem<26><6> , \mem<26><5> , \mem<26><4> , \mem<26><3> , \mem<26><2> ,
         \mem<26><1> , \mem<26><0> , \mem<27><7> , \mem<27><6> , \mem<27><5> ,
         \mem<27><4> , \mem<27><3> , \mem<27><2> , \mem<27><1> , \mem<27><0> ,
         \mem<28><7> , \mem<28><6> , \mem<28><5> , \mem<28><4> , \mem<28><3> ,
         \mem<28><2> , \mem<28><1> , \mem<28><0> , \mem<29><7> , \mem<29><6> ,
         \mem<29><5> , \mem<29><4> , \mem<29><3> , \mem<29><2> , \mem<29><1> ,
         \mem<29><0> , \mem<30><7> , \mem<30><6> , \mem<30><5> , \mem<30><4> ,
         \mem<30><3> , \mem<30><2> , \mem<30><1> , \mem<30><0> , \mem<31><7> ,
         \mem<31><6> , \mem<31><5> , \mem<31><4> , \mem<31><3> , \mem<31><2> ,
         \mem<31><1> , \mem<31><0> , \mem<32><7> , \mem<32><6> , \mem<32><5> ,
         \mem<32><4> , \mem<32><3> , \mem<32><2> , \mem<32><1> , \mem<32><0> ,
         \data_out_1c<15> , \data_out_1c<14> , \data_out_1c<13> ,
         \data_out_1c<12> , \data_out_1c<11> , \data_out_1c<10> ,
         \data_out_1c<9> , \data_out_1c<8> , rd2, wr2, rd3, wr3, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n50, n150, n189, n289, n348, n372, n379,
         n381, n386, n387, n401, n402, n408, n409, n421, n422, n434, n435,
         n447, n448, n460, n461, n473, n474, n486, n487, n507, n508, n522,
         n523, n537, n538, n552, n553, n567, n568, n582, n583, n591, n592,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839;

  DFFPOSX1 \mem_reg<0><7>  ( .D(n1048), .CLK(clk), .Q(\mem<0><7> ) );
  DFFPOSX1 \mem_reg<0><6>  ( .D(n1049), .CLK(clk), .Q(\mem<0><6> ) );
  DFFPOSX1 \mem_reg<0><5>  ( .D(n1050), .CLK(clk), .Q(\mem<0><5> ) );
  DFFPOSX1 \mem_reg<0><4>  ( .D(n1051), .CLK(clk), .Q(\mem<0><4> ) );
  DFFPOSX1 \mem_reg<0><3>  ( .D(n1052), .CLK(clk), .Q(\mem<0><3> ) );
  DFFPOSX1 \mem_reg<0><2>  ( .D(n1053), .CLK(clk), .Q(\mem<0><2> ) );
  DFFPOSX1 \mem_reg<0><1>  ( .D(n1054), .CLK(clk), .Q(\mem<0><1> ) );
  DFFPOSX1 \mem_reg<0><0>  ( .D(n1055), .CLK(clk), .Q(\mem<0><0> ) );
  DFFPOSX1 \mem_reg<1><7>  ( .D(n1056), .CLK(clk), .Q(\mem<1><7> ) );
  DFFPOSX1 \mem_reg<1><6>  ( .D(n1057), .CLK(clk), .Q(\mem<1><6> ) );
  DFFPOSX1 \mem_reg<1><5>  ( .D(n1058), .CLK(clk), .Q(\mem<1><5> ) );
  DFFPOSX1 \mem_reg<1><4>  ( .D(n1059), .CLK(clk), .Q(\mem<1><4> ) );
  DFFPOSX1 \mem_reg<1><3>  ( .D(n1060), .CLK(clk), .Q(\mem<1><3> ) );
  DFFPOSX1 \mem_reg<1><2>  ( .D(n1061), .CLK(clk), .Q(\mem<1><2> ) );
  DFFPOSX1 \mem_reg<1><1>  ( .D(n1062), .CLK(clk), .Q(\mem<1><1> ) );
  DFFPOSX1 \mem_reg<1><0>  ( .D(n1063), .CLK(clk), .Q(\mem<1><0> ) );
  DFFPOSX1 \mem_reg<2><7>  ( .D(n1064), .CLK(clk), .Q(\mem<2><7> ) );
  DFFPOSX1 \mem_reg<2><6>  ( .D(n1065), .CLK(clk), .Q(\mem<2><6> ) );
  DFFPOSX1 \mem_reg<2><5>  ( .D(n1066), .CLK(clk), .Q(\mem<2><5> ) );
  DFFPOSX1 \mem_reg<2><4>  ( .D(n1067), .CLK(clk), .Q(\mem<2><4> ) );
  DFFPOSX1 \mem_reg<2><3>  ( .D(n1068), .CLK(clk), .Q(\mem<2><3> ) );
  DFFPOSX1 \mem_reg<2><2>  ( .D(n1069), .CLK(clk), .Q(\mem<2><2> ) );
  DFFPOSX1 \mem_reg<2><1>  ( .D(n1070), .CLK(clk), .Q(\mem<2><1> ) );
  DFFPOSX1 \mem_reg<2><0>  ( .D(n1071), .CLK(clk), .Q(\mem<2><0> ) );
  DFFPOSX1 \mem_reg<3><7>  ( .D(n1072), .CLK(clk), .Q(\mem<3><7> ) );
  DFFPOSX1 \mem_reg<3><6>  ( .D(n1073), .CLK(clk), .Q(\mem<3><6> ) );
  DFFPOSX1 \mem_reg<3><5>  ( .D(n1074), .CLK(clk), .Q(\mem<3><5> ) );
  DFFPOSX1 \mem_reg<3><4>  ( .D(n1075), .CLK(clk), .Q(\mem<3><4> ) );
  DFFPOSX1 \mem_reg<3><3>  ( .D(n1076), .CLK(clk), .Q(\mem<3><3> ) );
  DFFPOSX1 \mem_reg<3><2>  ( .D(n1077), .CLK(clk), .Q(\mem<3><2> ) );
  DFFPOSX1 \mem_reg<3><1>  ( .D(n1078), .CLK(clk), .Q(\mem<3><1> ) );
  DFFPOSX1 \mem_reg<3><0>  ( .D(n1079), .CLK(clk), .Q(\mem<3><0> ) );
  DFFPOSX1 \mem_reg<4><7>  ( .D(n1080), .CLK(clk), .Q(\mem<4><7> ) );
  DFFPOSX1 \mem_reg<4><6>  ( .D(n1081), .CLK(clk), .Q(\mem<4><6> ) );
  DFFPOSX1 \mem_reg<4><5>  ( .D(n1082), .CLK(clk), .Q(\mem<4><5> ) );
  DFFPOSX1 \mem_reg<4><4>  ( .D(n1083), .CLK(clk), .Q(\mem<4><4> ) );
  DFFPOSX1 \mem_reg<4><3>  ( .D(n1084), .CLK(clk), .Q(\mem<4><3> ) );
  DFFPOSX1 \mem_reg<4><2>  ( .D(n1085), .CLK(clk), .Q(\mem<4><2> ) );
  DFFPOSX1 \mem_reg<4><1>  ( .D(n1086), .CLK(clk), .Q(\mem<4><1> ) );
  DFFPOSX1 \mem_reg<4><0>  ( .D(n1087), .CLK(clk), .Q(\mem<4><0> ) );
  DFFPOSX1 \mem_reg<5><7>  ( .D(n1088), .CLK(clk), .Q(\mem<5><7> ) );
  DFFPOSX1 \mem_reg<5><6>  ( .D(n1089), .CLK(clk), .Q(\mem<5><6> ) );
  DFFPOSX1 \mem_reg<5><5>  ( .D(n1090), .CLK(clk), .Q(\mem<5><5> ) );
  DFFPOSX1 \mem_reg<5><4>  ( .D(n1091), .CLK(clk), .Q(\mem<5><4> ) );
  DFFPOSX1 \mem_reg<5><3>  ( .D(n1092), .CLK(clk), .Q(\mem<5><3> ) );
  DFFPOSX1 \mem_reg<5><2>  ( .D(n1093), .CLK(clk), .Q(\mem<5><2> ) );
  DFFPOSX1 \mem_reg<5><1>  ( .D(n1094), .CLK(clk), .Q(\mem<5><1> ) );
  DFFPOSX1 \mem_reg<5><0>  ( .D(n1095), .CLK(clk), .Q(\mem<5><0> ) );
  DFFPOSX1 \mem_reg<6><7>  ( .D(n1096), .CLK(clk), .Q(\mem<6><7> ) );
  DFFPOSX1 \mem_reg<6><6>  ( .D(n1097), .CLK(clk), .Q(\mem<6><6> ) );
  DFFPOSX1 \mem_reg<6><5>  ( .D(n1098), .CLK(clk), .Q(\mem<6><5> ) );
  DFFPOSX1 \mem_reg<6><4>  ( .D(n1099), .CLK(clk), .Q(\mem<6><4> ) );
  DFFPOSX1 \mem_reg<6><3>  ( .D(n1100), .CLK(clk), .Q(\mem<6><3> ) );
  DFFPOSX1 \mem_reg<6><2>  ( .D(n1101), .CLK(clk), .Q(\mem<6><2> ) );
  DFFPOSX1 \mem_reg<6><1>  ( .D(n1102), .CLK(clk), .Q(\mem<6><1> ) );
  DFFPOSX1 \mem_reg<6><0>  ( .D(n1103), .CLK(clk), .Q(\mem<6><0> ) );
  DFFPOSX1 \mem_reg<7><7>  ( .D(n1104), .CLK(clk), .Q(\mem<7><7> ) );
  DFFPOSX1 \mem_reg<7><6>  ( .D(n1105), .CLK(clk), .Q(\mem<7><6> ) );
  DFFPOSX1 \mem_reg<7><5>  ( .D(n1106), .CLK(clk), .Q(\mem<7><5> ) );
  DFFPOSX1 \mem_reg<7><4>  ( .D(n1107), .CLK(clk), .Q(\mem<7><4> ) );
  DFFPOSX1 \mem_reg<7><3>  ( .D(n1108), .CLK(clk), .Q(\mem<7><3> ) );
  DFFPOSX1 \mem_reg<7><2>  ( .D(n1109), .CLK(clk), .Q(\mem<7><2> ) );
  DFFPOSX1 \mem_reg<7><1>  ( .D(n1110), .CLK(clk), .Q(\mem<7><1> ) );
  DFFPOSX1 \mem_reg<7><0>  ( .D(n1111), .CLK(clk), .Q(\mem<7><0> ) );
  DFFPOSX1 \mem_reg<8><7>  ( .D(n1112), .CLK(clk), .Q(\mem<8><7> ) );
  DFFPOSX1 \mem_reg<8><6>  ( .D(n1113), .CLK(clk), .Q(\mem<8><6> ) );
  DFFPOSX1 \mem_reg<8><5>  ( .D(n1114), .CLK(clk), .Q(\mem<8><5> ) );
  DFFPOSX1 \mem_reg<8><4>  ( .D(n1115), .CLK(clk), .Q(\mem<8><4> ) );
  DFFPOSX1 \mem_reg<8><3>  ( .D(n1116), .CLK(clk), .Q(\mem<8><3> ) );
  DFFPOSX1 \mem_reg<8><2>  ( .D(n1117), .CLK(clk), .Q(\mem<8><2> ) );
  DFFPOSX1 \mem_reg<8><1>  ( .D(n1118), .CLK(clk), .Q(\mem<8><1> ) );
  DFFPOSX1 \mem_reg<8><0>  ( .D(n1119), .CLK(clk), .Q(\mem<8><0> ) );
  DFFPOSX1 \mem_reg<9><7>  ( .D(n1120), .CLK(clk), .Q(\mem<9><7> ) );
  DFFPOSX1 \mem_reg<9><6>  ( .D(n1121), .CLK(clk), .Q(\mem<9><6> ) );
  DFFPOSX1 \mem_reg<9><5>  ( .D(n1122), .CLK(clk), .Q(\mem<9><5> ) );
  DFFPOSX1 \mem_reg<9><4>  ( .D(n1123), .CLK(clk), .Q(\mem<9><4> ) );
  DFFPOSX1 \mem_reg<9><3>  ( .D(n1124), .CLK(clk), .Q(\mem<9><3> ) );
  DFFPOSX1 \mem_reg<9><2>  ( .D(n1125), .CLK(clk), .Q(\mem<9><2> ) );
  DFFPOSX1 \mem_reg<9><1>  ( .D(n1126), .CLK(clk), .Q(\mem<9><1> ) );
  DFFPOSX1 \mem_reg<9><0>  ( .D(n1127), .CLK(clk), .Q(\mem<9><0> ) );
  DFFPOSX1 \mem_reg<10><7>  ( .D(n1128), .CLK(clk), .Q(\mem<10><7> ) );
  DFFPOSX1 \mem_reg<10><6>  ( .D(n1129), .CLK(clk), .Q(\mem<10><6> ) );
  DFFPOSX1 \mem_reg<10><5>  ( .D(n1130), .CLK(clk), .Q(\mem<10><5> ) );
  DFFPOSX1 \mem_reg<10><4>  ( .D(n1131), .CLK(clk), .Q(\mem<10><4> ) );
  DFFPOSX1 \mem_reg<10><3>  ( .D(n1132), .CLK(clk), .Q(\mem<10><3> ) );
  DFFPOSX1 \mem_reg<10><2>  ( .D(n1133), .CLK(clk), .Q(\mem<10><2> ) );
  DFFPOSX1 \mem_reg<10><1>  ( .D(n1134), .CLK(clk), .Q(\mem<10><1> ) );
  DFFPOSX1 \mem_reg<10><0>  ( .D(n1135), .CLK(clk), .Q(\mem<10><0> ) );
  DFFPOSX1 \mem_reg<11><7>  ( .D(n1136), .CLK(clk), .Q(\mem<11><7> ) );
  DFFPOSX1 \mem_reg<11><6>  ( .D(n1137), .CLK(clk), .Q(\mem<11><6> ) );
  DFFPOSX1 \mem_reg<11><5>  ( .D(n1138), .CLK(clk), .Q(\mem<11><5> ) );
  DFFPOSX1 \mem_reg<11><4>  ( .D(n1139), .CLK(clk), .Q(\mem<11><4> ) );
  DFFPOSX1 \mem_reg<11><3>  ( .D(n1140), .CLK(clk), .Q(\mem<11><3> ) );
  DFFPOSX1 \mem_reg<11><2>  ( .D(n1141), .CLK(clk), .Q(\mem<11><2> ) );
  DFFPOSX1 \mem_reg<11><1>  ( .D(n1142), .CLK(clk), .Q(\mem<11><1> ) );
  DFFPOSX1 \mem_reg<11><0>  ( .D(n1143), .CLK(clk), .Q(\mem<11><0> ) );
  DFFPOSX1 \mem_reg<12><7>  ( .D(n1144), .CLK(clk), .Q(\mem<12><7> ) );
  DFFPOSX1 \mem_reg<12><6>  ( .D(n1145), .CLK(clk), .Q(\mem<12><6> ) );
  DFFPOSX1 \mem_reg<12><5>  ( .D(n1146), .CLK(clk), .Q(\mem<12><5> ) );
  DFFPOSX1 \mem_reg<12><4>  ( .D(n1147), .CLK(clk), .Q(\mem<12><4> ) );
  DFFPOSX1 \mem_reg<12><3>  ( .D(n1148), .CLK(clk), .Q(\mem<12><3> ) );
  DFFPOSX1 \mem_reg<12><2>  ( .D(n1149), .CLK(clk), .Q(\mem<12><2> ) );
  DFFPOSX1 \mem_reg<12><1>  ( .D(n1150), .CLK(clk), .Q(\mem<12><1> ) );
  DFFPOSX1 \mem_reg<12><0>  ( .D(n1151), .CLK(clk), .Q(\mem<12><0> ) );
  DFFPOSX1 \mem_reg<13><7>  ( .D(n1152), .CLK(clk), .Q(\mem<13><7> ) );
  DFFPOSX1 \mem_reg<13><6>  ( .D(n1153), .CLK(clk), .Q(\mem<13><6> ) );
  DFFPOSX1 \mem_reg<13><5>  ( .D(n1154), .CLK(clk), .Q(\mem<13><5> ) );
  DFFPOSX1 \mem_reg<13><4>  ( .D(n1155), .CLK(clk), .Q(\mem<13><4> ) );
  DFFPOSX1 \mem_reg<13><3>  ( .D(n1156), .CLK(clk), .Q(\mem<13><3> ) );
  DFFPOSX1 \mem_reg<13><2>  ( .D(n1157), .CLK(clk), .Q(\mem<13><2> ) );
  DFFPOSX1 \mem_reg<13><1>  ( .D(n1158), .CLK(clk), .Q(\mem<13><1> ) );
  DFFPOSX1 \mem_reg<13><0>  ( .D(n1159), .CLK(clk), .Q(\mem<13><0> ) );
  DFFPOSX1 \mem_reg<14><7>  ( .D(n1160), .CLK(clk), .Q(\mem<14><7> ) );
  DFFPOSX1 \mem_reg<14><6>  ( .D(n1161), .CLK(clk), .Q(\mem<14><6> ) );
  DFFPOSX1 \mem_reg<14><5>  ( .D(n1162), .CLK(clk), .Q(\mem<14><5> ) );
  DFFPOSX1 \mem_reg<14><4>  ( .D(n1163), .CLK(clk), .Q(\mem<14><4> ) );
  DFFPOSX1 \mem_reg<14><3>  ( .D(n1164), .CLK(clk), .Q(\mem<14><3> ) );
  DFFPOSX1 \mem_reg<14><2>  ( .D(n1165), .CLK(clk), .Q(\mem<14><2> ) );
  DFFPOSX1 \mem_reg<14><1>  ( .D(n1166), .CLK(clk), .Q(\mem<14><1> ) );
  DFFPOSX1 \mem_reg<14><0>  ( .D(n1167), .CLK(clk), .Q(\mem<14><0> ) );
  DFFPOSX1 \mem_reg<15><7>  ( .D(n1168), .CLK(clk), .Q(\mem<15><7> ) );
  DFFPOSX1 \mem_reg<15><6>  ( .D(n1169), .CLK(clk), .Q(\mem<15><6> ) );
  DFFPOSX1 \mem_reg<15><5>  ( .D(n1170), .CLK(clk), .Q(\mem<15><5> ) );
  DFFPOSX1 \mem_reg<15><4>  ( .D(n1171), .CLK(clk), .Q(\mem<15><4> ) );
  DFFPOSX1 \mem_reg<15><3>  ( .D(n1172), .CLK(clk), .Q(\mem<15><3> ) );
  DFFPOSX1 \mem_reg<15><2>  ( .D(n1173), .CLK(clk), .Q(\mem<15><2> ) );
  DFFPOSX1 \mem_reg<15><1>  ( .D(n1174), .CLK(clk), .Q(\mem<15><1> ) );
  DFFPOSX1 \mem_reg<15><0>  ( .D(n1175), .CLK(clk), .Q(\mem<15><0> ) );
  DFFPOSX1 \mem_reg<16><7>  ( .D(n1176), .CLK(clk), .Q(\mem<16><7> ) );
  DFFPOSX1 \mem_reg<16><6>  ( .D(n1177), .CLK(clk), .Q(\mem<16><6> ) );
  DFFPOSX1 \mem_reg<16><5>  ( .D(n1178), .CLK(clk), .Q(\mem<16><5> ) );
  DFFPOSX1 \mem_reg<16><4>  ( .D(n1179), .CLK(clk), .Q(\mem<16><4> ) );
  DFFPOSX1 \mem_reg<16><3>  ( .D(n1180), .CLK(clk), .Q(\mem<16><3> ) );
  DFFPOSX1 \mem_reg<16><2>  ( .D(n1181), .CLK(clk), .Q(\mem<16><2> ) );
  DFFPOSX1 \mem_reg<16><1>  ( .D(n1182), .CLK(clk), .Q(\mem<16><1> ) );
  DFFPOSX1 \mem_reg<16><0>  ( .D(n1183), .CLK(clk), .Q(\mem<16><0> ) );
  DFFPOSX1 \mem_reg<17><7>  ( .D(n1184), .CLK(clk), .Q(\mem<17><7> ) );
  DFFPOSX1 \mem_reg<17><6>  ( .D(n1185), .CLK(clk), .Q(\mem<17><6> ) );
  DFFPOSX1 \mem_reg<17><5>  ( .D(n1186), .CLK(clk), .Q(\mem<17><5> ) );
  DFFPOSX1 \mem_reg<17><4>  ( .D(n1187), .CLK(clk), .Q(\mem<17><4> ) );
  DFFPOSX1 \mem_reg<17><3>  ( .D(n1188), .CLK(clk), .Q(\mem<17><3> ) );
  DFFPOSX1 \mem_reg<17><2>  ( .D(n1189), .CLK(clk), .Q(\mem<17><2> ) );
  DFFPOSX1 \mem_reg<17><1>  ( .D(n1190), .CLK(clk), .Q(\mem<17><1> ) );
  DFFPOSX1 \mem_reg<17><0>  ( .D(n1191), .CLK(clk), .Q(\mem<17><0> ) );
  DFFPOSX1 \mem_reg<18><7>  ( .D(n1192), .CLK(clk), .Q(\mem<18><7> ) );
  DFFPOSX1 \mem_reg<18><6>  ( .D(n1193), .CLK(clk), .Q(\mem<18><6> ) );
  DFFPOSX1 \mem_reg<18><5>  ( .D(n1194), .CLK(clk), .Q(\mem<18><5> ) );
  DFFPOSX1 \mem_reg<18><4>  ( .D(n1195), .CLK(clk), .Q(\mem<18><4> ) );
  DFFPOSX1 \mem_reg<18><3>  ( .D(n1196), .CLK(clk), .Q(\mem<18><3> ) );
  DFFPOSX1 \mem_reg<18><2>  ( .D(n1197), .CLK(clk), .Q(\mem<18><2> ) );
  DFFPOSX1 \mem_reg<18><1>  ( .D(n1198), .CLK(clk), .Q(\mem<18><1> ) );
  DFFPOSX1 \mem_reg<18><0>  ( .D(n1199), .CLK(clk), .Q(\mem<18><0> ) );
  DFFPOSX1 \mem_reg<19><7>  ( .D(n1200), .CLK(clk), .Q(\mem<19><7> ) );
  DFFPOSX1 \mem_reg<19><6>  ( .D(n1201), .CLK(clk), .Q(\mem<19><6> ) );
  DFFPOSX1 \mem_reg<19><5>  ( .D(n1202), .CLK(clk), .Q(\mem<19><5> ) );
  DFFPOSX1 \mem_reg<19><4>  ( .D(n1203), .CLK(clk), .Q(\mem<19><4> ) );
  DFFPOSX1 \mem_reg<19><3>  ( .D(n1204), .CLK(clk), .Q(\mem<19><3> ) );
  DFFPOSX1 \mem_reg<19><2>  ( .D(n1205), .CLK(clk), .Q(\mem<19><2> ) );
  DFFPOSX1 \mem_reg<19><1>  ( .D(n1206), .CLK(clk), .Q(\mem<19><1> ) );
  DFFPOSX1 \mem_reg<19><0>  ( .D(n1207), .CLK(clk), .Q(\mem<19><0> ) );
  DFFPOSX1 \mem_reg<20><7>  ( .D(n1208), .CLK(clk), .Q(\mem<20><7> ) );
  DFFPOSX1 \mem_reg<20><6>  ( .D(n1209), .CLK(clk), .Q(\mem<20><6> ) );
  DFFPOSX1 \mem_reg<20><5>  ( .D(n1210), .CLK(clk), .Q(\mem<20><5> ) );
  DFFPOSX1 \mem_reg<20><4>  ( .D(n1211), .CLK(clk), .Q(\mem<20><4> ) );
  DFFPOSX1 \mem_reg<20><3>  ( .D(n1212), .CLK(clk), .Q(\mem<20><3> ) );
  DFFPOSX1 \mem_reg<20><2>  ( .D(n1213), .CLK(clk), .Q(\mem<20><2> ) );
  DFFPOSX1 \mem_reg<20><1>  ( .D(n1214), .CLK(clk), .Q(\mem<20><1> ) );
  DFFPOSX1 \mem_reg<20><0>  ( .D(n1215), .CLK(clk), .Q(\mem<20><0> ) );
  DFFPOSX1 \mem_reg<21><7>  ( .D(n1216), .CLK(clk), .Q(\mem<21><7> ) );
  DFFPOSX1 \mem_reg<21><6>  ( .D(n1217), .CLK(clk), .Q(\mem<21><6> ) );
  DFFPOSX1 \mem_reg<21><5>  ( .D(n1218), .CLK(clk), .Q(\mem<21><5> ) );
  DFFPOSX1 \mem_reg<21><4>  ( .D(n1219), .CLK(clk), .Q(\mem<21><4> ) );
  DFFPOSX1 \mem_reg<21><3>  ( .D(n1220), .CLK(clk), .Q(\mem<21><3> ) );
  DFFPOSX1 \mem_reg<21><2>  ( .D(n1221), .CLK(clk), .Q(\mem<21><2> ) );
  DFFPOSX1 \mem_reg<21><1>  ( .D(n1222), .CLK(clk), .Q(\mem<21><1> ) );
  DFFPOSX1 \mem_reg<21><0>  ( .D(n1223), .CLK(clk), .Q(\mem<21><0> ) );
  DFFPOSX1 \mem_reg<22><7>  ( .D(n1224), .CLK(clk), .Q(\mem<22><7> ) );
  DFFPOSX1 \mem_reg<22><6>  ( .D(n1225), .CLK(clk), .Q(\mem<22><6> ) );
  DFFPOSX1 \mem_reg<22><5>  ( .D(n1226), .CLK(clk), .Q(\mem<22><5> ) );
  DFFPOSX1 \mem_reg<22><4>  ( .D(n1227), .CLK(clk), .Q(\mem<22><4> ) );
  DFFPOSX1 \mem_reg<22><3>  ( .D(n1228), .CLK(clk), .Q(\mem<22><3> ) );
  DFFPOSX1 \mem_reg<22><2>  ( .D(n1229), .CLK(clk), .Q(\mem<22><2> ) );
  DFFPOSX1 \mem_reg<22><1>  ( .D(n1230), .CLK(clk), .Q(\mem<22><1> ) );
  DFFPOSX1 \mem_reg<22><0>  ( .D(n1231), .CLK(clk), .Q(\mem<22><0> ) );
  DFFPOSX1 \mem_reg<23><7>  ( .D(n1232), .CLK(clk), .Q(\mem<23><7> ) );
  DFFPOSX1 \mem_reg<23><6>  ( .D(n1233), .CLK(clk), .Q(\mem<23><6> ) );
  DFFPOSX1 \mem_reg<23><5>  ( .D(n1234), .CLK(clk), .Q(\mem<23><5> ) );
  DFFPOSX1 \mem_reg<23><4>  ( .D(n1235), .CLK(clk), .Q(\mem<23><4> ) );
  DFFPOSX1 \mem_reg<23><3>  ( .D(n1236), .CLK(clk), .Q(\mem<23><3> ) );
  DFFPOSX1 \mem_reg<23><2>  ( .D(n1237), .CLK(clk), .Q(\mem<23><2> ) );
  DFFPOSX1 \mem_reg<23><1>  ( .D(n1238), .CLK(clk), .Q(\mem<23><1> ) );
  DFFPOSX1 \mem_reg<23><0>  ( .D(n1239), .CLK(clk), .Q(\mem<23><0> ) );
  DFFPOSX1 \mem_reg<24><7>  ( .D(n1240), .CLK(clk), .Q(\mem<24><7> ) );
  DFFPOSX1 \mem_reg<24><6>  ( .D(n1241), .CLK(clk), .Q(\mem<24><6> ) );
  DFFPOSX1 \mem_reg<24><5>  ( .D(n1242), .CLK(clk), .Q(\mem<24><5> ) );
  DFFPOSX1 \mem_reg<24><4>  ( .D(n1243), .CLK(clk), .Q(\mem<24><4> ) );
  DFFPOSX1 \mem_reg<24><3>  ( .D(n1244), .CLK(clk), .Q(\mem<24><3> ) );
  DFFPOSX1 \mem_reg<24><2>  ( .D(n1245), .CLK(clk), .Q(\mem<24><2> ) );
  DFFPOSX1 \mem_reg<24><1>  ( .D(n1246), .CLK(clk), .Q(\mem<24><1> ) );
  DFFPOSX1 \mem_reg<24><0>  ( .D(n1247), .CLK(clk), .Q(\mem<24><0> ) );
  DFFPOSX1 \mem_reg<25><7>  ( .D(n1248), .CLK(clk), .Q(\mem<25><7> ) );
  DFFPOSX1 \mem_reg<25><6>  ( .D(n1249), .CLK(clk), .Q(\mem<25><6> ) );
  DFFPOSX1 \mem_reg<25><5>  ( .D(n1250), .CLK(clk), .Q(\mem<25><5> ) );
  DFFPOSX1 \mem_reg<25><4>  ( .D(n1251), .CLK(clk), .Q(\mem<25><4> ) );
  DFFPOSX1 \mem_reg<25><3>  ( .D(n1252), .CLK(clk), .Q(\mem<25><3> ) );
  DFFPOSX1 \mem_reg<25><2>  ( .D(n1253), .CLK(clk), .Q(\mem<25><2> ) );
  DFFPOSX1 \mem_reg<25><1>  ( .D(n1254), .CLK(clk), .Q(\mem<25><1> ) );
  DFFPOSX1 \mem_reg<25><0>  ( .D(n1255), .CLK(clk), .Q(\mem<25><0> ) );
  DFFPOSX1 \mem_reg<26><7>  ( .D(n1256), .CLK(clk), .Q(\mem<26><7> ) );
  DFFPOSX1 \mem_reg<26><6>  ( .D(n1257), .CLK(clk), .Q(\mem<26><6> ) );
  DFFPOSX1 \mem_reg<26><5>  ( .D(n1258), .CLK(clk), .Q(\mem<26><5> ) );
  DFFPOSX1 \mem_reg<26><4>  ( .D(n1259), .CLK(clk), .Q(\mem<26><4> ) );
  DFFPOSX1 \mem_reg<26><3>  ( .D(n1260), .CLK(clk), .Q(\mem<26><3> ) );
  DFFPOSX1 \mem_reg<26><2>  ( .D(n1261), .CLK(clk), .Q(\mem<26><2> ) );
  DFFPOSX1 \mem_reg<26><1>  ( .D(n1262), .CLK(clk), .Q(\mem<26><1> ) );
  DFFPOSX1 \mem_reg<26><0>  ( .D(n1263), .CLK(clk), .Q(\mem<26><0> ) );
  DFFPOSX1 \mem_reg<27><7>  ( .D(n1264), .CLK(clk), .Q(\mem<27><7> ) );
  DFFPOSX1 \mem_reg<27><6>  ( .D(n1265), .CLK(clk), .Q(\mem<27><6> ) );
  DFFPOSX1 \mem_reg<27><5>  ( .D(n1266), .CLK(clk), .Q(\mem<27><5> ) );
  DFFPOSX1 \mem_reg<27><4>  ( .D(n1267), .CLK(clk), .Q(\mem<27><4> ) );
  DFFPOSX1 \mem_reg<27><3>  ( .D(n1268), .CLK(clk), .Q(\mem<27><3> ) );
  DFFPOSX1 \mem_reg<27><2>  ( .D(n1269), .CLK(clk), .Q(\mem<27><2> ) );
  DFFPOSX1 \mem_reg<27><1>  ( .D(n1270), .CLK(clk), .Q(\mem<27><1> ) );
  DFFPOSX1 \mem_reg<27><0>  ( .D(n1271), .CLK(clk), .Q(\mem<27><0> ) );
  DFFPOSX1 \mem_reg<28><7>  ( .D(n1272), .CLK(clk), .Q(\mem<28><7> ) );
  DFFPOSX1 \mem_reg<28><6>  ( .D(n1273), .CLK(clk), .Q(\mem<28><6> ) );
  DFFPOSX1 \mem_reg<28><5>  ( .D(n1274), .CLK(clk), .Q(\mem<28><5> ) );
  DFFPOSX1 \mem_reg<28><4>  ( .D(n1275), .CLK(clk), .Q(\mem<28><4> ) );
  DFFPOSX1 \mem_reg<28><3>  ( .D(n1276), .CLK(clk), .Q(\mem<28><3> ) );
  DFFPOSX1 \mem_reg<28><2>  ( .D(n1277), .CLK(clk), .Q(\mem<28><2> ) );
  DFFPOSX1 \mem_reg<28><1>  ( .D(n1278), .CLK(clk), .Q(\mem<28><1> ) );
  DFFPOSX1 \mem_reg<28><0>  ( .D(n1279), .CLK(clk), .Q(\mem<28><0> ) );
  DFFPOSX1 \mem_reg<29><7>  ( .D(n1280), .CLK(clk), .Q(\mem<29><7> ) );
  DFFPOSX1 \mem_reg<29><6>  ( .D(n1281), .CLK(clk), .Q(\mem<29><6> ) );
  DFFPOSX1 \mem_reg<29><5>  ( .D(n1282), .CLK(clk), .Q(\mem<29><5> ) );
  DFFPOSX1 \mem_reg<29><4>  ( .D(n1283), .CLK(clk), .Q(\mem<29><4> ) );
  DFFPOSX1 \mem_reg<29><3>  ( .D(n1284), .CLK(clk), .Q(\mem<29><3> ) );
  DFFPOSX1 \mem_reg<29><2>  ( .D(n1285), .CLK(clk), .Q(\mem<29><2> ) );
  DFFPOSX1 \mem_reg<29><1>  ( .D(n1286), .CLK(clk), .Q(\mem<29><1> ) );
  DFFPOSX1 \mem_reg<29><0>  ( .D(n1287), .CLK(clk), .Q(\mem<29><0> ) );
  DFFPOSX1 \mem_reg<30><7>  ( .D(n1288), .CLK(clk), .Q(\mem<30><7> ) );
  DFFPOSX1 \mem_reg<30><6>  ( .D(n1289), .CLK(clk), .Q(\mem<30><6> ) );
  DFFPOSX1 \mem_reg<30><5>  ( .D(n1290), .CLK(clk), .Q(\mem<30><5> ) );
  DFFPOSX1 \mem_reg<30><4>  ( .D(n1291), .CLK(clk), .Q(\mem<30><4> ) );
  DFFPOSX1 \mem_reg<30><3>  ( .D(n1292), .CLK(clk), .Q(\mem<30><3> ) );
  DFFPOSX1 \mem_reg<30><2>  ( .D(n1293), .CLK(clk), .Q(\mem<30><2> ) );
  DFFPOSX1 \mem_reg<30><1>  ( .D(n1294), .CLK(clk), .Q(\mem<30><1> ) );
  DFFPOSX1 \mem_reg<30><0>  ( .D(n1295), .CLK(clk), .Q(\mem<30><0> ) );
  DFFPOSX1 \mem_reg<31><7>  ( .D(n1296), .CLK(clk), .Q(\mem<31><7> ) );
  DFFPOSX1 \mem_reg<31><6>  ( .D(n1297), .CLK(clk), .Q(\mem<31><6> ) );
  DFFPOSX1 \mem_reg<31><5>  ( .D(n1298), .CLK(clk), .Q(\mem<31><5> ) );
  DFFPOSX1 \mem_reg<31><4>  ( .D(n1299), .CLK(clk), .Q(\mem<31><4> ) );
  DFFPOSX1 \mem_reg<31><3>  ( .D(n1300), .CLK(clk), .Q(\mem<31><3> ) );
  DFFPOSX1 \mem_reg<31><2>  ( .D(n1301), .CLK(clk), .Q(\mem<31><2> ) );
  DFFPOSX1 \mem_reg<31><1>  ( .D(n1302), .CLK(clk), .Q(\mem<31><1> ) );
  DFFPOSX1 \mem_reg<31><0>  ( .D(n1303), .CLK(clk), .Q(\mem<31><0> ) );
  DFFPOSX1 \mem_reg<32><7>  ( .D(n1304), .CLK(clk), .Q(\mem<32><7> ) );
  DFFPOSX1 \mem_reg<32><6>  ( .D(n1305), .CLK(clk), .Q(\mem<32><6> ) );
  DFFPOSX1 \mem_reg<32><5>  ( .D(n1306), .CLK(clk), .Q(\mem<32><5> ) );
  DFFPOSX1 \mem_reg<32><4>  ( .D(n1307), .CLK(clk), .Q(\mem<32><4> ) );
  DFFPOSX1 \mem_reg<32><3>  ( .D(n1308), .CLK(clk), .Q(\mem<32><3> ) );
  DFFPOSX1 \mem_reg<32><2>  ( .D(n1309), .CLK(clk), .Q(\mem<32><2> ) );
  DFFPOSX1 \mem_reg<32><1>  ( .D(n1310), .CLK(clk), .Q(\mem<32><1> ) );
  DFFPOSX1 \mem_reg<32><0>  ( .D(n1311), .CLK(clk), .Q(\mem<32><0> ) );
  AND2X2 U9 ( .A(n1479), .B(n1478), .Y(n1480) );
  AND2X2 U10 ( .A(n1474), .B(n1473), .Y(n1475) );
  AND2X2 U11 ( .A(n1468), .B(n1467), .Y(n1469) );
  AND2X2 U12 ( .A(n1463), .B(n1462), .Y(n1464) );
  AND2X2 U13 ( .A(n1457), .B(n1456), .Y(n1458) );
  AND2X2 U14 ( .A(n1452), .B(n1451), .Y(n1453) );
  AND2X2 U15 ( .A(n1446), .B(n1445), .Y(n1447) );
  AND2X2 U16 ( .A(n1441), .B(n1440), .Y(n1442) );
  AND2X2 U17 ( .A(n1435), .B(n1434), .Y(n1436) );
  AND2X2 U18 ( .A(n1430), .B(n1429), .Y(n1431) );
  AND2X2 U19 ( .A(n1424), .B(n1423), .Y(n1425) );
  AND2X2 U20 ( .A(n1419), .B(n1418), .Y(n1420) );
  AND2X2 U21 ( .A(n1413), .B(n1412), .Y(n1414) );
  AND2X2 U22 ( .A(n1408), .B(n1407), .Y(n1409) );
  AND2X2 U30 ( .A(n1328), .B(n1028), .Y(n1633) );
  AND2X2 U31 ( .A(n1327), .B(n1028), .Y(n1788) );
  AND2X2 U32 ( .A(n1328), .B(\addr_1c<0> ), .Y(n1653) );
  AND2X2 U33 ( .A(n1327), .B(\addr_1c<0> ), .Y(n1808) );
  AND2X2 U34 ( .A(n1322), .B(n1321), .Y(n1323) );
  AND2X2 U45 ( .A(n1315), .B(n1314), .Y(n1316) );
  NOR3X1 U94 ( .A(n1024), .B(rd), .C(n963), .Y(wr0) );
  NOR3X1 U95 ( .A(n1025), .B(wr), .C(n963), .Y(rd0) );
  OAI21X1 U96 ( .A(n1011), .B(n1040), .C(n1838), .Y(n1311) );
  NAND2X1 U97 ( .A(\mem<32><0> ), .B(n1011), .Y(n1838) );
  OAI21X1 U98 ( .A(n1011), .B(n1041), .C(n1837), .Y(n1310) );
  NAND2X1 U99 ( .A(\mem<32><1> ), .B(n1011), .Y(n1837) );
  OAI21X1 U100 ( .A(n1011), .B(n1042), .C(n1836), .Y(n1309) );
  NAND2X1 U101 ( .A(\mem<32><2> ), .B(n1011), .Y(n1836) );
  OAI21X1 U102 ( .A(n1011), .B(n1043), .C(n1835), .Y(n1308) );
  NAND2X1 U103 ( .A(\mem<32><3> ), .B(n1011), .Y(n1835) );
  OAI21X1 U104 ( .A(n1011), .B(n1044), .C(n1834), .Y(n1307) );
  NAND2X1 U105 ( .A(\mem<32><4> ), .B(n1011), .Y(n1834) );
  OAI21X1 U106 ( .A(n1011), .B(n1045), .C(n1833), .Y(n1306) );
  NAND2X1 U107 ( .A(\mem<32><5> ), .B(n1011), .Y(n1833) );
  OAI21X1 U108 ( .A(n1011), .B(n1046), .C(n1832), .Y(n1305) );
  NAND2X1 U109 ( .A(\mem<32><6> ), .B(n1011), .Y(n1832) );
  OAI21X1 U110 ( .A(n1011), .B(n1047), .C(n1831), .Y(n1304) );
  NAND2X1 U111 ( .A(\mem<32><7> ), .B(n1011), .Y(n1831) );
  NAND3X1 U112 ( .A(n1012), .B(n1829), .C(n965), .Y(n1839) );
  OAI21X1 U113 ( .A(n6), .B(n1032), .C(n1828), .Y(n1303) );
  NAND2X1 U114 ( .A(\mem<31><0> ), .B(n6), .Y(n1828) );
  OAI21X1 U115 ( .A(n6), .B(n1033), .C(n1827), .Y(n1302) );
  NAND2X1 U116 ( .A(\mem<31><1> ), .B(n6), .Y(n1827) );
  OAI21X1 U117 ( .A(n6), .B(n1034), .C(n1826), .Y(n1301) );
  NAND2X1 U118 ( .A(\mem<31><2> ), .B(n6), .Y(n1826) );
  OAI21X1 U119 ( .A(n6), .B(n1035), .C(n1825), .Y(n1300) );
  NAND2X1 U120 ( .A(\mem<31><3> ), .B(n6), .Y(n1825) );
  OAI21X1 U121 ( .A(n6), .B(n1036), .C(n1824), .Y(n1299) );
  NAND2X1 U122 ( .A(\mem<31><4> ), .B(n6), .Y(n1824) );
  OAI21X1 U123 ( .A(n6), .B(n1037), .C(n1823), .Y(n1298) );
  NAND2X1 U124 ( .A(\mem<31><5> ), .B(n6), .Y(n1823) );
  OAI21X1 U125 ( .A(n6), .B(n1038), .C(n1822), .Y(n1297) );
  NAND2X1 U126 ( .A(\mem<31><6> ), .B(n6), .Y(n1822) );
  OAI21X1 U127 ( .A(n6), .B(n1039), .C(n1821), .Y(n1296) );
  NAND2X1 U128 ( .A(\mem<31><7> ), .B(n6), .Y(n1821) );
  OAI21X1 U130 ( .A(n1040), .B(n1010), .C(n1817), .Y(n1295) );
  NAND2X1 U131 ( .A(\mem<30><0> ), .B(n1010), .Y(n1817) );
  OAI21X1 U132 ( .A(n1041), .B(n1009), .C(n1816), .Y(n1294) );
  NAND2X1 U133 ( .A(\mem<30><1> ), .B(n1010), .Y(n1816) );
  OAI21X1 U134 ( .A(n1042), .B(n1009), .C(n1815), .Y(n1293) );
  NAND2X1 U135 ( .A(\mem<30><2> ), .B(n1010), .Y(n1815) );
  OAI21X1 U136 ( .A(n1043), .B(n1009), .C(n1814), .Y(n1292) );
  NAND2X1 U137 ( .A(\mem<30><3> ), .B(n1010), .Y(n1814) );
  OAI21X1 U138 ( .A(n1044), .B(n1009), .C(n1813), .Y(n1291) );
  NAND2X1 U139 ( .A(\mem<30><4> ), .B(n1010), .Y(n1813) );
  OAI21X1 U140 ( .A(n1045), .B(n1009), .C(n1812), .Y(n1290) );
  NAND2X1 U141 ( .A(\mem<30><5> ), .B(n1010), .Y(n1812) );
  OAI21X1 U142 ( .A(n1046), .B(n1009), .C(n1811), .Y(n1289) );
  NAND2X1 U143 ( .A(\mem<30><6> ), .B(n1010), .Y(n1811) );
  OAI21X1 U144 ( .A(n1047), .B(n1009), .C(n1810), .Y(n1288) );
  NAND2X1 U145 ( .A(\mem<30><7> ), .B(n1010), .Y(n1810) );
  NAND3X1 U146 ( .A(n1809), .B(n1830), .C(n1808), .Y(n1818) );
  OAI21X1 U147 ( .A(n1032), .B(n1008), .C(n1806), .Y(n1287) );
  NAND2X1 U148 ( .A(\mem<29><0> ), .B(n1008), .Y(n1806) );
  OAI21X1 U149 ( .A(n1033), .B(n1008), .C(n1805), .Y(n1286) );
  NAND2X1 U150 ( .A(\mem<29><1> ), .B(n1008), .Y(n1805) );
  OAI21X1 U151 ( .A(n1034), .B(n1008), .C(n1804), .Y(n1285) );
  NAND2X1 U152 ( .A(\mem<29><2> ), .B(n1008), .Y(n1804) );
  OAI21X1 U153 ( .A(n1035), .B(n1008), .C(n1803), .Y(n1284) );
  NAND2X1 U154 ( .A(\mem<29><3> ), .B(n1008), .Y(n1803) );
  OAI21X1 U155 ( .A(n1036), .B(n1008), .C(n1802), .Y(n1283) );
  NAND2X1 U156 ( .A(\mem<29><4> ), .B(n1008), .Y(n1802) );
  OAI21X1 U157 ( .A(n1037), .B(n1008), .C(n1801), .Y(n1282) );
  NAND2X1 U158 ( .A(\mem<29><5> ), .B(n1008), .Y(n1801) );
  OAI21X1 U159 ( .A(n1038), .B(n1008), .C(n1800), .Y(n1281) );
  NAND2X1 U160 ( .A(\mem<29><6> ), .B(n1008), .Y(n1800) );
  OAI21X1 U161 ( .A(n1039), .B(n1008), .C(n1799), .Y(n1280) );
  NAND2X1 U162 ( .A(\mem<29><7> ), .B(n1008), .Y(n1799) );
  NAND3X1 U163 ( .A(n973), .B(n1013), .C(n1798), .Y(n1807) );
  OAI21X1 U164 ( .A(n1040), .B(n1007), .C(n1796), .Y(n1279) );
  NAND2X1 U165 ( .A(\mem<28><0> ), .B(n1007), .Y(n1796) );
  OAI21X1 U166 ( .A(n1041), .B(n1006), .C(n1795), .Y(n1278) );
  NAND2X1 U167 ( .A(\mem<28><1> ), .B(n1007), .Y(n1795) );
  OAI21X1 U168 ( .A(n1042), .B(n1006), .C(n1794), .Y(n1277) );
  NAND2X1 U169 ( .A(\mem<28><2> ), .B(n1007), .Y(n1794) );
  OAI21X1 U170 ( .A(n1043), .B(n1006), .C(n1793), .Y(n1276) );
  NAND2X1 U171 ( .A(\mem<28><3> ), .B(n1007), .Y(n1793) );
  OAI21X1 U172 ( .A(n1044), .B(n1006), .C(n1792), .Y(n1275) );
  NAND2X1 U173 ( .A(\mem<28><4> ), .B(n1007), .Y(n1792) );
  OAI21X1 U174 ( .A(n1045), .B(n1006), .C(n1791), .Y(n1274) );
  NAND2X1 U175 ( .A(\mem<28><5> ), .B(n1007), .Y(n1791) );
  OAI21X1 U176 ( .A(n1046), .B(n1006), .C(n1790), .Y(n1273) );
  NAND2X1 U177 ( .A(\mem<28><6> ), .B(n1007), .Y(n1790) );
  OAI21X1 U178 ( .A(n1047), .B(n1006), .C(n1789), .Y(n1272) );
  NAND2X1 U179 ( .A(\mem<28><7> ), .B(n1007), .Y(n1789) );
  NAND3X1 U180 ( .A(n1809), .B(n1830), .C(n1788), .Y(n1797) );
  OAI21X1 U181 ( .A(n1032), .B(n1005), .C(n1786), .Y(n1271) );
  NAND2X1 U182 ( .A(\mem<27><0> ), .B(n1005), .Y(n1786) );
  OAI21X1 U183 ( .A(n1033), .B(n1005), .C(n1785), .Y(n1270) );
  NAND2X1 U184 ( .A(\mem<27><1> ), .B(n1005), .Y(n1785) );
  OAI21X1 U185 ( .A(n1034), .B(n1005), .C(n1784), .Y(n1269) );
  NAND2X1 U186 ( .A(\mem<27><2> ), .B(n1005), .Y(n1784) );
  OAI21X1 U187 ( .A(n1035), .B(n1005), .C(n1783), .Y(n1268) );
  NAND2X1 U188 ( .A(\mem<27><3> ), .B(n1005), .Y(n1783) );
  OAI21X1 U189 ( .A(n1036), .B(n1005), .C(n1782), .Y(n1267) );
  NAND2X1 U190 ( .A(\mem<27><4> ), .B(n1005), .Y(n1782) );
  OAI21X1 U191 ( .A(n1037), .B(n1005), .C(n1781), .Y(n1266) );
  NAND2X1 U192 ( .A(\mem<27><5> ), .B(n1005), .Y(n1781) );
  OAI21X1 U193 ( .A(n1038), .B(n1005), .C(n1780), .Y(n1265) );
  NAND2X1 U194 ( .A(\mem<27><6> ), .B(n1005), .Y(n1780) );
  OAI21X1 U195 ( .A(n1039), .B(n1005), .C(n1779), .Y(n1264) );
  NAND2X1 U196 ( .A(\mem<27><7> ), .B(n1005), .Y(n1779) );
  NAND3X1 U197 ( .A(n973), .B(n1012), .C(n1778), .Y(n1787) );
  OAI21X1 U198 ( .A(n1040), .B(n1004), .C(n1776), .Y(n1263) );
  NAND2X1 U199 ( .A(\mem<26><0> ), .B(n1004), .Y(n1776) );
  OAI21X1 U200 ( .A(n1041), .B(n1003), .C(n1775), .Y(n1262) );
  NAND2X1 U201 ( .A(\mem<26><1> ), .B(n1004), .Y(n1775) );
  OAI21X1 U202 ( .A(n1042), .B(n1003), .C(n1774), .Y(n1261) );
  NAND2X1 U203 ( .A(\mem<26><2> ), .B(n1004), .Y(n1774) );
  OAI21X1 U204 ( .A(n1043), .B(n1003), .C(n1773), .Y(n1260) );
  NAND2X1 U205 ( .A(\mem<26><3> ), .B(n1004), .Y(n1773) );
  OAI21X1 U206 ( .A(n1044), .B(n1003), .C(n1772), .Y(n1259) );
  NAND2X1 U207 ( .A(\mem<26><4> ), .B(n1004), .Y(n1772) );
  OAI21X1 U208 ( .A(n1045), .B(n1003), .C(n1771), .Y(n1258) );
  NAND2X1 U209 ( .A(\mem<26><5> ), .B(n1004), .Y(n1771) );
  OAI21X1 U210 ( .A(n1046), .B(n1003), .C(n1770), .Y(n1257) );
  NAND2X1 U211 ( .A(\mem<26><6> ), .B(n1004), .Y(n1770) );
  OAI21X1 U212 ( .A(n1047), .B(n1003), .C(n1769), .Y(n1256) );
  NAND2X1 U213 ( .A(\mem<26><7> ), .B(n1004), .Y(n1769) );
  NAND3X1 U214 ( .A(n1808), .B(n1013), .C(n1768), .Y(n1777) );
  OAI21X1 U215 ( .A(n1032), .B(n1002), .C(n1766), .Y(n1255) );
  NAND2X1 U216 ( .A(\mem<25><0> ), .B(n1002), .Y(n1766) );
  OAI21X1 U217 ( .A(n1033), .B(n1002), .C(n1765), .Y(n1254) );
  NAND2X1 U218 ( .A(\mem<25><1> ), .B(n1002), .Y(n1765) );
  OAI21X1 U219 ( .A(n1034), .B(n1002), .C(n1764), .Y(n1253) );
  NAND2X1 U220 ( .A(\mem<25><2> ), .B(n1002), .Y(n1764) );
  OAI21X1 U221 ( .A(n1035), .B(n1002), .C(n1763), .Y(n1252) );
  NAND2X1 U222 ( .A(\mem<25><3> ), .B(n1002), .Y(n1763) );
  OAI21X1 U223 ( .A(n1036), .B(n1002), .C(n1762), .Y(n1251) );
  NAND2X1 U224 ( .A(\mem<25><4> ), .B(n1002), .Y(n1762) );
  OAI21X1 U225 ( .A(n1037), .B(n1002), .C(n1761), .Y(n1250) );
  NAND2X1 U226 ( .A(\mem<25><5> ), .B(n1002), .Y(n1761) );
  OAI21X1 U227 ( .A(n1038), .B(n1002), .C(n1760), .Y(n1249) );
  NAND2X1 U228 ( .A(\mem<25><6> ), .B(n1002), .Y(n1760) );
  OAI21X1 U229 ( .A(n1039), .B(n1002), .C(n1759), .Y(n1248) );
  NAND2X1 U230 ( .A(\mem<25><7> ), .B(n1002), .Y(n1759) );
  NAND3X1 U231 ( .A(n973), .B(n1013), .C(n1758), .Y(n1767) );
  OAI21X1 U232 ( .A(n1040), .B(n1001), .C(n1756), .Y(n1247) );
  NAND2X1 U233 ( .A(\mem<24><0> ), .B(n1001), .Y(n1756) );
  OAI21X1 U234 ( .A(n1041), .B(n1000), .C(n1755), .Y(n1246) );
  NAND2X1 U235 ( .A(\mem<24><1> ), .B(n1001), .Y(n1755) );
  OAI21X1 U236 ( .A(n1042), .B(n1000), .C(n1754), .Y(n1245) );
  NAND2X1 U237 ( .A(\mem<24><2> ), .B(n1001), .Y(n1754) );
  OAI21X1 U238 ( .A(n1043), .B(n1000), .C(n1753), .Y(n1244) );
  NAND2X1 U239 ( .A(\mem<24><3> ), .B(n1001), .Y(n1753) );
  OAI21X1 U240 ( .A(n1044), .B(n1000), .C(n1752), .Y(n1243) );
  NAND2X1 U241 ( .A(\mem<24><4> ), .B(n1001), .Y(n1752) );
  OAI21X1 U242 ( .A(n1045), .B(n1000), .C(n1751), .Y(n1242) );
  NAND2X1 U243 ( .A(\mem<24><5> ), .B(n1001), .Y(n1751) );
  OAI21X1 U244 ( .A(n1046), .B(n1000), .C(n1750), .Y(n1241) );
  NAND2X1 U245 ( .A(\mem<24><6> ), .B(n1001), .Y(n1750) );
  OAI21X1 U246 ( .A(n1047), .B(n1000), .C(n1749), .Y(n1240) );
  NAND2X1 U247 ( .A(\mem<24><7> ), .B(n1001), .Y(n1749) );
  NAND3X1 U248 ( .A(n1788), .B(n1013), .C(n1768), .Y(n1757) );
  OAI21X1 U249 ( .A(n1032), .B(n999), .C(n1747), .Y(n1239) );
  NAND2X1 U250 ( .A(\mem<23><0> ), .B(n999), .Y(n1747) );
  OAI21X1 U251 ( .A(n1033), .B(n999), .C(n1746), .Y(n1238) );
  NAND2X1 U252 ( .A(\mem<23><1> ), .B(n999), .Y(n1746) );
  OAI21X1 U253 ( .A(n1034), .B(n999), .C(n1745), .Y(n1237) );
  NAND2X1 U254 ( .A(\mem<23><2> ), .B(n999), .Y(n1745) );
  OAI21X1 U255 ( .A(n1035), .B(n999), .C(n1744), .Y(n1236) );
  NAND2X1 U256 ( .A(\mem<23><3> ), .B(n999), .Y(n1744) );
  OAI21X1 U257 ( .A(n1036), .B(n999), .C(n1743), .Y(n1235) );
  NAND2X1 U258 ( .A(\mem<23><4> ), .B(n999), .Y(n1743) );
  OAI21X1 U259 ( .A(n1037), .B(n999), .C(n1742), .Y(n1234) );
  NAND2X1 U260 ( .A(\mem<23><5> ), .B(n999), .Y(n1742) );
  OAI21X1 U261 ( .A(n1038), .B(n999), .C(n1741), .Y(n1233) );
  NAND2X1 U262 ( .A(\mem<23><6> ), .B(n999), .Y(n1741) );
  OAI21X1 U263 ( .A(n1039), .B(n999), .C(n1740), .Y(n1232) );
  NAND2X1 U264 ( .A(\mem<23><7> ), .B(n999), .Y(n1740) );
  NAND3X1 U265 ( .A(n973), .B(n1013), .C(n1739), .Y(n1748) );
  OAI21X1 U266 ( .A(n1040), .B(n998), .C(n1737), .Y(n1231) );
  NAND2X1 U267 ( .A(\mem<22><0> ), .B(n998), .Y(n1737) );
  OAI21X1 U268 ( .A(n1041), .B(n998), .C(n1736), .Y(n1230) );
  NAND2X1 U269 ( .A(\mem<22><1> ), .B(n998), .Y(n1736) );
  OAI21X1 U270 ( .A(n1042), .B(n998), .C(n1735), .Y(n1229) );
  NAND2X1 U271 ( .A(\mem<22><2> ), .B(n998), .Y(n1735) );
  OAI21X1 U272 ( .A(n1043), .B(n998), .C(n1734), .Y(n1228) );
  NAND2X1 U273 ( .A(\mem<22><3> ), .B(n998), .Y(n1734) );
  OAI21X1 U274 ( .A(n1044), .B(n998), .C(n1733), .Y(n1227) );
  NAND2X1 U275 ( .A(\mem<22><4> ), .B(n998), .Y(n1733) );
  OAI21X1 U276 ( .A(n1045), .B(n998), .C(n1732), .Y(n1226) );
  NAND2X1 U277 ( .A(\mem<22><5> ), .B(n998), .Y(n1732) );
  OAI21X1 U278 ( .A(n1046), .B(n998), .C(n1731), .Y(n1225) );
  NAND2X1 U279 ( .A(\mem<22><6> ), .B(n998), .Y(n1731) );
  OAI21X1 U280 ( .A(n1047), .B(n998), .C(n1730), .Y(n1224) );
  NAND2X1 U281 ( .A(\mem<22><7> ), .B(n998), .Y(n1730) );
  NAND3X1 U282 ( .A(n1808), .B(n1013), .C(n969), .Y(n1738) );
  OAI21X1 U283 ( .A(n1032), .B(n997), .C(n1728), .Y(n1223) );
  NAND2X1 U284 ( .A(\mem<21><0> ), .B(n997), .Y(n1728) );
  OAI21X1 U285 ( .A(n1033), .B(n997), .C(n1727), .Y(n1222) );
  NAND2X1 U286 ( .A(\mem<21><1> ), .B(n997), .Y(n1727) );
  OAI21X1 U287 ( .A(n1034), .B(n997), .C(n1726), .Y(n1221) );
  NAND2X1 U288 ( .A(\mem<21><2> ), .B(n997), .Y(n1726) );
  OAI21X1 U289 ( .A(n1035), .B(n997), .C(n1725), .Y(n1220) );
  NAND2X1 U290 ( .A(\mem<21><3> ), .B(n997), .Y(n1725) );
  OAI21X1 U291 ( .A(n1036), .B(n997), .C(n1724), .Y(n1219) );
  NAND2X1 U292 ( .A(\mem<21><4> ), .B(n997), .Y(n1724) );
  OAI21X1 U293 ( .A(n1037), .B(n997), .C(n1723), .Y(n1218) );
  NAND2X1 U294 ( .A(\mem<21><5> ), .B(n997), .Y(n1723) );
  OAI21X1 U295 ( .A(n1038), .B(n997), .C(n1722), .Y(n1217) );
  NAND2X1 U296 ( .A(\mem<21><6> ), .B(n997), .Y(n1722) );
  OAI21X1 U297 ( .A(n1039), .B(n997), .C(n1721), .Y(n1216) );
  NAND2X1 U298 ( .A(\mem<21><7> ), .B(n997), .Y(n1721) );
  NAND3X1 U299 ( .A(n973), .B(n1013), .C(n1720), .Y(n1729) );
  OAI21X1 U300 ( .A(n1040), .B(n996), .C(n1718), .Y(n1215) );
  NAND2X1 U301 ( .A(\mem<20><0> ), .B(n996), .Y(n1718) );
  OAI21X1 U302 ( .A(n1041), .B(n996), .C(n1717), .Y(n1214) );
  NAND2X1 U303 ( .A(\mem<20><1> ), .B(n996), .Y(n1717) );
  OAI21X1 U304 ( .A(n1042), .B(n996), .C(n1716), .Y(n1213) );
  NAND2X1 U305 ( .A(\mem<20><2> ), .B(n996), .Y(n1716) );
  OAI21X1 U306 ( .A(n1043), .B(n996), .C(n1715), .Y(n1212) );
  NAND2X1 U307 ( .A(\mem<20><3> ), .B(n996), .Y(n1715) );
  OAI21X1 U308 ( .A(n1044), .B(n996), .C(n1714), .Y(n1211) );
  NAND2X1 U309 ( .A(\mem<20><4> ), .B(n996), .Y(n1714) );
  OAI21X1 U310 ( .A(n1045), .B(n996), .C(n1713), .Y(n1210) );
  NAND2X1 U311 ( .A(\mem<20><5> ), .B(n996), .Y(n1713) );
  OAI21X1 U312 ( .A(n1046), .B(n996), .C(n1712), .Y(n1209) );
  NAND2X1 U313 ( .A(\mem<20><6> ), .B(n996), .Y(n1712) );
  OAI21X1 U314 ( .A(n1047), .B(n996), .C(n1711), .Y(n1208) );
  NAND2X1 U315 ( .A(\mem<20><7> ), .B(n996), .Y(n1711) );
  NAND3X1 U316 ( .A(n1788), .B(n1013), .C(n969), .Y(n1719) );
  OAI21X1 U317 ( .A(n1032), .B(n995), .C(n1709), .Y(n1207) );
  NAND2X1 U318 ( .A(\mem<19><0> ), .B(n995), .Y(n1709) );
  OAI21X1 U319 ( .A(n1033), .B(n995), .C(n1708), .Y(n1206) );
  NAND2X1 U320 ( .A(\mem<19><1> ), .B(n995), .Y(n1708) );
  OAI21X1 U321 ( .A(n1034), .B(n995), .C(n1707), .Y(n1205) );
  NAND2X1 U322 ( .A(\mem<19><2> ), .B(n995), .Y(n1707) );
  OAI21X1 U323 ( .A(n1035), .B(n995), .C(n1706), .Y(n1204) );
  NAND2X1 U324 ( .A(\mem<19><3> ), .B(n995), .Y(n1706) );
  OAI21X1 U325 ( .A(n1036), .B(n995), .C(n1705), .Y(n1203) );
  NAND2X1 U326 ( .A(\mem<19><4> ), .B(n995), .Y(n1705) );
  OAI21X1 U327 ( .A(n1037), .B(n995), .C(n1704), .Y(n1202) );
  NAND2X1 U328 ( .A(\mem<19><5> ), .B(n995), .Y(n1704) );
  OAI21X1 U329 ( .A(n1038), .B(n995), .C(n1703), .Y(n1201) );
  NAND2X1 U330 ( .A(\mem<19><6> ), .B(n995), .Y(n1703) );
  OAI21X1 U331 ( .A(n1039), .B(n995), .C(n1702), .Y(n1200) );
  NAND2X1 U332 ( .A(\mem<19><7> ), .B(n995), .Y(n1702) );
  NAND3X1 U333 ( .A(n973), .B(n1013), .C(n1701), .Y(n1710) );
  OAI21X1 U334 ( .A(n1040), .B(n994), .C(n1699), .Y(n1199) );
  NAND2X1 U335 ( .A(\mem<18><0> ), .B(n994), .Y(n1699) );
  OAI21X1 U336 ( .A(n1041), .B(n994), .C(n1698), .Y(n1198) );
  NAND2X1 U337 ( .A(\mem<18><1> ), .B(n994), .Y(n1698) );
  OAI21X1 U338 ( .A(n1042), .B(n994), .C(n1697), .Y(n1197) );
  NAND2X1 U339 ( .A(\mem<18><2> ), .B(n994), .Y(n1697) );
  OAI21X1 U340 ( .A(n1043), .B(n994), .C(n1696), .Y(n1196) );
  NAND2X1 U341 ( .A(\mem<18><3> ), .B(n994), .Y(n1696) );
  OAI21X1 U342 ( .A(n1044), .B(n994), .C(n1695), .Y(n1195) );
  NAND2X1 U343 ( .A(\mem<18><4> ), .B(n994), .Y(n1695) );
  OAI21X1 U344 ( .A(n1045), .B(n994), .C(n1694), .Y(n1194) );
  NAND2X1 U345 ( .A(\mem<18><5> ), .B(n994), .Y(n1694) );
  OAI21X1 U346 ( .A(n1046), .B(n994), .C(n1693), .Y(n1193) );
  NAND2X1 U347 ( .A(\mem<18><6> ), .B(n994), .Y(n1693) );
  OAI21X1 U348 ( .A(n1047), .B(n994), .C(n1692), .Y(n1192) );
  NAND2X1 U349 ( .A(\mem<18><7> ), .B(n994), .Y(n1692) );
  NAND3X1 U350 ( .A(n1808), .B(n1013), .C(n967), .Y(n1700) );
  OAI21X1 U351 ( .A(n1032), .B(n993), .C(n1690), .Y(n1191) );
  NAND2X1 U352 ( .A(\mem<17><0> ), .B(n993), .Y(n1690) );
  OAI21X1 U353 ( .A(n1033), .B(n993), .C(n1689), .Y(n1190) );
  NAND2X1 U354 ( .A(\mem<17><1> ), .B(n993), .Y(n1689) );
  OAI21X1 U355 ( .A(n1034), .B(n993), .C(n1688), .Y(n1189) );
  NAND2X1 U356 ( .A(\mem<17><2> ), .B(n993), .Y(n1688) );
  OAI21X1 U357 ( .A(n1035), .B(n993), .C(n1687), .Y(n1188) );
  NAND2X1 U358 ( .A(\mem<17><3> ), .B(n993), .Y(n1687) );
  OAI21X1 U359 ( .A(n1036), .B(n993), .C(n1686), .Y(n1187) );
  NAND2X1 U360 ( .A(\mem<17><4> ), .B(n993), .Y(n1686) );
  OAI21X1 U361 ( .A(n1037), .B(n993), .C(n1685), .Y(n1186) );
  NAND2X1 U362 ( .A(\mem<17><5> ), .B(n993), .Y(n1685) );
  OAI21X1 U363 ( .A(n1038), .B(n993), .C(n1684), .Y(n1185) );
  NAND2X1 U364 ( .A(\mem<17><6> ), .B(n993), .Y(n1684) );
  OAI21X1 U365 ( .A(n1039), .B(n993), .C(n1683), .Y(n1184) );
  NAND2X1 U366 ( .A(\mem<17><7> ), .B(n993), .Y(n1683) );
  NAND3X1 U367 ( .A(n973), .B(n1013), .C(n1682), .Y(n1691) );
  OAI21X1 U368 ( .A(n1040), .B(n992), .C(n1680), .Y(n1183) );
  NAND2X1 U369 ( .A(\mem<16><0> ), .B(n992), .Y(n1680) );
  OAI21X1 U370 ( .A(n1041), .B(n992), .C(n1679), .Y(n1182) );
  NAND2X1 U371 ( .A(\mem<16><1> ), .B(n992), .Y(n1679) );
  OAI21X1 U372 ( .A(n1042), .B(n992), .C(n1678), .Y(n1181) );
  NAND2X1 U373 ( .A(\mem<16><2> ), .B(n992), .Y(n1678) );
  OAI21X1 U374 ( .A(n1043), .B(n992), .C(n1677), .Y(n1180) );
  NAND2X1 U375 ( .A(\mem<16><3> ), .B(n992), .Y(n1677) );
  OAI21X1 U376 ( .A(n1044), .B(n992), .C(n1676), .Y(n1179) );
  NAND2X1 U377 ( .A(\mem<16><4> ), .B(n992), .Y(n1676) );
  OAI21X1 U378 ( .A(n1045), .B(n992), .C(n1675), .Y(n1178) );
  NAND2X1 U379 ( .A(\mem<16><5> ), .B(n992), .Y(n1675) );
  OAI21X1 U380 ( .A(n1046), .B(n992), .C(n1674), .Y(n1177) );
  NAND2X1 U381 ( .A(\mem<16><6> ), .B(n992), .Y(n1674) );
  OAI21X1 U382 ( .A(n1047), .B(n992), .C(n1673), .Y(n1176) );
  NAND2X1 U383 ( .A(\mem<16><7> ), .B(n992), .Y(n1673) );
  NAND3X1 U384 ( .A(n1788), .B(n1013), .C(n967), .Y(n1681) );
  OAI21X1 U385 ( .A(n1032), .B(n991), .C(n1671), .Y(n1175) );
  NAND2X1 U386 ( .A(\mem<15><0> ), .B(n991), .Y(n1671) );
  OAI21X1 U387 ( .A(n1033), .B(n991), .C(n1670), .Y(n1174) );
  NAND2X1 U388 ( .A(\mem<15><1> ), .B(n991), .Y(n1670) );
  OAI21X1 U389 ( .A(n1034), .B(n991), .C(n1669), .Y(n1173) );
  NAND2X1 U390 ( .A(\mem<15><2> ), .B(n991), .Y(n1669) );
  OAI21X1 U391 ( .A(n1035), .B(n991), .C(n1668), .Y(n1172) );
  NAND2X1 U392 ( .A(\mem<15><3> ), .B(n991), .Y(n1668) );
  OAI21X1 U393 ( .A(n1036), .B(n991), .C(n1667), .Y(n1171) );
  NAND2X1 U394 ( .A(\mem<15><4> ), .B(n991), .Y(n1667) );
  OAI21X1 U395 ( .A(n1037), .B(n991), .C(n1666), .Y(n1170) );
  NAND2X1 U396 ( .A(\mem<15><5> ), .B(n991), .Y(n1666) );
  OAI21X1 U397 ( .A(n1038), .B(n991), .C(n1665), .Y(n1169) );
  NAND2X1 U398 ( .A(\mem<15><6> ), .B(n991), .Y(n1665) );
  OAI21X1 U399 ( .A(n1039), .B(n991), .C(n1664), .Y(n1168) );
  NAND2X1 U400 ( .A(\mem<15><7> ), .B(n991), .Y(n1664) );
  NAND3X1 U401 ( .A(n973), .B(n1013), .C(n1663), .Y(n1672) );
  OAI21X1 U402 ( .A(n1040), .B(n990), .C(n1661), .Y(n1167) );
  NAND2X1 U403 ( .A(\mem<14><0> ), .B(n990), .Y(n1661) );
  OAI21X1 U404 ( .A(n1041), .B(n989), .C(n1660), .Y(n1166) );
  NAND2X1 U405 ( .A(\mem<14><1> ), .B(n990), .Y(n1660) );
  OAI21X1 U406 ( .A(n1042), .B(n989), .C(n1659), .Y(n1165) );
  NAND2X1 U407 ( .A(\mem<14><2> ), .B(n990), .Y(n1659) );
  OAI21X1 U408 ( .A(n1043), .B(n989), .C(n1658), .Y(n1164) );
  NAND2X1 U409 ( .A(\mem<14><3> ), .B(n990), .Y(n1658) );
  OAI21X1 U410 ( .A(n1044), .B(n989), .C(n1657), .Y(n1163) );
  NAND2X1 U411 ( .A(\mem<14><4> ), .B(n990), .Y(n1657) );
  OAI21X1 U412 ( .A(n1045), .B(n989), .C(n1656), .Y(n1162) );
  NAND2X1 U413 ( .A(\mem<14><5> ), .B(n990), .Y(n1656) );
  OAI21X1 U414 ( .A(n1046), .B(n989), .C(n1655), .Y(n1161) );
  NAND2X1 U415 ( .A(\mem<14><6> ), .B(n990), .Y(n1655) );
  OAI21X1 U416 ( .A(n1047), .B(n989), .C(n1654), .Y(n1160) );
  NAND2X1 U417 ( .A(\mem<14><7> ), .B(n990), .Y(n1654) );
  NAND3X1 U418 ( .A(n1809), .B(n1012), .C(n1653), .Y(n1662) );
  OAI21X1 U419 ( .A(n1032), .B(n988), .C(n1651), .Y(n1159) );
  NAND2X1 U420 ( .A(\mem<13><0> ), .B(n988), .Y(n1651) );
  OAI21X1 U421 ( .A(n1033), .B(n988), .C(n1650), .Y(n1158) );
  NAND2X1 U422 ( .A(\mem<13><1> ), .B(n988), .Y(n1650) );
  OAI21X1 U423 ( .A(n1034), .B(n988), .C(n1649), .Y(n1157) );
  NAND2X1 U424 ( .A(\mem<13><2> ), .B(n988), .Y(n1649) );
  OAI21X1 U425 ( .A(n1035), .B(n988), .C(n1648), .Y(n1156) );
  NAND2X1 U426 ( .A(\mem<13><3> ), .B(n988), .Y(n1648) );
  OAI21X1 U427 ( .A(n1036), .B(n988), .C(n1647), .Y(n1155) );
  NAND2X1 U428 ( .A(\mem<13><4> ), .B(n988), .Y(n1647) );
  OAI21X1 U429 ( .A(n1037), .B(n988), .C(n1646), .Y(n1154) );
  NAND2X1 U430 ( .A(\mem<13><5> ), .B(n988), .Y(n1646) );
  OAI21X1 U431 ( .A(n1038), .B(n988), .C(n1645), .Y(n1153) );
  NAND2X1 U432 ( .A(\mem<13><6> ), .B(n988), .Y(n1645) );
  OAI21X1 U433 ( .A(n1039), .B(n988), .C(n1644), .Y(n1152) );
  NAND2X1 U434 ( .A(\mem<13><7> ), .B(n988), .Y(n1644) );
  NAND3X1 U435 ( .A(n973), .B(n1012), .C(n1643), .Y(n1652) );
  OAI21X1 U436 ( .A(n1040), .B(n987), .C(n1641), .Y(n1151) );
  NAND2X1 U437 ( .A(\mem<12><0> ), .B(n987), .Y(n1641) );
  OAI21X1 U438 ( .A(n1041), .B(n986), .C(n1640), .Y(n1150) );
  NAND2X1 U439 ( .A(\mem<12><1> ), .B(n987), .Y(n1640) );
  OAI21X1 U440 ( .A(n1042), .B(n986), .C(n1639), .Y(n1149) );
  NAND2X1 U441 ( .A(\mem<12><2> ), .B(n987), .Y(n1639) );
  OAI21X1 U442 ( .A(n1043), .B(n986), .C(n1638), .Y(n1148) );
  NAND2X1 U443 ( .A(\mem<12><3> ), .B(n987), .Y(n1638) );
  OAI21X1 U444 ( .A(n1044), .B(n986), .C(n1637), .Y(n1147) );
  NAND2X1 U445 ( .A(\mem<12><4> ), .B(n987), .Y(n1637) );
  OAI21X1 U446 ( .A(n1045), .B(n986), .C(n1636), .Y(n1146) );
  NAND2X1 U447 ( .A(\mem<12><5> ), .B(n987), .Y(n1636) );
  OAI21X1 U448 ( .A(n1046), .B(n986), .C(n1635), .Y(n1145) );
  NAND2X1 U449 ( .A(\mem<12><6> ), .B(n987), .Y(n1635) );
  OAI21X1 U450 ( .A(n1047), .B(n986), .C(n1634), .Y(n1144) );
  NAND2X1 U451 ( .A(\mem<12><7> ), .B(n987), .Y(n1634) );
  NAND3X1 U452 ( .A(n1809), .B(n1012), .C(n1633), .Y(n1642) );
  OAI21X1 U453 ( .A(n1032), .B(n985), .C(n1630), .Y(n1143) );
  NAND2X1 U454 ( .A(\mem<11><0> ), .B(n985), .Y(n1630) );
  OAI21X1 U455 ( .A(n1033), .B(n985), .C(n1629), .Y(n1142) );
  NAND2X1 U456 ( .A(\mem<11><1> ), .B(n985), .Y(n1629) );
  OAI21X1 U457 ( .A(n1034), .B(n985), .C(n1628), .Y(n1141) );
  NAND2X1 U458 ( .A(\mem<11><2> ), .B(n985), .Y(n1628) );
  OAI21X1 U459 ( .A(n1035), .B(n985), .C(n1627), .Y(n1140) );
  NAND2X1 U460 ( .A(\mem<11><3> ), .B(n985), .Y(n1627) );
  OAI21X1 U461 ( .A(n1036), .B(n985), .C(n1626), .Y(n1139) );
  NAND2X1 U462 ( .A(\mem<11><4> ), .B(n985), .Y(n1626) );
  OAI21X1 U463 ( .A(n1037), .B(n985), .C(n1625), .Y(n1138) );
  NAND2X1 U464 ( .A(\mem<11><5> ), .B(n985), .Y(n1625) );
  OAI21X1 U465 ( .A(n1038), .B(n985), .C(n1624), .Y(n1137) );
  NAND2X1 U466 ( .A(\mem<11><6> ), .B(n985), .Y(n1624) );
  OAI21X1 U467 ( .A(n1039), .B(n985), .C(n1623), .Y(n1136) );
  NAND2X1 U468 ( .A(\mem<11><7> ), .B(n985), .Y(n1623) );
  NAND3X1 U469 ( .A(n973), .B(n1012), .C(n1622), .Y(n1631) );
  OAI21X1 U470 ( .A(n1040), .B(n984), .C(n1620), .Y(n1135) );
  NAND2X1 U471 ( .A(\mem<10><0> ), .B(n984), .Y(n1620) );
  OAI21X1 U472 ( .A(n1041), .B(n983), .C(n1619), .Y(n1134) );
  NAND2X1 U473 ( .A(\mem<10><1> ), .B(n984), .Y(n1619) );
  OAI21X1 U474 ( .A(n1042), .B(n983), .C(n1618), .Y(n1133) );
  NAND2X1 U475 ( .A(\mem<10><2> ), .B(n984), .Y(n1618) );
  OAI21X1 U476 ( .A(n1043), .B(n983), .C(n1617), .Y(n1132) );
  NAND2X1 U477 ( .A(\mem<10><3> ), .B(n984), .Y(n1617) );
  OAI21X1 U478 ( .A(n1044), .B(n983), .C(n1616), .Y(n1131) );
  NAND2X1 U479 ( .A(\mem<10><4> ), .B(n984), .Y(n1616) );
  OAI21X1 U480 ( .A(n1045), .B(n983), .C(n1615), .Y(n1130) );
  NAND2X1 U481 ( .A(\mem<10><5> ), .B(n984), .Y(n1615) );
  OAI21X1 U482 ( .A(n1046), .B(n983), .C(n1614), .Y(n1129) );
  NAND2X1 U483 ( .A(\mem<10><6> ), .B(n984), .Y(n1614) );
  OAI21X1 U484 ( .A(n1047), .B(n983), .C(n1613), .Y(n1128) );
  NAND2X1 U485 ( .A(\mem<10><7> ), .B(n984), .Y(n1613) );
  NAND3X1 U486 ( .A(n1768), .B(n1012), .C(n1653), .Y(n1621) );
  OAI21X1 U487 ( .A(n1032), .B(n982), .C(n1611), .Y(n1127) );
  NAND2X1 U488 ( .A(\mem<9><0> ), .B(n982), .Y(n1611) );
  OAI21X1 U489 ( .A(n1033), .B(n982), .C(n1610), .Y(n1126) );
  NAND2X1 U490 ( .A(\mem<9><1> ), .B(n982), .Y(n1610) );
  OAI21X1 U491 ( .A(n1034), .B(n982), .C(n1609), .Y(n1125) );
  NAND2X1 U492 ( .A(\mem<9><2> ), .B(n982), .Y(n1609) );
  OAI21X1 U493 ( .A(n1035), .B(n982), .C(n1608), .Y(n1124) );
  NAND2X1 U494 ( .A(\mem<9><3> ), .B(n982), .Y(n1608) );
  OAI21X1 U495 ( .A(n1036), .B(n982), .C(n1607), .Y(n1123) );
  NAND2X1 U496 ( .A(\mem<9><4> ), .B(n982), .Y(n1607) );
  OAI21X1 U497 ( .A(n1037), .B(n982), .C(n1606), .Y(n1122) );
  NAND2X1 U498 ( .A(\mem<9><5> ), .B(n982), .Y(n1606) );
  OAI21X1 U499 ( .A(n1038), .B(n982), .C(n1605), .Y(n1121) );
  NAND2X1 U500 ( .A(\mem<9><6> ), .B(n982), .Y(n1605) );
  OAI21X1 U501 ( .A(n1039), .B(n982), .C(n1604), .Y(n1120) );
  NAND2X1 U502 ( .A(\mem<9><7> ), .B(n982), .Y(n1604) );
  NAND3X1 U503 ( .A(n973), .B(n1012), .C(n1603), .Y(n1612) );
  OAI21X1 U504 ( .A(n1040), .B(n981), .C(n1601), .Y(n1119) );
  NAND2X1 U505 ( .A(\mem<8><0> ), .B(n981), .Y(n1601) );
  OAI21X1 U506 ( .A(n1041), .B(n980), .C(n1600), .Y(n1118) );
  NAND2X1 U507 ( .A(\mem<8><1> ), .B(n981), .Y(n1600) );
  OAI21X1 U508 ( .A(n1042), .B(n980), .C(n1599), .Y(n1117) );
  NAND2X1 U509 ( .A(\mem<8><2> ), .B(n981), .Y(n1599) );
  OAI21X1 U510 ( .A(n1043), .B(n980), .C(n1598), .Y(n1116) );
  NAND2X1 U511 ( .A(\mem<8><3> ), .B(n981), .Y(n1598) );
  OAI21X1 U512 ( .A(n1044), .B(n980), .C(n1597), .Y(n1115) );
  NAND2X1 U513 ( .A(\mem<8><4> ), .B(n981), .Y(n1597) );
  OAI21X1 U514 ( .A(n1045), .B(n980), .C(n1596), .Y(n1114) );
  NAND2X1 U515 ( .A(\mem<8><5> ), .B(n981), .Y(n1596) );
  OAI21X1 U516 ( .A(n1046), .B(n980), .C(n1595), .Y(n1113) );
  NAND2X1 U517 ( .A(\mem<8><6> ), .B(n981), .Y(n1595) );
  OAI21X1 U518 ( .A(n1047), .B(n980), .C(n1594), .Y(n1112) );
  NAND2X1 U519 ( .A(\mem<8><7> ), .B(n981), .Y(n1594) );
  NAND3X1 U520 ( .A(n1768), .B(n1012), .C(n1633), .Y(n1602) );
  OAI21X1 U521 ( .A(n1032), .B(n979), .C(n1591), .Y(n1111) );
  NAND2X1 U522 ( .A(\mem<7><0> ), .B(n979), .Y(n1591) );
  OAI21X1 U523 ( .A(n1033), .B(n979), .C(n1590), .Y(n1110) );
  NAND2X1 U524 ( .A(\mem<7><1> ), .B(n979), .Y(n1590) );
  OAI21X1 U525 ( .A(n1034), .B(n979), .C(n1589), .Y(n1109) );
  NAND2X1 U526 ( .A(\mem<7><2> ), .B(n979), .Y(n1589) );
  OAI21X1 U527 ( .A(n1035), .B(n979), .C(n1588), .Y(n1108) );
  NAND2X1 U528 ( .A(\mem<7><3> ), .B(n979), .Y(n1588) );
  OAI21X1 U529 ( .A(n1036), .B(n979), .C(n1587), .Y(n1107) );
  NAND2X1 U530 ( .A(\mem<7><4> ), .B(n979), .Y(n1587) );
  OAI21X1 U531 ( .A(n1037), .B(n979), .C(n1586), .Y(n1106) );
  NAND2X1 U532 ( .A(\mem<7><5> ), .B(n979), .Y(n1586) );
  OAI21X1 U533 ( .A(n1038), .B(n979), .C(n1585), .Y(n1105) );
  NAND2X1 U534 ( .A(\mem<7><6> ), .B(n979), .Y(n1585) );
  OAI21X1 U535 ( .A(n1039), .B(n979), .C(n1584), .Y(n1104) );
  NAND2X1 U536 ( .A(\mem<7><7> ), .B(n979), .Y(n1584) );
  NAND3X1 U537 ( .A(n973), .B(n1012), .C(n1583), .Y(n1592) );
  OAI21X1 U538 ( .A(n1040), .B(n978), .C(n1581), .Y(n1103) );
  NAND2X1 U539 ( .A(\mem<6><0> ), .B(n978), .Y(n1581) );
  OAI21X1 U540 ( .A(n1041), .B(n978), .C(n1580), .Y(n1102) );
  NAND2X1 U541 ( .A(\mem<6><1> ), .B(n978), .Y(n1580) );
  OAI21X1 U542 ( .A(n1042), .B(n978), .C(n1579), .Y(n1101) );
  NAND2X1 U543 ( .A(\mem<6><2> ), .B(n978), .Y(n1579) );
  OAI21X1 U544 ( .A(n1043), .B(n978), .C(n1578), .Y(n1100) );
  NAND2X1 U545 ( .A(\mem<6><3> ), .B(n978), .Y(n1578) );
  OAI21X1 U546 ( .A(n1044), .B(n978), .C(n1577), .Y(n1099) );
  NAND2X1 U547 ( .A(\mem<6><4> ), .B(n978), .Y(n1577) );
  OAI21X1 U548 ( .A(n1045), .B(n978), .C(n1576), .Y(n1098) );
  NAND2X1 U549 ( .A(\mem<6><5> ), .B(n978), .Y(n1576) );
  OAI21X1 U550 ( .A(n1046), .B(n978), .C(n1575), .Y(n1097) );
  NAND2X1 U551 ( .A(\mem<6><6> ), .B(n978), .Y(n1575) );
  OAI21X1 U552 ( .A(n1047), .B(n978), .C(n1574), .Y(n1096) );
  NAND2X1 U553 ( .A(\mem<6><7> ), .B(n978), .Y(n1574) );
  NAND3X1 U554 ( .A(n969), .B(n1012), .C(n1653), .Y(n1582) );
  OAI21X1 U555 ( .A(n1032), .B(n977), .C(n1572), .Y(n1095) );
  NAND2X1 U556 ( .A(\mem<5><0> ), .B(n977), .Y(n1572) );
  OAI21X1 U557 ( .A(n1033), .B(n977), .C(n1571), .Y(n1094) );
  NAND2X1 U558 ( .A(\mem<5><1> ), .B(n977), .Y(n1571) );
  OAI21X1 U559 ( .A(n1034), .B(n977), .C(n1570), .Y(n1093) );
  NAND2X1 U560 ( .A(\mem<5><2> ), .B(n977), .Y(n1570) );
  OAI21X1 U561 ( .A(n1035), .B(n977), .C(n1569), .Y(n1092) );
  NAND2X1 U562 ( .A(\mem<5><3> ), .B(n977), .Y(n1569) );
  OAI21X1 U563 ( .A(n1036), .B(n977), .C(n1568), .Y(n1091) );
  NAND2X1 U564 ( .A(\mem<5><4> ), .B(n977), .Y(n1568) );
  OAI21X1 U565 ( .A(n1037), .B(n977), .C(n1567), .Y(n1090) );
  NAND2X1 U566 ( .A(\mem<5><5> ), .B(n977), .Y(n1567) );
  OAI21X1 U567 ( .A(n1038), .B(n977), .C(n1566), .Y(n1089) );
  NAND2X1 U568 ( .A(\mem<5><6> ), .B(n977), .Y(n1566) );
  OAI21X1 U569 ( .A(n1039), .B(n977), .C(n1565), .Y(n1088) );
  NAND2X1 U570 ( .A(\mem<5><7> ), .B(n977), .Y(n1565) );
  NAND3X1 U571 ( .A(n973), .B(n1012), .C(n1564), .Y(n1573) );
  OAI21X1 U572 ( .A(n1040), .B(n976), .C(n1562), .Y(n1087) );
  NAND2X1 U573 ( .A(\mem<4><0> ), .B(n976), .Y(n1562) );
  OAI21X1 U574 ( .A(n1041), .B(n976), .C(n1561), .Y(n1086) );
  NAND2X1 U575 ( .A(\mem<4><1> ), .B(n976), .Y(n1561) );
  OAI21X1 U576 ( .A(n1042), .B(n976), .C(n1560), .Y(n1085) );
  NAND2X1 U577 ( .A(\mem<4><2> ), .B(n976), .Y(n1560) );
  OAI21X1 U578 ( .A(n1043), .B(n976), .C(n1559), .Y(n1084) );
  NAND2X1 U579 ( .A(\mem<4><3> ), .B(n976), .Y(n1559) );
  OAI21X1 U580 ( .A(n1044), .B(n976), .C(n1558), .Y(n1083) );
  NAND2X1 U581 ( .A(\mem<4><4> ), .B(n976), .Y(n1558) );
  OAI21X1 U582 ( .A(n1045), .B(n976), .C(n1557), .Y(n1082) );
  NAND2X1 U583 ( .A(\mem<4><5> ), .B(n976), .Y(n1557) );
  OAI21X1 U584 ( .A(n1046), .B(n976), .C(n1556), .Y(n1081) );
  NAND2X1 U585 ( .A(\mem<4><6> ), .B(n976), .Y(n1556) );
  OAI21X1 U586 ( .A(n1047), .B(n976), .C(n1555), .Y(n1080) );
  NAND2X1 U587 ( .A(\mem<4><7> ), .B(n976), .Y(n1555) );
  NAND3X1 U588 ( .A(n969), .B(n1012), .C(n1633), .Y(n1563) );
  OAI21X1 U590 ( .A(n1032), .B(n975), .C(n1552), .Y(n1079) );
  NAND2X1 U591 ( .A(\mem<3><0> ), .B(n975), .Y(n1552) );
  OAI21X1 U592 ( .A(n1033), .B(n975), .C(n1551), .Y(n1078) );
  NAND2X1 U593 ( .A(\mem<3><1> ), .B(n975), .Y(n1551) );
  OAI21X1 U594 ( .A(n1034), .B(n975), .C(n1550), .Y(n1077) );
  NAND2X1 U595 ( .A(\mem<3><2> ), .B(n975), .Y(n1550) );
  OAI21X1 U596 ( .A(n1035), .B(n975), .C(n1549), .Y(n1076) );
  NAND2X1 U597 ( .A(\mem<3><3> ), .B(n975), .Y(n1549) );
  OAI21X1 U598 ( .A(n1036), .B(n975), .C(n1548), .Y(n1075) );
  NAND2X1 U599 ( .A(\mem<3><4> ), .B(n975), .Y(n1548) );
  OAI21X1 U600 ( .A(n1037), .B(n975), .C(n1547), .Y(n1074) );
  NAND2X1 U601 ( .A(\mem<3><5> ), .B(n975), .Y(n1547) );
  OAI21X1 U602 ( .A(n1038), .B(n975), .C(n1546), .Y(n1073) );
  NAND2X1 U603 ( .A(\mem<3><6> ), .B(n975), .Y(n1546) );
  OAI21X1 U604 ( .A(n1039), .B(n975), .C(n1545), .Y(n1072) );
  NAND2X1 U605 ( .A(\mem<3><7> ), .B(n975), .Y(n1545) );
  NAND3X1 U606 ( .A(n973), .B(n1012), .C(n1544), .Y(n1553) );
  OAI21X1 U607 ( .A(n1040), .B(n974), .C(n1542), .Y(n1071) );
  NAND2X1 U608 ( .A(\mem<2><0> ), .B(n974), .Y(n1542) );
  OAI21X1 U609 ( .A(n1041), .B(n974), .C(n1541), .Y(n1070) );
  NAND2X1 U610 ( .A(\mem<2><1> ), .B(n974), .Y(n1541) );
  OAI21X1 U611 ( .A(n1042), .B(n974), .C(n1540), .Y(n1069) );
  NAND2X1 U612 ( .A(\mem<2><2> ), .B(n974), .Y(n1540) );
  OAI21X1 U613 ( .A(n1043), .B(n974), .C(n1539), .Y(n1068) );
  NAND2X1 U614 ( .A(\mem<2><3> ), .B(n974), .Y(n1539) );
  OAI21X1 U615 ( .A(n1044), .B(n974), .C(n1538), .Y(n1067) );
  NAND2X1 U616 ( .A(\mem<2><4> ), .B(n974), .Y(n1538) );
  OAI21X1 U617 ( .A(n1045), .B(n974), .C(n1537), .Y(n1066) );
  NAND2X1 U618 ( .A(\mem<2><5> ), .B(n974), .Y(n1537) );
  OAI21X1 U619 ( .A(n1046), .B(n974), .C(n1536), .Y(n1065) );
  NAND2X1 U620 ( .A(\mem<2><6> ), .B(n974), .Y(n1536) );
  OAI21X1 U621 ( .A(n1047), .B(n974), .C(n1535), .Y(n1064) );
  NAND2X1 U622 ( .A(\mem<2><7> ), .B(n974), .Y(n1535) );
  NAND3X1 U623 ( .A(n967), .B(n1012), .C(n1653), .Y(n1543) );
  OAI21X1 U624 ( .A(n1032), .B(n8), .C(n1534), .Y(n1063) );
  NAND2X1 U625 ( .A(\mem<1><0> ), .B(n8), .Y(n1534) );
  OAI21X1 U626 ( .A(n1033), .B(n8), .C(n1533), .Y(n1062) );
  NAND2X1 U627 ( .A(\mem<1><1> ), .B(n8), .Y(n1533) );
  OAI21X1 U628 ( .A(n1034), .B(n8), .C(n1532), .Y(n1061) );
  NAND2X1 U629 ( .A(\mem<1><2> ), .B(n8), .Y(n1532) );
  OAI21X1 U630 ( .A(n1035), .B(n8), .C(n1531), .Y(n1060) );
  NAND2X1 U631 ( .A(\mem<1><3> ), .B(n8), .Y(n1531) );
  OAI21X1 U632 ( .A(n1036), .B(n8), .C(n1530), .Y(n1059) );
  NAND2X1 U633 ( .A(\mem<1><4> ), .B(n8), .Y(n1530) );
  OAI21X1 U634 ( .A(n1037), .B(n8), .C(n1529), .Y(n1058) );
  NAND2X1 U635 ( .A(\mem<1><5> ), .B(n8), .Y(n1529) );
  OAI21X1 U636 ( .A(n1038), .B(n8), .C(n1528), .Y(n1057) );
  NAND2X1 U637 ( .A(\mem<1><6> ), .B(n8), .Y(n1528) );
  OAI21X1 U638 ( .A(n1039), .B(n8), .C(n1527), .Y(n1056) );
  NAND2X1 U639 ( .A(\mem<1><7> ), .B(n8), .Y(n1527) );
  NOR2X1 U641 ( .A(n964), .B(\addr_1c<4> ), .Y(n1820) );
  OAI21X1 U642 ( .A(n1040), .B(n972), .C(n1524), .Y(n1055) );
  NAND2X1 U643 ( .A(\mem<0><0> ), .B(n972), .Y(n1524) );
  OAI21X1 U644 ( .A(n1041), .B(n972), .C(n1523), .Y(n1054) );
  NAND2X1 U645 ( .A(\mem<0><1> ), .B(n972), .Y(n1523) );
  OAI21X1 U646 ( .A(n1042), .B(n972), .C(n1522), .Y(n1053) );
  NAND2X1 U647 ( .A(\mem<0><2> ), .B(n972), .Y(n1522) );
  OAI21X1 U648 ( .A(n1043), .B(n972), .C(n1521), .Y(n1052) );
  NAND2X1 U649 ( .A(\mem<0><3> ), .B(n972), .Y(n1521) );
  OAI21X1 U650 ( .A(n1044), .B(n972), .C(n1520), .Y(n1051) );
  NAND2X1 U651 ( .A(\mem<0><4> ), .B(n972), .Y(n1520) );
  OAI21X1 U652 ( .A(n1045), .B(n972), .C(n1519), .Y(n1050) );
  NAND2X1 U653 ( .A(\mem<0><5> ), .B(n972), .Y(n1519) );
  OAI21X1 U654 ( .A(n1046), .B(n972), .C(n1518), .Y(n1049) );
  NAND2X1 U655 ( .A(\mem<0><6> ), .B(n972), .Y(n1518) );
  OAI21X1 U656 ( .A(n1047), .B(n972), .C(n1517), .Y(n1048) );
  NAND2X1 U657 ( .A(\mem<0><7> ), .B(n972), .Y(n1517) );
  NAND3X1 U658 ( .A(n967), .B(n1013), .C(n1633), .Y(n1525) );
  NOR3X1 U661 ( .A(n1513), .B(\addr_1c<7> ), .C(\addr_1c<6> ), .Y(n1514) );
  NOR3X1 U662 ( .A(n1512), .B(\addr_1c<11> ), .C(\addr_1c<10> ), .Y(n1515) );
  AOI21X1 U663 ( .A(n461), .B(n1511), .C(n963), .Y(n1840) );
  OAI21X1 U665 ( .A(rd), .B(n1510), .C(wr), .Y(n1511) );
  NAND3X1 U667 ( .A(n1509), .B(n1027), .C(n1508), .Y(n1510) );
  NOR3X1 U668 ( .A(rd1), .B(rd3), .C(rd2), .Y(n1508) );
  NOR2X1 U669 ( .A(wr3), .B(wr2), .Y(n1509) );
  AOI21X1 U670 ( .A(n448), .B(n1506), .C(n1026), .Y(\data_out_1c<9> ) );
  NOR3X1 U671 ( .A(n2), .B(n1505), .C(n4), .Y(n1506) );
  AOI22X1 U673 ( .A(\mem<16><1> ), .B(n1788), .C(\mem<0><1> ), .D(n1633), .Y(
        n1503) );
  AOI22X1 U674 ( .A(\mem<18><1> ), .B(n1808), .C(\mem<2><1> ), .D(n1653), .Y(
        n1504) );
  AOI22X1 U676 ( .A(\mem<20><1> ), .B(n1788), .C(\mem<4><1> ), .D(n1633), .Y(
        n1501) );
  AOI22X1 U677 ( .A(\mem<22><1> ), .B(n1808), .C(\mem<6><1> ), .D(n1653), .Y(
        n1502) );
  AOI22X1 U678 ( .A(n1593), .B(n892), .C(n1632), .D(n932), .Y(n1507) );
  AOI22X1 U680 ( .A(\mem<28><1> ), .B(n1788), .C(\mem<12><1> ), .D(n1633), .Y(
        n1499) );
  AOI22X1 U681 ( .A(\mem<30><1> ), .B(n1808), .C(\mem<14><1> ), .D(n1653), .Y(
        n1500) );
  AOI22X1 U683 ( .A(\mem<24><1> ), .B(n1788), .C(\mem<8><1> ), .D(n1633), .Y(
        n1497) );
  AOI22X1 U684 ( .A(\mem<26><1> ), .B(n1808), .C(\mem<10><1> ), .D(n1653), .Y(
        n1498) );
  AOI21X1 U685 ( .A(n447), .B(n1495), .C(n1026), .Y(\data_out_1c<8> ) );
  NOR3X1 U686 ( .A(n939), .B(n1493), .C(n950), .Y(n1495) );
  AOI21X1 U687 ( .A(n1491), .B(n1490), .C(n971), .Y(n1492) );
  AOI22X1 U688 ( .A(\mem<16><0> ), .B(n1788), .C(\mem<0><0> ), .D(n1633), .Y(
        n1490) );
  AOI22X1 U689 ( .A(\mem<18><0> ), .B(n1808), .C(\mem<2><0> ), .D(n1653), .Y(
        n1491) );
  AOI21X1 U690 ( .A(n1489), .B(n1488), .C(n970), .Y(n1494) );
  AOI22X1 U691 ( .A(\mem<20><0> ), .B(n1788), .C(\mem<4><0> ), .D(n1633), .Y(
        n1488) );
  AOI22X1 U692 ( .A(\mem<22><0> ), .B(n1808), .C(\mem<6><0> ), .D(n1653), .Y(
        n1489) );
  AOI22X1 U693 ( .A(n1593), .B(n890), .C(n1632), .D(n930), .Y(n1496) );
  AOI22X1 U695 ( .A(\mem<28><0> ), .B(n1788), .C(\mem<12><0> ), .D(n1633), .Y(
        n1486) );
  AOI22X1 U696 ( .A(\mem<30><0> ), .B(n1808), .C(\mem<14><0> ), .D(n1653), .Y(
        n1487) );
  AOI22X1 U698 ( .A(\mem<24><0> ), .B(n1788), .C(\mem<8><0> ), .D(n1633), .Y(
        n1484) );
  AOI22X1 U699 ( .A(\mem<26><0> ), .B(n1808), .C(\mem<10><0> ), .D(n1653), .Y(
        n1485) );
  OAI21X1 U700 ( .A(n23), .B(n50), .C(rd1), .Y(n1483) );
  AOI22X1 U702 ( .A(\mem<17><7> ), .B(n1682), .C(\mem<19><7> ), .D(n1701), .Y(
        n1478) );
  AOI22X1 U703 ( .A(\mem<21><7> ), .B(n1720), .C(\mem<23><7> ), .D(n1739), .Y(
        n1479) );
  AOI22X1 U704 ( .A(\mem<25><7> ), .B(n1758), .C(\mem<27><7> ), .D(n1778), .Y(
        n1481) );
  AOI22X1 U705 ( .A(\mem<29><7> ), .B(n1798), .C(\mem<31><7> ), .D(n1819), .Y(
        n1482) );
  AOI22X1 U707 ( .A(\mem<1><7> ), .B(n1526), .C(\mem<3><7> ), .D(n1544), .Y(
        n1473) );
  AOI22X1 U708 ( .A(\mem<5><7> ), .B(n1564), .C(\mem<7><7> ), .D(n1583), .Y(
        n1474) );
  AOI22X1 U709 ( .A(\mem<9><7> ), .B(n1603), .C(\mem<11><7> ), .D(n1622), .Y(
        n1476) );
  AOI22X1 U710 ( .A(\mem<13><7> ), .B(n1643), .C(\mem<15><7> ), .D(n1663), .Y(
        n1477) );
  OAI21X1 U711 ( .A(n21), .B(n37), .C(rd1), .Y(n1472) );
  AOI22X1 U713 ( .A(\mem<17><6> ), .B(n1682), .C(\mem<19><6> ), .D(n1701), .Y(
        n1467) );
  AOI22X1 U714 ( .A(\mem<21><6> ), .B(n1720), .C(\mem<23><6> ), .D(n1739), .Y(
        n1468) );
  AOI22X1 U715 ( .A(\mem<25><6> ), .B(n1758), .C(\mem<27><6> ), .D(n1778), .Y(
        n1470) );
  AOI22X1 U716 ( .A(\mem<29><6> ), .B(n1798), .C(\mem<31><6> ), .D(n1819), .Y(
        n1471) );
  AOI22X1 U718 ( .A(\mem<1><6> ), .B(n1526), .C(\mem<3><6> ), .D(n1544), .Y(
        n1462) );
  AOI22X1 U719 ( .A(\mem<5><6> ), .B(n1564), .C(\mem<7><6> ), .D(n1583), .Y(
        n1463) );
  AOI22X1 U720 ( .A(\mem<9><6> ), .B(n1603), .C(\mem<11><6> ), .D(n1622), .Y(
        n1465) );
  AOI22X1 U721 ( .A(\mem<13><6> ), .B(n1643), .C(\mem<15><6> ), .D(n1663), .Y(
        n1466) );
  OAI21X1 U722 ( .A(n19), .B(n35), .C(rd1), .Y(n1461) );
  AOI22X1 U724 ( .A(\mem<17><5> ), .B(n1682), .C(\mem<19><5> ), .D(n1701), .Y(
        n1456) );
  AOI22X1 U725 ( .A(\mem<21><5> ), .B(n1720), .C(\mem<23><5> ), .D(n1739), .Y(
        n1457) );
  AOI22X1 U726 ( .A(\mem<25><5> ), .B(n1758), .C(\mem<27><5> ), .D(n1778), .Y(
        n1459) );
  AOI22X1 U727 ( .A(\mem<29><5> ), .B(n1798), .C(\mem<31><5> ), .D(n1819), .Y(
        n1460) );
  AOI22X1 U729 ( .A(\mem<1><5> ), .B(n1526), .C(\mem<3><5> ), .D(n1544), .Y(
        n1451) );
  AOI22X1 U730 ( .A(\mem<5><5> ), .B(n1564), .C(\mem<7><5> ), .D(n1583), .Y(
        n1452) );
  AOI22X1 U731 ( .A(\mem<9><5> ), .B(n1603), .C(\mem<11><5> ), .D(n1622), .Y(
        n1454) );
  AOI22X1 U732 ( .A(\mem<13><5> ), .B(n1643), .C(\mem<15><5> ), .D(n1663), .Y(
        n1455) );
  OAI21X1 U733 ( .A(n17), .B(n33), .C(rd1), .Y(n1450) );
  AOI22X1 U735 ( .A(\mem<17><4> ), .B(n1682), .C(\mem<19><4> ), .D(n1701), .Y(
        n1445) );
  AOI22X1 U736 ( .A(\mem<21><4> ), .B(n1720), .C(\mem<23><4> ), .D(n1739), .Y(
        n1446) );
  AOI22X1 U737 ( .A(\mem<25><4> ), .B(n1758), .C(\mem<27><4> ), .D(n1778), .Y(
        n1448) );
  AOI22X1 U738 ( .A(\mem<29><4> ), .B(n1798), .C(\mem<31><4> ), .D(n1819), .Y(
        n1449) );
  AOI22X1 U740 ( .A(\mem<1><4> ), .B(n1526), .C(\mem<3><4> ), .D(n1544), .Y(
        n1440) );
  AOI22X1 U741 ( .A(\mem<5><4> ), .B(n1564), .C(\mem<7><4> ), .D(n1583), .Y(
        n1441) );
  AOI22X1 U742 ( .A(\mem<9><4> ), .B(n1603), .C(\mem<11><4> ), .D(n1622), .Y(
        n1443) );
  AOI22X1 U743 ( .A(\mem<13><4> ), .B(n1643), .C(\mem<15><4> ), .D(n1663), .Y(
        n1444) );
  OAI21X1 U744 ( .A(n15), .B(n31), .C(rd1), .Y(n1439) );
  AOI22X1 U746 ( .A(\mem<17><3> ), .B(n1682), .C(\mem<19><3> ), .D(n1701), .Y(
        n1434) );
  AOI22X1 U747 ( .A(\mem<21><3> ), .B(n1720), .C(\mem<23><3> ), .D(n1739), .Y(
        n1435) );
  AOI22X1 U748 ( .A(\mem<25><3> ), .B(n1758), .C(\mem<27><3> ), .D(n1778), .Y(
        n1437) );
  AOI22X1 U749 ( .A(\mem<29><3> ), .B(n1798), .C(\mem<31><3> ), .D(n1819), .Y(
        n1438) );
  AOI22X1 U751 ( .A(\mem<1><3> ), .B(n1526), .C(\mem<3><3> ), .D(n1544), .Y(
        n1429) );
  AOI22X1 U752 ( .A(\mem<5><3> ), .B(n1564), .C(\mem<7><3> ), .D(n1583), .Y(
        n1430) );
  AOI22X1 U753 ( .A(\mem<9><3> ), .B(n1603), .C(\mem<11><3> ), .D(n1622), .Y(
        n1432) );
  AOI22X1 U754 ( .A(\mem<13><3> ), .B(n1643), .C(\mem<15><3> ), .D(n1663), .Y(
        n1433) );
  OAI21X1 U755 ( .A(n13), .B(n29), .C(rd1), .Y(n1428) );
  AOI22X1 U757 ( .A(\mem<17><2> ), .B(n1682), .C(\mem<19><2> ), .D(n1701), .Y(
        n1423) );
  AOI22X1 U758 ( .A(\mem<21><2> ), .B(n1720), .C(\mem<23><2> ), .D(n1739), .Y(
        n1424) );
  AOI22X1 U759 ( .A(\mem<25><2> ), .B(n1758), .C(\mem<27><2> ), .D(n1778), .Y(
        n1426) );
  AOI22X1 U760 ( .A(\mem<29><2> ), .B(n1798), .C(\mem<31><2> ), .D(n1819), .Y(
        n1427) );
  AOI22X1 U762 ( .A(\mem<1><2> ), .B(n1526), .C(\mem<3><2> ), .D(n1544), .Y(
        n1418) );
  AOI22X1 U763 ( .A(\mem<5><2> ), .B(n1564), .C(\mem<7><2> ), .D(n1583), .Y(
        n1419) );
  AOI22X1 U764 ( .A(\mem<9><2> ), .B(n1603), .C(\mem<11><2> ), .D(n1622), .Y(
        n1421) );
  AOI22X1 U765 ( .A(\mem<13><2> ), .B(n1643), .C(\mem<15><2> ), .D(n1663), .Y(
        n1422) );
  OAI21X1 U766 ( .A(n11), .B(n27), .C(rd1), .Y(n1417) );
  AOI22X1 U768 ( .A(\mem<17><1> ), .B(n1682), .C(\mem<19><1> ), .D(n1701), .Y(
        n1412) );
  AOI22X1 U769 ( .A(\mem<21><1> ), .B(n1720), .C(\mem<23><1> ), .D(n1739), .Y(
        n1413) );
  AOI22X1 U770 ( .A(\mem<25><1> ), .B(n1758), .C(\mem<27><1> ), .D(n1778), .Y(
        n1415) );
  AOI22X1 U771 ( .A(\mem<29><1> ), .B(n1798), .C(\mem<31><1> ), .D(n1819), .Y(
        n1416) );
  AOI22X1 U773 ( .A(\mem<1><1> ), .B(n1526), .C(\mem<3><1> ), .D(n1544), .Y(
        n1407) );
  AOI22X1 U774 ( .A(\mem<5><1> ), .B(n1564), .C(\mem<7><1> ), .D(n1583), .Y(
        n1408) );
  AOI22X1 U775 ( .A(\mem<9><1> ), .B(n1603), .C(\mem<11><1> ), .D(n1622), .Y(
        n1410) );
  AOI22X1 U776 ( .A(\mem<13><1> ), .B(n1643), .C(\mem<15><1> ), .D(n1663), .Y(
        n1411) );
  AOI21X1 U777 ( .A(n435), .B(n1405), .C(n1026), .Y(\data_out_1c<15> ) );
  NOR3X1 U778 ( .A(n938), .B(n1403), .C(n949), .Y(n1405) );
  AOI21X1 U779 ( .A(n1401), .B(n1400), .C(n971), .Y(n1402) );
  AOI22X1 U780 ( .A(\mem<16><7> ), .B(n1788), .C(\mem<0><7> ), .D(n1633), .Y(
        n1400) );
  AOI22X1 U781 ( .A(\mem<18><7> ), .B(n1808), .C(\mem<2><7> ), .D(n1653), .Y(
        n1401) );
  AOI21X1 U782 ( .A(n1399), .B(n1398), .C(n970), .Y(n1404) );
  AOI22X1 U783 ( .A(\mem<20><7> ), .B(n1788), .C(\mem<4><7> ), .D(n1633), .Y(
        n1398) );
  AOI22X1 U784 ( .A(\mem<22><7> ), .B(n1808), .C(\mem<6><7> ), .D(n1653), .Y(
        n1399) );
  AOI22X1 U785 ( .A(n1593), .B(n888), .C(n1632), .D(n928), .Y(n1406) );
  AOI22X1 U787 ( .A(\mem<28><7> ), .B(n1788), .C(\mem<12><7> ), .D(n1633), .Y(
        n1396) );
  AOI22X1 U788 ( .A(\mem<30><7> ), .B(n1808), .C(\mem<14><7> ), .D(n1653), .Y(
        n1397) );
  AOI22X1 U790 ( .A(\mem<24><7> ), .B(n1788), .C(\mem<8><7> ), .D(n1633), .Y(
        n1394) );
  AOI22X1 U791 ( .A(\mem<26><7> ), .B(n1808), .C(\mem<10><7> ), .D(n1653), .Y(
        n1395) );
  AOI21X1 U792 ( .A(n434), .B(n1392), .C(n1026), .Y(\data_out_1c<14> ) );
  NOR3X1 U793 ( .A(n937), .B(n1390), .C(n948), .Y(n1392) );
  AOI21X1 U794 ( .A(n1388), .B(n1387), .C(n971), .Y(n1389) );
  AOI22X1 U795 ( .A(\mem<16><6> ), .B(n1788), .C(\mem<0><6> ), .D(n1633), .Y(
        n1387) );
  AOI22X1 U796 ( .A(\mem<18><6> ), .B(n1808), .C(\mem<2><6> ), .D(n1653), .Y(
        n1388) );
  AOI21X1 U797 ( .A(n1386), .B(n1385), .C(n970), .Y(n1391) );
  AOI22X1 U798 ( .A(\mem<20><6> ), .B(n1788), .C(\mem<4><6> ), .D(n1633), .Y(
        n1385) );
  AOI22X1 U799 ( .A(\mem<22><6> ), .B(n1808), .C(\mem<6><6> ), .D(n1653), .Y(
        n1386) );
  AOI22X1 U800 ( .A(n1593), .B(n886), .C(n1632), .D(n926), .Y(n1393) );
  AOI22X1 U802 ( .A(\mem<28><6> ), .B(n1788), .C(\mem<12><6> ), .D(n1633), .Y(
        n1383) );
  AOI22X1 U803 ( .A(\mem<30><6> ), .B(n1808), .C(\mem<14><6> ), .D(n1653), .Y(
        n1384) );
  AOI22X1 U805 ( .A(\mem<24><6> ), .B(n1788), .C(\mem<8><6> ), .D(n1633), .Y(
        n1381) );
  AOI22X1 U806 ( .A(\mem<26><6> ), .B(n1808), .C(\mem<10><6> ), .D(n1653), .Y(
        n1382) );
  AOI21X1 U807 ( .A(n422), .B(n1379), .C(n1026), .Y(\data_out_1c<13> ) );
  NOR3X1 U808 ( .A(n936), .B(n1377), .C(n947), .Y(n1379) );
  AOI21X1 U809 ( .A(n1375), .B(n1374), .C(n971), .Y(n1376) );
  AOI22X1 U810 ( .A(\mem<16><5> ), .B(n1788), .C(\mem<0><5> ), .D(n1633), .Y(
        n1374) );
  AOI22X1 U811 ( .A(\mem<18><5> ), .B(n1808), .C(\mem<2><5> ), .D(n1653), .Y(
        n1375) );
  AOI21X1 U812 ( .A(n1373), .B(n1372), .C(n970), .Y(n1378) );
  AOI22X1 U813 ( .A(\mem<20><5> ), .B(n1788), .C(\mem<4><5> ), .D(n1633), .Y(
        n1372) );
  AOI22X1 U814 ( .A(\mem<22><5> ), .B(n1808), .C(\mem<6><5> ), .D(n1653), .Y(
        n1373) );
  AOI22X1 U815 ( .A(n1593), .B(n884), .C(n1632), .D(n924), .Y(n1380) );
  AOI22X1 U817 ( .A(\mem<28><5> ), .B(n1788), .C(\mem<12><5> ), .D(n1633), .Y(
        n1370) );
  AOI22X1 U818 ( .A(\mem<30><5> ), .B(n1808), .C(\mem<14><5> ), .D(n1653), .Y(
        n1371) );
  AOI22X1 U820 ( .A(\mem<24><5> ), .B(n1788), .C(\mem<8><5> ), .D(n1633), .Y(
        n1368) );
  AOI22X1 U821 ( .A(\mem<26><5> ), .B(n1808), .C(\mem<10><5> ), .D(n1653), .Y(
        n1369) );
  AOI21X1 U822 ( .A(n421), .B(n1366), .C(n1026), .Y(\data_out_1c<12> ) );
  NOR3X1 U823 ( .A(n935), .B(n1364), .C(n946), .Y(n1366) );
  AOI21X1 U824 ( .A(n1362), .B(n1361), .C(n971), .Y(n1363) );
  AOI22X1 U825 ( .A(\mem<16><4> ), .B(n1788), .C(\mem<0><4> ), .D(n1633), .Y(
        n1361) );
  AOI22X1 U826 ( .A(\mem<18><4> ), .B(n1808), .C(\mem<2><4> ), .D(n1653), .Y(
        n1362) );
  AOI21X1 U827 ( .A(n1360), .B(n1359), .C(n970), .Y(n1365) );
  AOI22X1 U828 ( .A(\mem<20><4> ), .B(n1788), .C(\mem<4><4> ), .D(n1633), .Y(
        n1359) );
  AOI22X1 U829 ( .A(\mem<22><4> ), .B(n1808), .C(\mem<6><4> ), .D(n1653), .Y(
        n1360) );
  AOI22X1 U830 ( .A(n1593), .B(n882), .C(n1632), .D(n922), .Y(n1367) );
  AOI22X1 U832 ( .A(\mem<28><4> ), .B(n1788), .C(\mem<12><4> ), .D(n1633), .Y(
        n1357) );
  AOI22X1 U833 ( .A(\mem<30><4> ), .B(n1808), .C(\mem<14><4> ), .D(n1653), .Y(
        n1358) );
  AOI22X1 U835 ( .A(\mem<24><4> ), .B(n1788), .C(\mem<8><4> ), .D(n1633), .Y(
        n1355) );
  AOI22X1 U836 ( .A(\mem<26><4> ), .B(n1808), .C(\mem<10><4> ), .D(n1653), .Y(
        n1356) );
  AOI21X1 U837 ( .A(n409), .B(n1353), .C(n1026), .Y(\data_out_1c<11> ) );
  NOR3X1 U838 ( .A(n934), .B(n1351), .C(n945), .Y(n1353) );
  AOI21X1 U839 ( .A(n1349), .B(n1348), .C(n971), .Y(n1350) );
  AOI22X1 U840 ( .A(\mem<16><3> ), .B(n1788), .C(\mem<0><3> ), .D(n1633), .Y(
        n1348) );
  AOI22X1 U841 ( .A(\mem<18><3> ), .B(n1808), .C(\mem<2><3> ), .D(n1653), .Y(
        n1349) );
  AOI21X1 U842 ( .A(n1347), .B(n1346), .C(n970), .Y(n1352) );
  AOI22X1 U843 ( .A(\mem<20><3> ), .B(n1788), .C(\mem<4><3> ), .D(n1633), .Y(
        n1346) );
  AOI22X1 U844 ( .A(\mem<22><3> ), .B(n1808), .C(\mem<6><3> ), .D(n1653), .Y(
        n1347) );
  AOI22X1 U845 ( .A(n1593), .B(n880), .C(n1632), .D(n920), .Y(n1354) );
  AOI22X1 U847 ( .A(\mem<28><3> ), .B(n1788), .C(\mem<12><3> ), .D(n1633), .Y(
        n1344) );
  AOI22X1 U848 ( .A(\mem<30><3> ), .B(n1808), .C(\mem<14><3> ), .D(n1653), .Y(
        n1345) );
  AOI22X1 U850 ( .A(\mem<24><3> ), .B(n1788), .C(\mem<8><3> ), .D(n1633), .Y(
        n1342) );
  AOI22X1 U851 ( .A(\mem<26><3> ), .B(n1808), .C(\mem<10><3> ), .D(n1653), .Y(
        n1343) );
  AOI21X1 U852 ( .A(n408), .B(n1340), .C(n1026), .Y(\data_out_1c<10> ) );
  NOR3X1 U853 ( .A(n933), .B(n1338), .C(n944), .Y(n1340) );
  AOI21X1 U854 ( .A(n1336), .B(n1335), .C(n971), .Y(n1337) );
  AOI22X1 U855 ( .A(\mem<16><2> ), .B(n1788), .C(\mem<0><2> ), .D(n1633), .Y(
        n1335) );
  AOI22X1 U856 ( .A(\mem<18><2> ), .B(n1808), .C(\mem<2><2> ), .D(n1653), .Y(
        n1336) );
  AOI21X1 U857 ( .A(n1334), .B(n1333), .C(n970), .Y(n1339) );
  AOI22X1 U858 ( .A(\mem<20><2> ), .B(n1788), .C(\mem<4><2> ), .D(n1633), .Y(
        n1333) );
  AOI22X1 U859 ( .A(\mem<22><2> ), .B(n1808), .C(\mem<6><2> ), .D(n1653), .Y(
        n1334) );
  AOI22X1 U860 ( .A(n1593), .B(n878), .C(n1632), .D(n918), .Y(n1341) );
  AOI22X1 U862 ( .A(\mem<28><2> ), .B(n1788), .C(\mem<12><2> ), .D(n1633), .Y(
        n1331) );
  AOI22X1 U863 ( .A(\mem<30><2> ), .B(n1808), .C(\mem<14><2> ), .D(n1653), .Y(
        n1332) );
  AOI22X1 U865 ( .A(\mem<24><2> ), .B(n1788), .C(\mem<8><2> ), .D(n1633), .Y(
        n1329) );
  AOI22X1 U866 ( .A(\mem<26><2> ), .B(n1808), .C(\mem<10><2> ), .D(n1653), .Y(
        n1330) );
  NOR2X1 U867 ( .A(\addr_1c<3> ), .B(\addr_1c<4> ), .Y(n1328) );
  NOR2X1 U868 ( .A(n1031), .B(\addr_1c<4> ), .Y(n1327) );
  OAI21X1 U869 ( .A(n9), .B(n25), .C(rd1), .Y(n1326) );
  AOI22X1 U871 ( .A(\mem<17><0> ), .B(n1682), .C(\mem<19><0> ), .D(n1701), .Y(
        n1321) );
  AOI22X1 U872 ( .A(\mem<21><0> ), .B(n1720), .C(\mem<23><0> ), .D(n1739), .Y(
        n1322) );
  AOI22X1 U873 ( .A(\mem<25><0> ), .B(n1758), .C(\mem<27><0> ), .D(n1778), .Y(
        n1324) );
  AOI22X1 U874 ( .A(\mem<29><0> ), .B(n1798), .C(\mem<31><0> ), .D(n1819), .Y(
        n1325) );
  AOI22X1 U876 ( .A(\mem<1><0> ), .B(n1526), .C(\mem<3><0> ), .D(n1544), .Y(
        n1314) );
  NAND2X1 U877 ( .A(n1029), .B(n1030), .Y(n1516) );
  AOI22X1 U878 ( .A(\mem<5><0> ), .B(n1564), .C(\mem<7><0> ), .D(n1583), .Y(
        n1315) );
  NAND2X1 U879 ( .A(\addr_1c<1> ), .B(n1030), .Y(n1554) );
  AOI22X1 U880 ( .A(\mem<9><0> ), .B(n1603), .C(\mem<11><0> ), .D(n1622), .Y(
        n1317) );
  AOI22X1 U881 ( .A(\mem<13><0> ), .B(n1643), .C(\mem<15><0> ), .D(n1663), .Y(
        n1318) );
  dff_50 ff0 ( .q(rd1), .d(rd0), .clk(clk), .rst(rst) );
  dff_49 ff1 ( .q(wr1), .d(wr0), .clk(clk), .rst(rst) );
  dff_48 \reg0[0]  ( .q(\addr_1c<0> ), .d(\addr<0> ), .clk(clk), .rst(rst) );
  dff_47 \reg0[1]  ( .q(\addr_1c<1> ), .d(\addr<1> ), .clk(clk), .rst(rst) );
  dff_46 \reg0[2]  ( .q(\addr_1c<2> ), .d(\addr<2> ), .clk(clk), .rst(rst) );
  dff_45 \reg0[3]  ( .q(\addr_1c<3> ), .d(\addr<3> ), .clk(clk), .rst(rst) );
  dff_44 \reg0[4]  ( .q(\addr_1c<4> ), .d(\addr<4> ), .clk(clk), .rst(rst) );
  dff_43 \reg0[5]  ( .q(\addr_1c<5> ), .d(\addr<5> ), .clk(clk), .rst(rst) );
  dff_42 \reg0[6]  ( .q(\addr_1c<6> ), .d(\addr<6> ), .clk(clk), .rst(rst) );
  dff_41 \reg0[7]  ( .q(\addr_1c<7> ), .d(\addr<7> ), .clk(clk), .rst(rst) );
  dff_40 \reg0[8]  ( .q(\addr_1c<8> ), .d(\addr<8> ), .clk(clk), .rst(rst) );
  dff_39 \reg0[9]  ( .q(\addr_1c<9> ), .d(\addr<9> ), .clk(clk), .rst(rst) );
  dff_38 \reg0[10]  ( .q(\addr_1c<10> ), .d(\addr<10> ), .clk(clk), .rst(rst)
         );
  dff_37 \reg0[11]  ( .q(\addr_1c<11> ), .d(\addr<11> ), .clk(clk), .rst(rst)
         );
  dff_36 \reg0[12]  ( .q(\addr_1c<12> ), .d(\addr<12> ), .clk(clk), .rst(rst)
         );
  dff_35 \reg1[0]  ( .q(\data_in_1c<0> ), .d(\data_in<0> ), .clk(clk), .rst(
        rst) );
  dff_34 \reg1[1]  ( .q(\data_in_1c<1> ), .d(\data_in<1> ), .clk(clk), .rst(
        rst) );
  dff_33 \reg1[2]  ( .q(\data_in_1c<2> ), .d(\data_in<2> ), .clk(clk), .rst(
        rst) );
  dff_32 \reg1[3]  ( .q(\data_in_1c<3> ), .d(\data_in<3> ), .clk(clk), .rst(
        rst) );
  dff_31 \reg1[4]  ( .q(\data_in_1c<4> ), .d(\data_in<4> ), .clk(clk), .rst(
        rst) );
  dff_30 \reg1[5]  ( .q(\data_in_1c<5> ), .d(\data_in<5> ), .clk(clk), .rst(
        rst) );
  dff_29 \reg1[6]  ( .q(\data_in_1c<6> ), .d(\data_in<6> ), .clk(clk), .rst(
        rst) );
  dff_28 \reg1[7]  ( .q(\data_in_1c<7> ), .d(\data_in<7> ), .clk(clk), .rst(
        rst) );
  dff_27 \reg1[8]  ( .q(\data_in_1c<8> ), .d(\data_in<8> ), .clk(clk), .rst(
        rst) );
  dff_26 \reg1[9]  ( .q(\data_in_1c<9> ), .d(\data_in<9> ), .clk(clk), .rst(
        rst) );
  dff_25 \reg1[10]  ( .q(\data_in_1c<10> ), .d(\data_in<10> ), .clk(clk), 
        .rst(rst) );
  dff_24 \reg1[11]  ( .q(\data_in_1c<11> ), .d(\data_in<11> ), .clk(clk), 
        .rst(rst) );
  dff_23 \reg1[12]  ( .q(\data_in_1c<12> ), .d(\data_in<12> ), .clk(clk), 
        .rst(rst) );
  dff_22 \reg1[13]  ( .q(\data_in_1c<13> ), .d(\data_in<13> ), .clk(clk), 
        .rst(rst) );
  dff_21 \reg1[14]  ( .q(\data_in_1c<14> ), .d(\data_in<14> ), .clk(clk), 
        .rst(rst) );
  dff_20 \reg1[15]  ( .q(\data_in_1c<15> ), .d(\data_in<15> ), .clk(clk), 
        .rst(rst) );
  dff_19 \reg2[0]  ( .q(\data_out<0> ), .d(n1023), .clk(clk), .rst(rst) );
  dff_18 \reg2[1]  ( .q(\data_out<1> ), .d(n1022), .clk(clk), .rst(rst) );
  dff_17 \reg2[2]  ( .q(\data_out<2> ), .d(n1021), .clk(clk), .rst(rst) );
  dff_16 \reg2[3]  ( .q(\data_out<3> ), .d(n1020), .clk(clk), .rst(rst) );
  dff_15 \reg2[4]  ( .q(\data_out<4> ), .d(n1019), .clk(clk), .rst(rst) );
  dff_14 \reg2[5]  ( .q(\data_out<5> ), .d(n1018), .clk(clk), .rst(rst) );
  dff_13 \reg2[6]  ( .q(\data_out<6> ), .d(n1017), .clk(clk), .rst(rst) );
  dff_12 \reg2[7]  ( .q(\data_out<7> ), .d(n1016), .clk(clk), .rst(rst) );
  dff_11 \reg2[8]  ( .q(\data_out<8> ), .d(\data_out_1c<8> ), .clk(clk), .rst(
        rst) );
  dff_10 \reg2[9]  ( .q(\data_out<9> ), .d(\data_out_1c<9> ), .clk(clk), .rst(
        rst) );
  dff_9 \reg2[10]  ( .q(\data_out<10> ), .d(\data_out_1c<10> ), .clk(clk), 
        .rst(rst) );
  dff_8 \reg2[11]  ( .q(\data_out<11> ), .d(\data_out_1c<11> ), .clk(clk), 
        .rst(rst) );
  dff_7 \reg2[12]  ( .q(\data_out<12> ), .d(\data_out_1c<12> ), .clk(clk), 
        .rst(rst) );
  dff_6 \reg2[13]  ( .q(\data_out<13> ), .d(\data_out_1c<13> ), .clk(clk), 
        .rst(rst) );
  dff_5 \reg2[14]  ( .q(\data_out<14> ), .d(\data_out_1c<14> ), .clk(clk), 
        .rst(rst) );
  dff_4 \reg2[15]  ( .q(\data_out<15> ), .d(\data_out_1c<15> ), .clk(clk), 
        .rst(rst) );
  dff_3 ff2 ( .q(rd2), .d(rd1), .clk(clk), .rst(rst) );
  dff_2 ff3 ( .q(wr2), .d(wr1), .clk(clk), .rst(rst) );
  dff_1 ff4 ( .q(rd3), .d(rd2), .clk(clk), .rst(rst) );
  dff_0 ff5 ( .q(wr3), .d(wr2), .clk(clk), .rst(rst) );
  INVX1 U2 ( .A(rd), .Y(n1025) );
  OR2X1 U3 ( .A(\addr_1c<5> ), .B(\addr_1c<12> ), .Y(n1512) );
  AND2X1 U4 ( .A(\addr_1c<4> ), .B(n1526), .Y(n1829) );
  INVX1 U5 ( .A(\addr_1c<3> ), .Y(n1031) );
  INVX1 U6 ( .A(\addr_1c<2> ), .Y(n1030) );
  OR2X1 U7 ( .A(\addr_1c<9> ), .B(\addr_1c<8> ), .Y(n1513) );
  AND2X1 U8 ( .A(n1632), .B(n965), .Y(n1809) );
  AND2X1 U23 ( .A(n1593), .B(n965), .Y(n1768) );
  INVX1 U24 ( .A(\addr_1c<0> ), .Y(n1028) );
  AND2X1 U25 ( .A(n1028), .B(n1031), .Y(n1312) );
  AND2X1 U26 ( .A(\addr_1c<0> ), .B(n1031), .Y(n1313) );
  AND2X1 U27 ( .A(\addr_1c<3> ), .B(\addr_1c<0> ), .Y(n1320) );
  AND2X1 U28 ( .A(\addr_1c<3> ), .B(n1028), .Y(n1319) );
  INVX1 U29 ( .A(\addr_1c<1> ), .Y(n1029) );
  INVX1 U35 ( .A(wr1), .Y(n1027) );
  AND2X1 U36 ( .A(n1593), .B(n1320), .Y(n1778) );
  AND2X1 U37 ( .A(n1593), .B(n1319), .Y(n1758) );
  AND2X1 U38 ( .A(n940), .B(n1320), .Y(n1739) );
  AND2X1 U39 ( .A(n940), .B(n1319), .Y(n1720) );
  AND2X1 U40 ( .A(n1320), .B(n951), .Y(n1701) );
  AND2X1 U41 ( .A(n1319), .B(n951), .Y(n1682) );
  AND2X1 U42 ( .A(n1313), .B(n1593), .Y(n1622) );
  AND2X1 U43 ( .A(n1593), .B(n1312), .Y(n1603) );
  AND2X1 U44 ( .A(n1313), .B(n940), .Y(n1583) );
  AND2X1 U46 ( .A(n940), .B(n1312), .Y(n1564) );
  OR2X1 U47 ( .A(n970), .B(n964), .Y(n968) );
  AND2X1 U48 ( .A(n1313), .B(n951), .Y(n1544) );
  AND2X1 U49 ( .A(wr1), .B(n1015), .Y(n1830) );
  OR2X1 U50 ( .A(n964), .B(n971), .Y(n966) );
  AND2X1 U51 ( .A(n1632), .B(n1312), .Y(n1643) );
  AND2X1 U52 ( .A(n1313), .B(n1632), .Y(n1663) );
  AND2X1 U53 ( .A(n1319), .B(n1632), .Y(n1798) );
  AND2X1 U54 ( .A(\addr_1c<2> ), .B(n1029), .Y(n1593) );
  AND2X1 U55 ( .A(\addr_1c<2> ), .B(\addr_1c<1> ), .Y(n1632) );
  BUFX2 U56 ( .A(n961), .Y(n1010) );
  BUFX2 U57 ( .A(n961), .Y(n1009) );
  BUFX2 U58 ( .A(n960), .Y(n1007) );
  BUFX2 U59 ( .A(n960), .Y(n1006) );
  BUFX2 U60 ( .A(n959), .Y(n1004) );
  BUFX2 U61 ( .A(n959), .Y(n1003) );
  BUFX2 U62 ( .A(n958), .Y(n1001) );
  BUFX2 U63 ( .A(n958), .Y(n1000) );
  BUFX2 U64 ( .A(n957), .Y(n990) );
  BUFX2 U65 ( .A(n957), .Y(n989) );
  BUFX2 U66 ( .A(n956), .Y(n987) );
  BUFX2 U67 ( .A(n956), .Y(n986) );
  BUFX2 U68 ( .A(n955), .Y(n984) );
  BUFX2 U69 ( .A(n955), .Y(n983) );
  BUFX2 U70 ( .A(n954), .Y(n981) );
  BUFX2 U71 ( .A(n954), .Y(n980) );
  INVX1 U72 ( .A(\data_in_1c<0> ), .Y(n1032) );
  INVX1 U73 ( .A(\data_in_1c<1> ), .Y(n1033) );
  INVX1 U74 ( .A(\data_in_1c<2> ), .Y(n1034) );
  INVX1 U75 ( .A(\data_in_1c<3> ), .Y(n1035) );
  INVX1 U76 ( .A(\data_in_1c<4> ), .Y(n1036) );
  INVX1 U77 ( .A(\data_in_1c<5> ), .Y(n1037) );
  INVX1 U78 ( .A(\data_in_1c<6> ), .Y(n1038) );
  INVX1 U79 ( .A(\data_in_1c<7> ), .Y(n1039) );
  INVX1 U80 ( .A(\data_in_1c<8> ), .Y(n1040) );
  INVX1 U81 ( .A(\data_in_1c<9> ), .Y(n1041) );
  INVX1 U82 ( .A(\data_in_1c<10> ), .Y(n1042) );
  INVX1 U83 ( .A(\data_in_1c<11> ), .Y(n1043) );
  INVX1 U84 ( .A(\data_in_1c<12> ), .Y(n1044) );
  INVX1 U85 ( .A(\data_in_1c<13> ), .Y(n1045) );
  INVX1 U86 ( .A(\data_in_1c<14> ), .Y(n1046) );
  INVX1 U87 ( .A(\data_in_1c<15> ), .Y(n1047) );
  AND2X1 U88 ( .A(n1829), .B(\mem<32><0> ), .Y(n1493) );
  AND2X1 U89 ( .A(n1829), .B(\mem<32><1> ), .Y(n1505) );
  AND2X1 U90 ( .A(n1829), .B(\mem<32><2> ), .Y(n1338) );
  AND2X1 U91 ( .A(n1829), .B(\mem<32><3> ), .Y(n1351) );
  AND2X1 U92 ( .A(n1829), .B(\mem<32><4> ), .Y(n1364) );
  AND2X1 U93 ( .A(n1829), .B(\mem<32><5> ), .Y(n1377) );
  AND2X1 U129 ( .A(n1829), .B(\mem<32><6> ), .Y(n1390) );
  AND2X1 U589 ( .A(n1829), .B(\mem<32><7> ), .Y(n1403) );
  INVX1 U640 ( .A(rd1), .Y(n1026) );
  INVX1 U659 ( .A(wr), .Y(n1024) );
  INVX1 U660 ( .A(n1326), .Y(n1023) );
  INVX1 U664 ( .A(n1417), .Y(n1022) );
  INVX1 U666 ( .A(n1428), .Y(n1021) );
  INVX1 U672 ( .A(n1439), .Y(n1020) );
  INVX1 U675 ( .A(n1450), .Y(n1019) );
  INVX1 U679 ( .A(n1461), .Y(n1018) );
  INVX1 U682 ( .A(n1472), .Y(n1017) );
  INVX1 U694 ( .A(n1483), .Y(n1016) );
  INVX1 U697 ( .A(n1830), .Y(n1014) );
  INVX1 U701 ( .A(rst), .Y(n1015) );
  INVX1 U706 ( .A(n1014), .Y(n1012) );
  INVX1 U712 ( .A(n1014), .Y(n1013) );
  AND2X1 U717 ( .A(n387), .B(n372), .Y(n1) );
  INVX1 U723 ( .A(n1), .Y(n2) );
  AND2X1 U728 ( .A(n402), .B(n381), .Y(n3) );
  INVX1 U734 ( .A(n3), .Y(n4) );
  AND2X1 U739 ( .A(n1819), .B(n189), .Y(n5) );
  INVX1 U745 ( .A(n5), .Y(n6) );
  AND2X1 U750 ( .A(n973), .B(n289), .Y(n7) );
  INVX1 U756 ( .A(n7), .Y(n8) );
  OR2X1 U761 ( .A(n486), .B(n10), .Y(n9) );
  OR2X1 U767 ( .A(n473), .B(n474), .Y(n10) );
  OR2X1 U772 ( .A(n508), .B(n12), .Y(n11) );
  OR2X1 U786 ( .A(n487), .B(n507), .Y(n12) );
  OR2X1 U789 ( .A(n537), .B(n14), .Y(n13) );
  OR2X1 U801 ( .A(n522), .B(n523), .Y(n14) );
  OR2X1 U804 ( .A(n553), .B(n16), .Y(n15) );
  OR2X1 U816 ( .A(n538), .B(n552), .Y(n16) );
  OR2X1 U819 ( .A(n582), .B(n18), .Y(n17) );
  OR2X1 U831 ( .A(n567), .B(n568), .Y(n18) );
  OR2X1 U834 ( .A(n592), .B(n20), .Y(n19) );
  OR2X1 U846 ( .A(n583), .B(n591), .Y(n20) );
  OR2X1 U849 ( .A(n873), .B(n22), .Y(n21) );
  OR2X1 U861 ( .A(n871), .B(n872), .Y(n22) );
  OR2X1 U864 ( .A(n876), .B(n24), .Y(n23) );
  OR2X1 U870 ( .A(n874), .B(n875), .Y(n24) );
  OR2X1 U875 ( .A(n895), .B(n26), .Y(n25) );
  OR2X1 U882 ( .A(n893), .B(n894), .Y(n26) );
  OR2X1 U883 ( .A(n898), .B(n28), .Y(n27) );
  OR2X1 U884 ( .A(n896), .B(n897), .Y(n28) );
  OR2X1 U885 ( .A(n901), .B(n30), .Y(n29) );
  OR2X1 U886 ( .A(n899), .B(n900), .Y(n30) );
  OR2X1 U887 ( .A(n904), .B(n32), .Y(n31) );
  OR2X1 U888 ( .A(n902), .B(n903), .Y(n32) );
  OR2X1 U889 ( .A(n907), .B(n34), .Y(n33) );
  OR2X1 U890 ( .A(n905), .B(n906), .Y(n34) );
  OR2X1 U891 ( .A(n910), .B(n36), .Y(n35) );
  OR2X1 U892 ( .A(n908), .B(n909), .Y(n36) );
  OR2X1 U893 ( .A(n913), .B(n38), .Y(n37) );
  OR2X1 U894 ( .A(n911), .B(n912), .Y(n38) );
  OR2X1 U895 ( .A(n916), .B(n150), .Y(n50) );
  OR2X1 U896 ( .A(n914), .B(n915), .Y(n150) );
  AND2X1 U897 ( .A(n973), .B(n1830), .Y(n189) );
  AND2X1 U898 ( .A(n1830), .B(n1526), .Y(n289) );
  AND2X1 U899 ( .A(n940), .B(n942), .Y(n348) );
  INVX1 U900 ( .A(n348), .Y(n372) );
  AND2X1 U901 ( .A(n951), .B(n953), .Y(n379) );
  INVX1 U902 ( .A(n379), .Y(n381) );
  AND2X1 U903 ( .A(n940), .B(n941), .Y(n386) );
  INVX1 U904 ( .A(n386), .Y(n387) );
  AND2X1 U905 ( .A(n951), .B(n952), .Y(n401) );
  INVX1 U906 ( .A(n401), .Y(n402) );
  BUFX2 U907 ( .A(n1341), .Y(n408) );
  BUFX2 U908 ( .A(n1354), .Y(n409) );
  BUFX2 U909 ( .A(n1367), .Y(n421) );
  BUFX2 U910 ( .A(n1380), .Y(n422) );
  BUFX2 U911 ( .A(n1393), .Y(n434) );
  BUFX2 U912 ( .A(n1406), .Y(n435) );
  BUFX2 U913 ( .A(n1496), .Y(n447) );
  BUFX2 U914 ( .A(n1507), .Y(n448) );
  AND2X2 U915 ( .A(rd), .B(n1510), .Y(n460) );
  INVX1 U916 ( .A(n460), .Y(n461) );
  INVX1 U917 ( .A(n1316), .Y(n473) );
  INVX1 U918 ( .A(n1317), .Y(n474) );
  INVX1 U919 ( .A(n1318), .Y(n486) );
  INVX1 U920 ( .A(n1409), .Y(n487) );
  INVX1 U921 ( .A(n1410), .Y(n507) );
  INVX1 U922 ( .A(n1411), .Y(n508) );
  INVX1 U923 ( .A(n1420), .Y(n522) );
  INVX1 U924 ( .A(n1421), .Y(n523) );
  INVX1 U925 ( .A(n1422), .Y(n537) );
  INVX1 U926 ( .A(n1431), .Y(n538) );
  INVX1 U927 ( .A(n1432), .Y(n552) );
  INVX1 U928 ( .A(n1433), .Y(n553) );
  INVX1 U929 ( .A(n1442), .Y(n567) );
  INVX1 U930 ( .A(n1443), .Y(n568) );
  INVX1 U931 ( .A(n1444), .Y(n582) );
  INVX1 U932 ( .A(n1453), .Y(n583) );
  INVX1 U933 ( .A(n1454), .Y(n591) );
  INVX1 U934 ( .A(n1455), .Y(n592) );
  INVX1 U935 ( .A(n1464), .Y(n871) );
  INVX1 U936 ( .A(n1465), .Y(n872) );
  INVX1 U937 ( .A(n1466), .Y(n873) );
  INVX1 U938 ( .A(n1475), .Y(n874) );
  INVX1 U939 ( .A(n1476), .Y(n875) );
  INVX1 U940 ( .A(n1477), .Y(n876) );
  AND2X2 U941 ( .A(n1330), .B(n1329), .Y(n877) );
  INVX1 U942 ( .A(n877), .Y(n878) );
  AND2X2 U943 ( .A(n1343), .B(n1342), .Y(n879) );
  INVX1 U944 ( .A(n879), .Y(n880) );
  AND2X2 U945 ( .A(n1356), .B(n1355), .Y(n881) );
  INVX1 U946 ( .A(n881), .Y(n882) );
  AND2X2 U947 ( .A(n1369), .B(n1368), .Y(n883) );
  INVX1 U948 ( .A(n883), .Y(n884) );
  AND2X2 U949 ( .A(n1382), .B(n1381), .Y(n885) );
  INVX1 U950 ( .A(n885), .Y(n886) );
  AND2X2 U951 ( .A(n1395), .B(n1394), .Y(n887) );
  INVX1 U952 ( .A(n887), .Y(n888) );
  AND2X2 U953 ( .A(n1485), .B(n1484), .Y(n889) );
  INVX1 U954 ( .A(n889), .Y(n890) );
  AND2X2 U955 ( .A(n1498), .B(n1497), .Y(n891) );
  INVX1 U956 ( .A(n891), .Y(n892) );
  INVX1 U957 ( .A(n1323), .Y(n893) );
  INVX1 U958 ( .A(n1324), .Y(n894) );
  INVX1 U959 ( .A(n1325), .Y(n895) );
  INVX1 U960 ( .A(n1414), .Y(n896) );
  INVX1 U961 ( .A(n1415), .Y(n897) );
  INVX1 U962 ( .A(n1416), .Y(n898) );
  INVX1 U963 ( .A(n1425), .Y(n899) );
  INVX1 U964 ( .A(n1426), .Y(n900) );
  INVX1 U965 ( .A(n1427), .Y(n901) );
  INVX1 U966 ( .A(n1436), .Y(n902) );
  INVX1 U967 ( .A(n1437), .Y(n903) );
  INVX1 U968 ( .A(n1438), .Y(n904) );
  INVX1 U969 ( .A(n1447), .Y(n905) );
  INVX1 U970 ( .A(n1448), .Y(n906) );
  INVX1 U971 ( .A(n1449), .Y(n907) );
  INVX1 U972 ( .A(n1458), .Y(n908) );
  INVX1 U973 ( .A(n1459), .Y(n909) );
  INVX1 U974 ( .A(n1460), .Y(n910) );
  INVX1 U975 ( .A(n1469), .Y(n911) );
  INVX1 U976 ( .A(n1470), .Y(n912) );
  INVX1 U977 ( .A(n1471), .Y(n913) );
  INVX1 U978 ( .A(n1480), .Y(n914) );
  INVX1 U979 ( .A(n1481), .Y(n915) );
  INVX1 U980 ( .A(n1482), .Y(n916) );
  AND2X2 U981 ( .A(n1332), .B(n1331), .Y(n917) );
  INVX1 U982 ( .A(n917), .Y(n918) );
  AND2X2 U983 ( .A(n1345), .B(n1344), .Y(n919) );
  INVX1 U984 ( .A(n919), .Y(n920) );
  AND2X2 U985 ( .A(n1358), .B(n1357), .Y(n921) );
  INVX1 U986 ( .A(n921), .Y(n922) );
  AND2X2 U987 ( .A(n1371), .B(n1370), .Y(n923) );
  INVX1 U988 ( .A(n923), .Y(n924) );
  AND2X2 U989 ( .A(n1384), .B(n1383), .Y(n925) );
  INVX1 U990 ( .A(n925), .Y(n926) );
  AND2X2 U991 ( .A(n1397), .B(n1396), .Y(n927) );
  INVX1 U992 ( .A(n927), .Y(n928) );
  AND2X2 U993 ( .A(n1487), .B(n1486), .Y(n929) );
  INVX1 U994 ( .A(n929), .Y(n930) );
  AND2X2 U995 ( .A(n1500), .B(n1499), .Y(n931) );
  INVX1 U996 ( .A(n931), .Y(n932) );
  BUFX2 U997 ( .A(n1339), .Y(n933) );
  BUFX2 U998 ( .A(n1352), .Y(n934) );
  BUFX2 U999 ( .A(n1365), .Y(n935) );
  BUFX2 U1000 ( .A(n1378), .Y(n936) );
  BUFX2 U1001 ( .A(n1391), .Y(n937) );
  BUFX2 U1002 ( .A(n1404), .Y(n938) );
  BUFX2 U1003 ( .A(n1494), .Y(n939) );
  INVX1 U1004 ( .A(n970), .Y(n940) );
  INVX1 U1005 ( .A(n1501), .Y(n941) );
  INVX1 U1006 ( .A(n1502), .Y(n942) );
  BUFX2 U1007 ( .A(n1554), .Y(n970) );
  BUFX2 U1008 ( .A(n1840), .Y(err) );
  BUFX2 U1009 ( .A(n1337), .Y(n944) );
  BUFX2 U1010 ( .A(n1350), .Y(n945) );
  BUFX2 U1011 ( .A(n1363), .Y(n946) );
  BUFX2 U1012 ( .A(n1376), .Y(n947) );
  BUFX2 U1013 ( .A(n1389), .Y(n948) );
  BUFX2 U1014 ( .A(n1402), .Y(n949) );
  BUFX2 U1015 ( .A(n1492), .Y(n950) );
  INVX1 U1016 ( .A(n971), .Y(n951) );
  INVX1 U1017 ( .A(n1503), .Y(n952) );
  INVX1 U1018 ( .A(n1504), .Y(n953) );
  BUFX2 U1019 ( .A(n1516), .Y(n971) );
  BUFX2 U1020 ( .A(n1525), .Y(n972) );
  BUFX2 U1021 ( .A(n1543), .Y(n974) );
  BUFX2 U1022 ( .A(n1553), .Y(n975) );
  BUFX2 U1023 ( .A(n1563), .Y(n976) );
  BUFX2 U1024 ( .A(n1573), .Y(n977) );
  BUFX2 U1025 ( .A(n1582), .Y(n978) );
  BUFX2 U1026 ( .A(n1592), .Y(n979) );
  BUFX2 U1027 ( .A(n1612), .Y(n982) );
  BUFX2 U1028 ( .A(n1631), .Y(n985) );
  BUFX2 U1029 ( .A(n1652), .Y(n988) );
  BUFX2 U1030 ( .A(n1672), .Y(n991) );
  BUFX2 U1031 ( .A(n1681), .Y(n992) );
  BUFX2 U1032 ( .A(n1691), .Y(n993) );
  BUFX2 U1033 ( .A(n1700), .Y(n994) );
  BUFX2 U1034 ( .A(n1710), .Y(n995) );
  BUFX2 U1035 ( .A(n1719), .Y(n996) );
  BUFX2 U1036 ( .A(n1729), .Y(n997) );
  BUFX2 U1037 ( .A(n1738), .Y(n998) );
  BUFX2 U1038 ( .A(n1748), .Y(n999) );
  BUFX2 U1039 ( .A(n1767), .Y(n1002) );
  BUFX2 U1040 ( .A(n1787), .Y(n1005) );
  BUFX2 U1041 ( .A(n1807), .Y(n1008) );
  BUFX2 U1042 ( .A(n1820), .Y(n973) );
  AND2X1 U1043 ( .A(n1632), .B(n1320), .Y(n1819) );
  BUFX2 U1044 ( .A(n1839), .Y(n1011) );
  BUFX2 U1045 ( .A(n1602), .Y(n954) );
  BUFX2 U1046 ( .A(n1621), .Y(n955) );
  BUFX2 U1047 ( .A(n1642), .Y(n956) );
  BUFX2 U1048 ( .A(n1662), .Y(n957) );
  BUFX2 U1049 ( .A(n1757), .Y(n958) );
  BUFX2 U1050 ( .A(n1777), .Y(n959) );
  BUFX2 U1051 ( .A(n1797), .Y(n960) );
  BUFX2 U1052 ( .A(n1818), .Y(n961) );
  AND2X1 U1053 ( .A(enable), .B(n1015), .Y(n962) );
  INVX1 U1054 ( .A(n962), .Y(n963) );
  INVX1 U1055 ( .A(n965), .Y(n964) );
  AND2X1 U1056 ( .A(n1515), .B(n1514), .Y(n965) );
  INVX1 U1057 ( .A(n966), .Y(n967) );
  INVX1 U1058 ( .A(n968), .Y(n969) );
  AND2X1 U1059 ( .A(n951), .B(n1312), .Y(n1526) );
endmodule


module dff_212 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_213 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_214 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_215 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_208 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_209 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_210 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_211 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_204 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_205 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_206 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_207 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module cache_cache_id0 ( enable, clk, rst, createdump, .tag_in({\tag_in<4> , 
        \tag_in<3> , \tag_in<2> , \tag_in<1> , \tag_in<0> }), .index({
        \index<7> , \index<6> , \index<5> , \index<4> , \index<3> , \index<2> , 
        \index<1> , \index<0> }), .offset({\offset<2> , \offset<1> , 
        \offset<0> }), .data_in({\data_in<15> , \data_in<14> , \data_in<13> , 
        \data_in<12> , \data_in<11> , \data_in<10> , \data_in<9> , 
        \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , 
        \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), comp, write, 
        valid_in, .tag_out({\tag_out<4> , \tag_out<3> , \tag_out<2> , 
        \tag_out<1> , \tag_out<0> }), .data_out({\data_out<15> , 
        \data_out<14> , \data_out<13> , \data_out<12> , \data_out<11> , 
        \data_out<10> , \data_out<9> , \data_out<8> , \data_out<7> , 
        \data_out<6> , \data_out<5> , \data_out<4> , \data_out<3> , 
        \data_out<2> , \data_out<1> , \data_out<0> }), hit, dirty, valid, err
 );
  input enable, clk, rst, createdump, \tag_in<4> , \tag_in<3> , \tag_in<2> ,
         \tag_in<1> , \tag_in<0> , \index<7> , \index<6> , \index<5> ,
         \index<4> , \index<3> , \index<2> , \index<1> , \index<0> ,
         \offset<2> , \offset<1> , \offset<0> , \data_in<15> , \data_in<14> ,
         \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> ,
         \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> ,
         \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> ,
         comp, write, valid_in;
  output \tag_out<4> , \tag_out<3> , \tag_out<2> , \tag_out<1> , \tag_out<0> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , hit,
         dirty, valid, err;
  wire   n197, n198, n199, n200, n201, \w0<15> , \w0<14> , \w0<13> , \w0<12> ,
         \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> ,
         \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> , \w1<15> , \w1<14> ,
         \w1<13> , \w1<12> , \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> ,
         \w1<6> , \w1<5> , \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> ,
         \w2<15> , \w2<14> , \w2<13> , \w2<12> , \w2<11> , \w2<10> , \w2<9> ,
         \w2<8> , \w2<7> , \w2<6> , \w2<5> , \w2<4> , \w2<3> , \w2<2> ,
         \w2<1> , \w2<0> , \w3<15> , \w3<14> , \w3<13> , \w3<12> , \w3<11> ,
         \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , \w3<4> ,
         \w3<3> , \w3<2> , \w3<1> , \w3<0> , dirtybit, validbit, n1, n3, n4,
         n5, n6, n7, n8, n9, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n29, n31, n33, n35, n37, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n83, n85,
         n87, n89, n91, n93, n95, n97, n99, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n124, n125, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195;

  memc_Size16_3 mem_w0 ( .data_out({\w0<15> , \w0<14> , \w0<13> , \w0<12> , 
        \w0<11> , \w0<10> , \w0<9> , \w0<8> , \w0<7> , \w0<6> , \w0<5> , 
        \w0<4> , \w0<3> , \w0<2> , \w0<1> , \w0<0> }), .addr({\index<7> , 
        \index<6> , \index<5> , n144, n142, n140, n8, n6}), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), .write(n21), .clk(clk), .rst(n136), 
        .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  memc_Size16_2 mem_w1 ( .data_out({\w1<15> , \w1<14> , \w1<13> , \w1<12> , 
        \w1<11> , \w1<10> , \w1<9> , \w1<8> , \w1<7> , \w1<6> , \w1<5> , 
        \w1<4> , \w1<3> , \w1<2> , \w1<1> , \w1<0> }), .addr({\index<7> , 
        \index<6> , \index<5> , n144, n142, n140, n8, n6}), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), .write(n121), .clk(clk), .rst(n136), 
        .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b0, 1'b1}) );
  memc_Size16_1 mem_w2 ( .data_out({\w2<15> , \w2<14> , \w2<13> , \w2<12> , 
        \w2<11> , \w2<10> , \w2<9> , \w2<8> , \w2<7> , \w2<6> , \w2<5> , 
        \w2<4> , \w2<3> , \w2<2> , \w2<1> , \w2<0> }), .addr({\index<7> , 
        \index<6> , \index<5> , n144, n142, n140, n8, n6}), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), .write(n19), .clk(clk), .rst(n136), 
        .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b1, 1'b0}) );
  memc_Size16_0 mem_w3 ( .data_out({\w3<15> , \w3<14> , \w3<13> , \w3<12> , 
        \w3<11> , \w3<10> , \w3<9> , \w3<8> , \w3<7> , \w3<6> , \w3<5> , 
        \w3<4> , \w3<3> , \w3<2> , \w3<1> , \w3<0> }), .addr({\index<7> , 
        \index<6> , \index<5> , n144, n142, n140, n8, n6}), .data_in({
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), .write(n120), .clk(clk), .rst(n136), 
        .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b1, 1'b1}) );
  memc_Size5 mem_tg ( .data_out({n197, n198, n199, n200, n201}), .addr({
        \index<7> , \index<6> , \index<5> , n144, n142, n140, n138, n129}), 
        .data_in({\tag_in<4> , \tag_in<3> , \tag_in<2> , \tag_in<1> , 
        \tag_in<0> }), .write(n17), .clk(clk), .rst(n136), .createdump(
        createdump), .file_id({1'b0, 1'b0, 1'b1, 1'b0, 1'b0}) );
  memc_Size1 mem_dr ( .data_out(dirtybit), .addr({\index<7> , \index<6> , 
        \index<5> , n144, n142, n140, n138, n6}), .data_in(n16), .write(n134), 
        .clk(clk), .rst(n136), .createdump(createdump), .file_id({1'b0, 1'b0, 
        1'b1, 1'b0, 1'b1}) );
  memv mem_vl ( .data_out(validbit), .addr({\index<7> , \index<6> , \index<5> , 
        n144, n142, n140, n8, n6}), .data_in(valid_in), .write(n132), .clk(clk), .rst(n136), .createdump(createdump), .file_id({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}) );
  BUFX2 U3 ( .A(n129), .Y(n1) );
  XOR2X1 U4 ( .A(n198), .B(\tag_in<3> ), .Y(n146) );
  BUFX2 U5 ( .A(n200), .Y(\tag_out<1> ) );
  AND2X2 U6 ( .A(n62), .B(n50), .Y(n75) );
  BUFX2 U7 ( .A(n192), .Y(n135) );
  INVX1 U8 ( .A(n119), .Y(n158) );
  INVX2 U9 ( .A(n102), .Y(n191) );
  INVX1 U10 ( .A(\index<4> ), .Y(n145) );
  INVX2 U11 ( .A(rst), .Y(n137) );
  INVX1 U12 ( .A(\offset<0> ), .Y(n125) );
  INVX1 U13 ( .A(n125), .Y(err) );
  INVX1 U14 ( .A(n22), .Y(n3) );
  XOR2X1 U15 ( .A(n201), .B(\tag_in<0> ), .Y(n148) );
  XOR2X1 U16 ( .A(n199), .B(\tag_in<2> ), .Y(n147) );
  OR2X1 U17 ( .A(n124), .B(n133), .Y(n159) );
  BUFX2 U18 ( .A(n23), .Y(n4) );
  INVX1 U19 ( .A(n1), .Y(n5) );
  INVX1 U20 ( .A(n5), .Y(n6) );
  INVX1 U21 ( .A(n138), .Y(n7) );
  INVX1 U22 ( .A(n7), .Y(n8) );
  XOR2X1 U23 ( .A(n200), .B(\tag_in<1> ), .Y(n149) );
  BUFX2 U24 ( .A(n150), .Y(n9) );
  BUFX2 U25 ( .A(n197), .Y(\tag_out<4> ) );
  OAI21X1 U26 ( .A(n152), .B(n112), .C(n26), .Y(n11) );
  INVX1 U27 ( .A(n133), .Y(n152) );
  BUFX2 U28 ( .A(n201), .Y(\tag_out<0> ) );
  BUFX2 U29 ( .A(n101), .Y(n13) );
  BUFX2 U30 ( .A(n151), .Y(n14) );
  INVX1 U31 ( .A(n22), .Y(n15) );
  INVX1 U32 ( .A(n14), .Y(n16) );
  AND2X2 U33 ( .A(n101), .B(n23), .Y(n17) );
  AND2X2 U34 ( .A(n150), .B(n4), .Y(n22) );
  OR2X2 U35 ( .A(n154), .B(n108), .Y(n18) );
  INVX1 U36 ( .A(n18), .Y(n19) );
  OR2X2 U37 ( .A(n154), .B(n111), .Y(n20) );
  INVX1 U38 ( .A(n20), .Y(n21) );
  AND2X2 U39 ( .A(enable), .B(n137), .Y(n23) );
  OR2X2 U40 ( .A(n154), .B(n119), .Y(n24) );
  OR2X2 U41 ( .A(n154), .B(n110), .Y(n25) );
  AND2X2 U42 ( .A(n4), .B(dirtybit), .Y(n26) );
  AND2X2 U43 ( .A(n69), .B(n63), .Y(n27) );
  INVX1 U44 ( .A(n27), .Y(\data_out<0> ) );
  AND2X2 U45 ( .A(n64), .B(n70), .Y(n29) );
  INVX1 U46 ( .A(n29), .Y(\data_out<1> ) );
  AND2X2 U47 ( .A(n71), .B(n65), .Y(n31) );
  INVX1 U48 ( .A(n31), .Y(\data_out<2> ) );
  AND2X2 U49 ( .A(n66), .B(n72), .Y(n33) );
  INVX1 U50 ( .A(n33), .Y(\data_out<3> ) );
  AND2X2 U51 ( .A(n67), .B(n73), .Y(n35) );
  INVX1 U52 ( .A(n35), .Y(\data_out<12> ) );
  AND2X2 U53 ( .A(n74), .B(n68), .Y(n37) );
  INVX1 U54 ( .A(n37), .Y(\data_out<15> ) );
  BUFX2 U55 ( .A(n170), .Y(n39) );
  BUFX2 U56 ( .A(n172), .Y(n40) );
  BUFX2 U57 ( .A(n174), .Y(n41) );
  BUFX2 U58 ( .A(n176), .Y(n42) );
  BUFX2 U59 ( .A(n178), .Y(n43) );
  BUFX2 U60 ( .A(n180), .Y(n44) );
  BUFX2 U61 ( .A(n182), .Y(n45) );
  BUFX2 U62 ( .A(n184), .Y(n46) );
  BUFX2 U63 ( .A(n188), .Y(n47) );
  BUFX2 U64 ( .A(n190), .Y(n48) );
  AND2X2 U65 ( .A(n197), .B(\tag_in<4> ), .Y(n49) );
  INVX1 U66 ( .A(n49), .Y(n50) );
  BUFX2 U67 ( .A(n169), .Y(n51) );
  BUFX2 U68 ( .A(n171), .Y(n52) );
  BUFX2 U69 ( .A(n173), .Y(n53) );
  BUFX2 U70 ( .A(n175), .Y(n54) );
  BUFX2 U71 ( .A(n177), .Y(n55) );
  BUFX2 U72 ( .A(n179), .Y(n56) );
  BUFX2 U73 ( .A(n181), .Y(n57) );
  BUFX2 U74 ( .A(n183), .Y(n58) );
  BUFX2 U75 ( .A(n187), .Y(n59) );
  BUFX2 U76 ( .A(n189), .Y(n60) );
  AND2X2 U77 ( .A(n130), .B(n131), .Y(n61) );
  INVX1 U78 ( .A(n61), .Y(n62) );
  BUFX2 U79 ( .A(n161), .Y(n63) );
  BUFX2 U80 ( .A(n163), .Y(n64) );
  BUFX2 U81 ( .A(n165), .Y(n65) );
  BUFX2 U82 ( .A(n167), .Y(n66) );
  BUFX2 U83 ( .A(n186), .Y(n67) );
  BUFX2 U84 ( .A(n193), .Y(n68) );
  BUFX2 U85 ( .A(n162), .Y(n69) );
  BUFX2 U86 ( .A(n164), .Y(n70) );
  BUFX2 U87 ( .A(n166), .Y(n71) );
  BUFX2 U88 ( .A(n168), .Y(n72) );
  BUFX2 U89 ( .A(n185), .Y(n73) );
  BUFX2 U90 ( .A(n194), .Y(n74) );
  INVX1 U91 ( .A(n75), .Y(n76) );
  OR2X2 U92 ( .A(n147), .B(n146), .Y(n77) );
  INVX1 U93 ( .A(n77), .Y(n78) );
  OR2X2 U94 ( .A(n149), .B(n148), .Y(n79) );
  INVX1 U95 ( .A(n79), .Y(n80) );
  AND2X2 U96 ( .A(n51), .B(n39), .Y(n81) );
  INVX1 U97 ( .A(n81), .Y(\data_out<4> ) );
  AND2X2 U98 ( .A(n40), .B(n52), .Y(n83) );
  INVX1 U99 ( .A(n83), .Y(\data_out<5> ) );
  AND2X2 U100 ( .A(n54), .B(n42), .Y(n85) );
  INVX1 U101 ( .A(n85), .Y(\data_out<7> ) );
  AND2X2 U102 ( .A(n43), .B(n55), .Y(n87) );
  INVX1 U103 ( .A(n87), .Y(\data_out<8> ) );
  AND2X2 U104 ( .A(n45), .B(n57), .Y(n89) );
  INVX1 U105 ( .A(n89), .Y(\data_out<10> ) );
  AND2X2 U106 ( .A(n46), .B(n58), .Y(n91) );
  INVX1 U107 ( .A(n91), .Y(\data_out<11> ) );
  AND2X2 U108 ( .A(n47), .B(n59), .Y(n93) );
  INVX1 U109 ( .A(n93), .Y(\data_out<13> ) );
  AND2X2 U110 ( .A(n48), .B(n60), .Y(n95) );
  INVX1 U111 ( .A(n95), .Y(\data_out<14> ) );
  AND2X2 U112 ( .A(n41), .B(n53), .Y(n97) );
  INVX1 U113 ( .A(n97), .Y(\data_out<6> ) );
  AND2X2 U114 ( .A(n56), .B(n44), .Y(n99) );
  INVX1 U115 ( .A(n99), .Y(\data_out<9> ) );
  AND2X2 U116 ( .A(n151), .B(write), .Y(n101) );
  INVX1 U117 ( .A(comp), .Y(n151) );
  OR2X1 U118 ( .A(n114), .B(n103), .Y(n102) );
  OR2X1 U119 ( .A(n113), .B(n159), .Y(n103) );
  OR2X1 U120 ( .A(n157), .B(n106), .Y(n104) );
  INVX1 U121 ( .A(n104), .Y(n105) );
  OR2X1 U122 ( .A(n115), .B(n159), .Y(n106) );
  AND2X2 U123 ( .A(\offset<2> ), .B(n157), .Y(n107) );
  INVX1 U124 ( .A(n107), .Y(n108) );
  AND2X2 U125 ( .A(n114), .B(\offset<1> ), .Y(n109) );
  INVX1 U126 ( .A(n109), .Y(n110) );
  OR2X2 U127 ( .A(\offset<1> ), .B(\offset<2> ), .Y(n111) );
  AND2X1 U128 ( .A(n16), .B(n117), .Y(n112) );
  INVX1 U129 ( .A(n157), .Y(n113) );
  INVX1 U130 ( .A(\offset<2> ), .Y(n114) );
  INVX1 U131 ( .A(\offset<1> ), .Y(n157) );
  INVX1 U132 ( .A(n114), .Y(n115) );
  INVX1 U133 ( .A(n159), .Y(n160) );
  AND2X1 U134 ( .A(n158), .B(n160), .Y(n116) );
  INVX1 U135 ( .A(n9), .Y(n117) );
  AND2X2 U136 ( .A(\offset<2> ), .B(\offset<1> ), .Y(n118) );
  INVX1 U137 ( .A(n118), .Y(n119) );
  INVX1 U138 ( .A(n24), .Y(n120) );
  INVX1 U139 ( .A(n25), .Y(n121) );
  INVX1 U140 ( .A(n22), .Y(n122) );
  INVX1 U141 ( .A(n11), .Y(dirty) );
  INVX1 U142 ( .A(n4), .Y(n124) );
  INVX4 U143 ( .A(n139), .Y(n138) );
  INVX1 U144 ( .A(\index<1> ), .Y(n139) );
  BUFX2 U145 ( .A(n198), .Y(\tag_out<3> ) );
  BUFX2 U146 ( .A(n199), .Y(\tag_out<2> ) );
  BUFX4 U147 ( .A(\index<0> ), .Y(n129) );
  INVX1 U148 ( .A(\tag_in<4> ), .Y(n130) );
  INVX1 U149 ( .A(n197), .Y(n131) );
  BUFX2 U150 ( .A(n17), .Y(n132) );
  BUFX2 U151 ( .A(write), .Y(n133) );
  INVX1 U152 ( .A(n132), .Y(n153) );
  INVX1 U153 ( .A(n122), .Y(hit) );
  OAI21X1 U154 ( .A(n15), .B(n152), .C(n153), .Y(n134) );
  INVX1 U155 ( .A(n156), .Y(n150) );
  INVX8 U156 ( .A(n137), .Y(n136) );
  INVX8 U157 ( .A(n141), .Y(n140) );
  INVX8 U158 ( .A(\index<2> ), .Y(n141) );
  INVX8 U159 ( .A(n143), .Y(n142) );
  INVX8 U160 ( .A(\index<3> ), .Y(n143) );
  INVX8 U161 ( .A(n145), .Y(n144) );
  NAND3X1 U162 ( .A(n76), .B(n78), .C(n80), .Y(n156) );
  OAI21X1 U163 ( .A(n152), .B(n3), .C(n153), .Y(n195) );
  INVX2 U164 ( .A(n195), .Y(n154) );
  INVX2 U165 ( .A(validbit), .Y(n155) );
  NOR3X1 U166 ( .A(n13), .B(n124), .C(n155), .Y(valid) );
  AOI22X1 U167 ( .A(n191), .B(\w2<0> ), .C(n116), .D(\w3<0> ), .Y(n162) );
  NOR3X1 U168 ( .A(\offset<2> ), .B(n159), .C(\offset<1> ), .Y(n192) );
  AOI22X1 U169 ( .A(n135), .B(\w0<0> ), .C(\w1<0> ), .D(n105), .Y(n161) );
  AOI22X1 U170 ( .A(n191), .B(\w2<1> ), .C(n116), .D(\w3<1> ), .Y(n164) );
  AOI22X1 U171 ( .A(n135), .B(\w0<1> ), .C(\w1<1> ), .D(n105), .Y(n163) );
  AOI22X1 U172 ( .A(n191), .B(\w2<2> ), .C(n116), .D(\w3<2> ), .Y(n166) );
  AOI22X1 U173 ( .A(n135), .B(\w0<2> ), .C(n105), .D(\w1<2> ), .Y(n165) );
  AOI22X1 U174 ( .A(n191), .B(\w2<3> ), .C(n116), .D(\w3<3> ), .Y(n168) );
  AOI22X1 U175 ( .A(n135), .B(\w0<3> ), .C(n105), .D(\w1<3> ), .Y(n167) );
  AOI22X1 U176 ( .A(n191), .B(\w2<4> ), .C(n116), .D(\w3<4> ), .Y(n170) );
  AOI22X1 U177 ( .A(n135), .B(\w0<4> ), .C(n105), .D(\w1<4> ), .Y(n169) );
  AOI22X1 U178 ( .A(n191), .B(\w2<5> ), .C(n116), .D(\w3<5> ), .Y(n172) );
  AOI22X1 U179 ( .A(n135), .B(\w0<5> ), .C(\w1<5> ), .D(n105), .Y(n171) );
  AOI22X1 U180 ( .A(n191), .B(\w2<6> ), .C(n116), .D(\w3<6> ), .Y(n174) );
  AOI22X1 U181 ( .A(n135), .B(\w0<6> ), .C(\w1<6> ), .D(n105), .Y(n173) );
  AOI22X1 U182 ( .A(n191), .B(\w2<7> ), .C(n116), .D(\w3<7> ), .Y(n176) );
  AOI22X1 U183 ( .A(n135), .B(\w0<7> ), .C(n105), .D(\w1<7> ), .Y(n175) );
  AOI22X1 U184 ( .A(n191), .B(\w2<8> ), .C(n116), .D(\w3<8> ), .Y(n178) );
  AOI22X1 U185 ( .A(n135), .B(\w0<8> ), .C(\w1<8> ), .D(n105), .Y(n177) );
  AOI22X1 U186 ( .A(n191), .B(\w2<9> ), .C(n116), .D(\w3<9> ), .Y(n180) );
  AOI22X1 U187 ( .A(n135), .B(\w0<9> ), .C(n105), .D(\w1<9> ), .Y(n179) );
  AOI22X1 U188 ( .A(n191), .B(\w2<10> ), .C(n116), .D(\w3<10> ), .Y(n182) );
  AOI22X1 U189 ( .A(n135), .B(\w0<10> ), .C(\w1<10> ), .D(n105), .Y(n181) );
  AOI22X1 U190 ( .A(n191), .B(\w2<11> ), .C(n116), .D(\w3<11> ), .Y(n184) );
  AOI22X1 U191 ( .A(n135), .B(\w0<11> ), .C(\w1<11> ), .D(n105), .Y(n183) );
  AOI22X1 U192 ( .A(n191), .B(\w2<12> ), .C(n116), .D(\w3<12> ), .Y(n186) );
  AOI22X1 U193 ( .A(n135), .B(\w0<12> ), .C(\w1<12> ), .D(n105), .Y(n185) );
  AOI22X1 U194 ( .A(n191), .B(\w2<13> ), .C(n116), .D(\w3<13> ), .Y(n188) );
  AOI22X1 U195 ( .A(n135), .B(\w0<13> ), .C(\w1<13> ), .D(n105), .Y(n187) );
  AOI22X1 U196 ( .A(n191), .B(\w2<14> ), .C(n116), .D(\w3<14> ), .Y(n190) );
  AOI22X1 U197 ( .A(n135), .B(\w0<14> ), .C(n105), .D(\w1<14> ), .Y(n189) );
  AOI22X1 U198 ( .A(n191), .B(\w2<15> ), .C(n116), .D(\w3<15> ), .Y(n194) );
  AOI22X1 U199 ( .A(n135), .B(\w0<15> ), .C(\w1<15> ), .D(n105), .Y(n193) );
endmodule


module four_bank_mem ( clk, rst, createdump, .addr({\addr<15> , \addr<14> , 
        \addr<13> , \addr<12> , \addr<11> , \addr<10> , \addr<9> , \addr<8> , 
        \addr<7> , \addr<6> , \addr<5> , \addr<4> , \addr<3> , \addr<2> , 
        \addr<1> , \addr<0> }), .data_in({\data_in<15> , \data_in<14> , 
        \data_in<13> , \data_in<12> , \data_in<11> , \data_in<10> , 
        \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , \data_in<5> , 
        \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> }), 
        wr, rd, .data_out({\data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), stall, .busy({\busy<3> , \busy<2> , \busy<1> , 
        \busy<0> }), err );
  input clk, rst, createdump, \addr<15> , \addr<14> , \addr<13> , \addr<12> ,
         \addr<11> , \addr<10> , \addr<9> , \addr<8> , \addr<7> , \addr<6> ,
         \addr<5> , \addr<4> , \addr<3> , \addr<2> , \addr<1> , \addr<0> ,
         \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , wr, rd;
  output \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> , stall,
         \busy<3> , \busy<2> , \busy<1> , \busy<0> , err;
  wire   \en<3> , \en<2> , \en<1> , \en<0> , \data0_out<15> , \data0_out<14> ,
         \data0_out<13> , \data0_out<12> , \data0_out<11> , \data0_out<10> ,
         \data0_out<9> , \data0_out<8> , \data0_out<7> , \data0_out<6> ,
         \data0_out<5> , \data0_out<4> , \data0_out<3> , \data0_out<2> ,
         \data0_out<1> , \data0_out<0> , err0, \data1_out<15> ,
         \data1_out<14> , \data1_out<13> , \data1_out<12> , \data1_out<11> ,
         \data1_out<10> , \data1_out<9> , \data1_out<8> , \data1_out<7> ,
         \data1_out<6> , \data1_out<5> , \data1_out<4> , \data1_out<3> ,
         \data1_out<2> , \data1_out<1> , \data1_out<0> , err1, \data2_out<15> ,
         \data2_out<14> , \data2_out<13> , \data2_out<12> , \data2_out<11> ,
         \data2_out<10> , \data2_out<9> , \data2_out<8> , \data2_out<7> ,
         \data2_out<6> , \data2_out<5> , \data2_out<4> , \data2_out<3> ,
         \data2_out<2> , \data2_out<1> , \data2_out<0> , err2, \data3_out<15> ,
         \data3_out<14> , \data3_out<13> , \data3_out<12> , \data3_out<11> ,
         \data3_out<10> , \data3_out<9> , \data3_out<8> , \data3_out<7> ,
         \data3_out<6> , \data3_out<5> , \data3_out<4> , \data3_out<3> ,
         \data3_out<2> , \data3_out<1> , \data3_out<0> , err3, \bsy0<3> ,
         \bsy0<2> , \bsy0<1> , \bsy0<0> , \bsy1<3> , \bsy1<2> , \bsy1<1> ,
         \bsy1<0> , \bsy2<3> , \bsy2<2> , \bsy2<1> , \bsy2<0> , n9, n10, n11,
         n13, n16, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n1, n2, n3, n4, n5, n6, n7,
         n8, n12, n14, n15, n17, n18, n19, n21, n55, n56, n57, n58, n59, n61,
         n63, n65, n67, n69, n71, n73, n75, n77, n79, n81, n83, n85, n87, n89,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106;

  NOR3X1 U9 ( .A(n92), .B(n93), .C(n5), .Y(stall) );
  OAI21X1 U11 ( .A(\addr<1> ), .B(n11), .C(n12), .Y(n10) );
  OAI21X1 U13 ( .A(\addr<1> ), .B(n13), .C(n8), .Y(n9) );
  AOI21X1 U15 ( .A(n15), .B(n16), .C(n92), .Y(err) );
  NOR3X1 U16 ( .A(err1), .B(err3), .C(err2), .Y(n16) );
  NOR3X1 U18 ( .A(n58), .B(\busy<3> ), .C(n92), .Y(\en<3> ) );
  NOR3X1 U20 ( .A(n56), .B(n92), .C(n106), .Y(\en<2> ) );
  NOR3X1 U22 ( .A(n21), .B(n92), .C(n105), .Y(\en<1> ) );
  NOR3X1 U24 ( .A(n18), .B(\busy<0> ), .C(n92), .Y(\en<0> ) );
  NOR2X1 U28 ( .A(\data3_out<9> ), .B(\data2_out<9> ), .Y(n23) );
  NOR2X1 U29 ( .A(\data1_out<9> ), .B(\data0_out<9> ), .Y(n22) );
  NOR2X1 U31 ( .A(\data3_out<8> ), .B(\data2_out<8> ), .Y(n25) );
  NOR2X1 U32 ( .A(\data1_out<8> ), .B(\data0_out<8> ), .Y(n24) );
  NOR2X1 U34 ( .A(\data3_out<7> ), .B(\data2_out<7> ), .Y(n27) );
  NOR2X1 U35 ( .A(\data1_out<7> ), .B(\data0_out<7> ), .Y(n26) );
  NOR2X1 U37 ( .A(\data3_out<6> ), .B(\data2_out<6> ), .Y(n29) );
  NOR2X1 U38 ( .A(\data1_out<6> ), .B(\data0_out<6> ), .Y(n28) );
  NOR2X1 U40 ( .A(\data3_out<5> ), .B(\data2_out<5> ), .Y(n31) );
  NOR2X1 U41 ( .A(\data1_out<5> ), .B(\data0_out<5> ), .Y(n30) );
  NOR2X1 U43 ( .A(\data3_out<4> ), .B(\data2_out<4> ), .Y(n33) );
  NOR2X1 U44 ( .A(\data1_out<4> ), .B(\data0_out<4> ), .Y(n32) );
  NOR2X1 U46 ( .A(\data3_out<3> ), .B(\data2_out<3> ), .Y(n35) );
  NOR2X1 U47 ( .A(\data1_out<3> ), .B(\data0_out<3> ), .Y(n34) );
  NOR2X1 U49 ( .A(\data3_out<2> ), .B(\data2_out<2> ), .Y(n37) );
  NOR2X1 U50 ( .A(\data1_out<2> ), .B(\data0_out<2> ), .Y(n36) );
  NOR2X1 U52 ( .A(\data3_out<1> ), .B(\data2_out<1> ), .Y(n39) );
  NOR2X1 U53 ( .A(\data1_out<1> ), .B(\data0_out<1> ), .Y(n38) );
  NOR2X1 U55 ( .A(\data3_out<15> ), .B(\data2_out<15> ), .Y(n41) );
  NOR2X1 U56 ( .A(\data1_out<15> ), .B(\data0_out<15> ), .Y(n40) );
  NOR2X1 U58 ( .A(\data3_out<14> ), .B(\data2_out<14> ), .Y(n43) );
  NOR2X1 U59 ( .A(\data1_out<14> ), .B(\data0_out<14> ), .Y(n42) );
  NOR2X1 U61 ( .A(\data3_out<13> ), .B(\data2_out<13> ), .Y(n45) );
  NOR2X1 U62 ( .A(\data1_out<13> ), .B(\data0_out<13> ), .Y(n44) );
  NOR2X1 U64 ( .A(\data3_out<12> ), .B(\data2_out<12> ), .Y(n47) );
  NOR2X1 U65 ( .A(\data1_out<12> ), .B(\data0_out<12> ), .Y(n46) );
  NOR2X1 U67 ( .A(\data3_out<11> ), .B(\data2_out<11> ), .Y(n49) );
  NOR2X1 U68 ( .A(\data1_out<11> ), .B(\data0_out<11> ), .Y(n48) );
  NOR2X1 U70 ( .A(\data3_out<10> ), .B(\data2_out<10> ), .Y(n51) );
  NOR2X1 U71 ( .A(\data1_out<10> ), .B(\data0_out<10> ), .Y(n50) );
  NOR2X1 U73 ( .A(\data3_out<0> ), .B(\data2_out<0> ), .Y(n53) );
  NOR2X1 U74 ( .A(\data1_out<0> ), .B(\data0_out<0> ), .Y(n52) );
  NOR3X1 U75 ( .A(\bsy0<3> ), .B(\bsy2<3> ), .C(\bsy1<3> ), .Y(n54) );
  NOR3X1 U76 ( .A(\bsy0<2> ), .B(\bsy2<2> ), .C(\bsy1<2> ), .Y(n11) );
  NOR3X1 U77 ( .A(\bsy0<1> ), .B(\bsy2<1> ), .C(\bsy1<1> ), .Y(n20) );
  NOR3X1 U78 ( .A(\bsy0<0> ), .B(\bsy2<0> ), .C(\bsy1<0> ), .Y(n13) );
  final_memory_3 m0 ( .data_out({\data0_out<15> , \data0_out<14> , 
        \data0_out<13> , \data0_out<12> , \data0_out<11> , \data0_out<10> , 
        \data0_out<9> , \data0_out<8> , \data0_out<7> , \data0_out<6> , 
        \data0_out<5> , \data0_out<4> , \data0_out<3> , \data0_out<2> , 
        \data0_out<1> , \data0_out<0> }), .err(err0), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , n103, n101, n99, n97, 
        n95}), .wr(wr), .rd(rd), .enable(\en<0> ), .create_dump(createdump), 
        .bank_id({1'b0, 1'b0}), .clk(clk), .rst(n93) );
  final_memory_2 m1 ( .data_out({\data1_out<15> , \data1_out<14> , 
        \data1_out<13> , \data1_out<12> , \data1_out<11> , \data1_out<10> , 
        \data1_out<9> , \data1_out<8> , \data1_out<7> , \data1_out<6> , 
        \data1_out<5> , \data1_out<4> , \data1_out<3> , \data1_out<2> , 
        \data1_out<1> , \data1_out<0> }), .err(err1), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , n103, n101, n99, n97, 
        n95}), .wr(wr), .rd(rd), .enable(\en<1> ), .create_dump(createdump), 
        .bank_id({1'b0, 1'b1}), .clk(clk), .rst(n93) );
  final_memory_1 m2 ( .data_out({\data2_out<15> , \data2_out<14> , 
        \data2_out<13> , \data2_out<12> , \data2_out<11> , \data2_out<10> , 
        \data2_out<9> , \data2_out<8> , \data2_out<7> , \data2_out<6> , 
        \data2_out<5> , \data2_out<4> , \data2_out<3> , \data2_out<2> , 
        \data2_out<1> , \data2_out<0> }), .err(err2), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , n103, n101, n99, n97, 
        n95}), .wr(wr), .rd(rd), .enable(\en<2> ), .create_dump(createdump), 
        .bank_id({1'b1, 1'b0}), .clk(clk), .rst(n93) );
  final_memory_0 m3 ( .data_out({\data3_out<15> , \data3_out<14> , 
        \data3_out<13> , \data3_out<12> , \data3_out<11> , \data3_out<10> , 
        \data3_out<9> , \data3_out<8> , \data3_out<7> , \data3_out<6> , 
        \data3_out<5> , \data3_out<4> , \data3_out<3> , \data3_out<2> , 
        \data3_out<1> , \data3_out<0> }), .err(err3), .data_in({\data_in<15> , 
        \data_in<14> , \data_in<13> , \data_in<12> , \data_in<11> , 
        \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , \data_in<6> , 
        \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , 
        \data_in<0> }), .addr({\addr<15> , \addr<14> , \addr<13> , \addr<12> , 
        \addr<11> , \addr<10> , \addr<9> , \addr<8> , n103, n101, n99, n97, 
        n95}), .wr(wr), .rd(rd), .enable(\en<3> ), .create_dump(createdump), 
        .bank_id({1'b1, 1'b1}), .clk(clk), .rst(n93) );
  dff_212 \b0[0]  ( .q(\bsy0<0> ), .d(\en<0> ), .clk(clk), .rst(n93) );
  dff_213 \b0[1]  ( .q(\bsy0<1> ), .d(\en<1> ), .clk(clk), .rst(n93) );
  dff_214 \b0[2]  ( .q(\bsy0<2> ), .d(\en<2> ), .clk(clk), .rst(n93) );
  dff_215 \b0[3]  ( .q(\bsy0<3> ), .d(\en<3> ), .clk(clk), .rst(n93) );
  dff_208 \b1[0]  ( .q(\bsy1<0> ), .d(\bsy0<0> ), .clk(clk), .rst(n93) );
  dff_209 \b1[1]  ( .q(\bsy1<1> ), .d(\bsy0<1> ), .clk(clk), .rst(n93) );
  dff_210 \b1[2]  ( .q(\bsy1<2> ), .d(\bsy0<2> ), .clk(clk), .rst(n93) );
  dff_211 \b1[3]  ( .q(\bsy1<3> ), .d(\bsy0<3> ), .clk(clk), .rst(n93) );
  dff_204 \b2[0]  ( .q(\bsy2<0> ), .d(\bsy1<0> ), .clk(clk), .rst(n93) );
  dff_205 \b2[1]  ( .q(\bsy2<1> ), .d(\bsy1<1> ), .clk(clk), .rst(n93) );
  dff_206 \b2[2]  ( .q(\bsy2<2> ), .d(\bsy1<2> ), .clk(clk), .rst(n93) );
  dff_207 \b2[3]  ( .q(\bsy2<3> ), .d(\bsy1<3> ), .clk(clk), .rst(n93) );
  INVX1 U3 ( .A(n13), .Y(\busy<0> ) );
  INVX1 U4 ( .A(n20), .Y(\busy<1> ) );
  INVX1 U5 ( .A(n54), .Y(\busy<3> ) );
  INVX1 U6 ( .A(n96), .Y(n95) );
  INVX1 U7 ( .A(n98), .Y(n97) );
  INVX1 U8 ( .A(n100), .Y(n99) );
  INVX1 U10 ( .A(\addr<5> ), .Y(n100) );
  INVX1 U12 ( .A(n102), .Y(n101) );
  INVX1 U14 ( .A(\addr<6> ), .Y(n102) );
  INVX1 U17 ( .A(n104), .Y(n103) );
  INVX1 U19 ( .A(\addr<7> ), .Y(n104) );
  OR2X1 U21 ( .A(rd), .B(wr), .Y(n91) );
  INVX1 U23 ( .A(rst), .Y(n94) );
  OR2X1 U25 ( .A(err0), .B(\addr<0> ), .Y(n14) );
  INVX1 U26 ( .A(n11), .Y(\busy<2> ) );
  INVX2 U27 ( .A(\addr<2> ), .Y(n106) );
  AND2X2 U30 ( .A(n9), .B(n106), .Y(n1) );
  INVX1 U33 ( .A(n1), .Y(n2) );
  AND2X2 U36 ( .A(n10), .B(\addr<2> ), .Y(n3) );
  INVX1 U39 ( .A(n3), .Y(n4) );
  AND2X2 U42 ( .A(n2), .B(n4), .Y(n5) );
  AND2X2 U45 ( .A(\addr<1> ), .B(\busy<3> ), .Y(n6) );
  AND2X2 U48 ( .A(\addr<1> ), .B(\busy<1> ), .Y(n7) );
  INVX1 U51 ( .A(n7), .Y(n8) );
  INVX1 U54 ( .A(n6), .Y(n12) );
  INVX1 U57 ( .A(n14), .Y(n15) );
  AND2X1 U60 ( .A(n105), .B(n106), .Y(n17) );
  INVX1 U63 ( .A(n17), .Y(n18) );
  AND2X1 U66 ( .A(n20), .B(n106), .Y(n19) );
  INVX1 U69 ( .A(n19), .Y(n21) );
  AND2X1 U72 ( .A(n11), .B(n105), .Y(n55) );
  INVX1 U79 ( .A(n55), .Y(n56) );
  INVX1 U80 ( .A(\addr<1> ), .Y(n105) );
  AND2X2 U81 ( .A(\addr<2> ), .B(\addr<1> ), .Y(n57) );
  INVX1 U82 ( .A(n57), .Y(n58) );
  AND2X2 U83 ( .A(n52), .B(n53), .Y(n59) );
  INVX1 U84 ( .A(n59), .Y(\data_out<0> ) );
  AND2X2 U85 ( .A(n50), .B(n51), .Y(n61) );
  INVX1 U86 ( .A(n61), .Y(\data_out<10> ) );
  AND2X2 U87 ( .A(n48), .B(n49), .Y(n63) );
  INVX1 U88 ( .A(n63), .Y(\data_out<11> ) );
  AND2X2 U89 ( .A(n46), .B(n47), .Y(n65) );
  INVX1 U90 ( .A(n65), .Y(\data_out<12> ) );
  AND2X2 U91 ( .A(n44), .B(n45), .Y(n67) );
  INVX1 U92 ( .A(n67), .Y(\data_out<13> ) );
  AND2X2 U93 ( .A(n42), .B(n43), .Y(n69) );
  INVX1 U94 ( .A(n69), .Y(\data_out<14> ) );
  AND2X2 U95 ( .A(n40), .B(n41), .Y(n71) );
  INVX1 U96 ( .A(n71), .Y(\data_out<15> ) );
  AND2X2 U97 ( .A(n38), .B(n39), .Y(n73) );
  INVX1 U98 ( .A(n73), .Y(\data_out<1> ) );
  AND2X2 U99 ( .A(n36), .B(n37), .Y(n75) );
  INVX1 U100 ( .A(n75), .Y(\data_out<2> ) );
  AND2X2 U101 ( .A(n34), .B(n35), .Y(n77) );
  INVX1 U102 ( .A(n77), .Y(\data_out<3> ) );
  AND2X2 U103 ( .A(n32), .B(n33), .Y(n79) );
  INVX1 U104 ( .A(n79), .Y(\data_out<4> ) );
  AND2X2 U105 ( .A(n30), .B(n31), .Y(n81) );
  INVX1 U106 ( .A(n81), .Y(\data_out<5> ) );
  AND2X2 U107 ( .A(n28), .B(n29), .Y(n83) );
  INVX1 U108 ( .A(n83), .Y(\data_out<6> ) );
  AND2X2 U109 ( .A(n26), .B(n27), .Y(n85) );
  INVX1 U110 ( .A(n85), .Y(\data_out<7> ) );
  AND2X2 U111 ( .A(n24), .B(n25), .Y(n87) );
  INVX1 U112 ( .A(n87), .Y(\data_out<8> ) );
  AND2X2 U113 ( .A(n22), .B(n23), .Y(n89) );
  INVX1 U114 ( .A(n89), .Y(\data_out<9> ) );
  INVX1 U115 ( .A(n91), .Y(n92) );
  INVX1 U116 ( .A(\addr<4> ), .Y(n98) );
  INVX1 U117 ( .A(\addr<3> ), .Y(n96) );
  INVX8 U118 ( .A(n94), .Y(n93) );
endmodule


module dff_264 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_263 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_245 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_246 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_247 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_248 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_249 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_250 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_251 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_252 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_253 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_254 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_255 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_256 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_257 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_258 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_259 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_260 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_262 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_229 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_230 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_231 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_232 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_233 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_234 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_235 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2, n3;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n2), .B(n3), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
endmodule


module dff_236 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_237 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_238 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2, n3;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n2), .B(n3), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n3) );
  INVX1 U5 ( .A(d), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n2) );
endmodule


module dff_239 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_240 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_241 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_242 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_243 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_244 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_261 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_224 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_225 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_226 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X2 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_227 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(d), .B(n1), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n1) );
endmodule


module dff_228 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1, n2;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  AND2X1 U3 ( .A(n1), .B(n2), .Y(N3) );
  INVX1 U4 ( .A(rst), .Y(n2) );
  BUFX2 U5 ( .A(d), .Y(n1) );
endmodule


module dff_221 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_222 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_223 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_216 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_217 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_218 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_219 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module dff_220 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   N3, n1;

  DFFPOSX1 state_reg ( .D(N3), .CLK(clk), .Q(q) );
  NOR2X1 U4 ( .A(rst), .B(n1), .Y(N3) );
  INVX1 U3 ( .A(d), .Y(n1) );
endmodule


module mem_system ( .DataOut({\DataOut<15> , \DataOut<14> , \DataOut<13> , 
        \DataOut<12> , \DataOut<11> , \DataOut<10> , \DataOut<9> , 
        \DataOut<8> , \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , 
        \DataOut<3> , \DataOut<2> , \DataOut<1> , \DataOut<0> }), Done, Stall, 
        CacheHit, err, .Addr({\Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , 
        \Addr<11> , \Addr<10> , \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , 
        \Addr<5> , \Addr<4> , \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> }), 
    .DataIn({\DataIn<15> , \DataIn<14> , \DataIn<13> , \DataIn<12> , 
        \DataIn<11> , \DataIn<10> , \DataIn<9> , \DataIn<8> , \DataIn<7> , 
        \DataIn<6> , \DataIn<5> , \DataIn<4> , \DataIn<3> , \DataIn<2> , 
        \DataIn<1> , \DataIn<0> }), Rd, Wr, createdump, clk, rst );
  input \Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , \Addr<11> , \Addr<10> ,
         \Addr<9> , \Addr<8> , \Addr<7> , \Addr<6> , \Addr<5> , \Addr<4> ,
         \Addr<3> , \Addr<2> , \Addr<1> , \Addr<0> , \DataIn<15> ,
         \DataIn<14> , \DataIn<13> , \DataIn<12> , \DataIn<11> , \DataIn<10> ,
         \DataIn<9> , \DataIn<8> , \DataIn<7> , \DataIn<6> , \DataIn<5> ,
         \DataIn<4> , \DataIn<3> , \DataIn<2> , \DataIn<1> , \DataIn<0> , Rd,
         Wr, createdump, clk, rst;
  output \DataOut<15> , \DataOut<14> , \DataOut<13> , \DataOut<12> ,
         \DataOut<11> , \DataOut<10> , \DataOut<9> , \DataOut<8> ,
         \DataOut<7> , \DataOut<6> , \DataOut<5> , \DataOut<4> , \DataOut<3> ,
         \DataOut<2> , \DataOut<1> , \DataOut<0> , Done, Stall, CacheHit, err;
  wire   \tagOut<4> , \tagOut<3> , \tagOut<2> , \tagOut<1> , \tagOut<0> ,
         \cacheDataOut<15> , \cacheDataOut<14> , \cacheDataOut<13> ,
         \cacheDataOut<12> , \cacheDataOut<11> , \cacheDataOut<10> ,
         \cacheDataOut<9> , \cacheDataOut<8> , \cacheDataOut<7> ,
         \cacheDataOut<6> , \cacheDataOut<5> , \cacheDataOut<4> ,
         \cacheDataOut<3> , \cacheDataOut<2> , \cacheDataOut<1> ,
         \cacheDataOut<0> , cacheHit, dirty, valid, \cacheOff<2> ,
         \cacheOff<0> , \cacheDataIn<15> , \cacheDataIn<14> ,
         \cacheDataIn<13> , \cacheDataIn<12> , \cacheDataIn<11> ,
         \cacheDataIn<10> , \cacheDataIn<9> , \cacheDataIn<8> ,
         \cacheDataIn<7> , \cacheDataIn<6> , \cacheDataIn<5> ,
         \cacheDataIn<4> , \cacheDataIn<3> , \cacheDataIn<2> ,
         \cacheDataIn<1> , \cacheDataIn<0> , memAddr_0, \memDataIn<15> ,
         \memDataIn<14> , \memDataIn<13> , \memDataIn<12> , \memDataIn<11> ,
         \memDataIn<10> , \memDataIn<9> , \memDataIn<8> , \memDataIn<7> ,
         \memDataIn<6> , \memDataIn<5> , \memDataIn<4> , \memDataIn<3> ,
         \memDataIn<2> , \memDataIn<1> , \memDataIn<0> , \memDataOut<15> ,
         \memDataOut<14> , \memDataOut<13> , \memDataOut<12> ,
         \memDataOut<11> , \memDataOut<10> , \memDataOut<9> , \memDataOut<8> ,
         \memDataOut<7> , \memDataOut<6> , \memDataOut<5> , \memDataOut<4> ,
         \memDataOut<3> , \memDataOut<2> , \memDataOut<1> , \memDataOut<0> ,
         memStall, doneWait_in, \memDataOut_flop<15> , \memDataOut_flop<14> ,
         \memDataOut_flop<13> , \memDataOut_flop<12> , \memDataOut_flop<11> ,
         \memDataOut_flop<10> , \memDataOut_flop<9> , \memDataOut_flop<8> ,
         \memDataOut_flop<7> , \memDataOut_flop<6> , \memDataOut_flop<5> ,
         \memDataOut_flop<4> , \memDataOut_flop<3> , \memDataOut_flop<2> ,
         \memDataOut_flop<1> , \memDataOut_flop<0> , waitMem_flop,
         \cacheDataOut_flop<15> , \cacheDataOut_flop<14> ,
         \cacheDataOut_flop<13> , \cacheDataOut_flop<12> ,
         \cacheDataOut_flop<11> , \cacheDataOut_flop<10> ,
         \cacheDataOut_flop<9> , \cacheDataOut_flop<8> ,
         \cacheDataOut_flop<7> , \cacheDataOut_flop<6> ,
         \cacheDataOut_flop<5> , \cacheDataOut_flop<4> ,
         \cacheDataOut_flop<3> , \cacheDataOut_flop<2> ,
         \cacheDataOut_flop<1> , \cacheDataOut_flop<0> , waitCacheHit_in,
         \nxtState<4> , \nxtState<2> , \nxtState<1> , \nxtState<0> ,
         \state<4> , \state<3> , \state<2> , \state<1> , \state<0> ,
         \wait4Cycles_flop<0> , \wait4Cycles_in<1> , \wait4Cycles_in<0> ,
         \nextEvictState_in<0> , \nxtEvict<4> , \nxtEvict<3> , \nxtEvict<2> ,
         \nxtEvict<1> , \nxtEvict<0> , n5, n9, n11, n192, n230, n235, n242,
         n245, n246, n247, n248, n250, n269, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797;

  XOR2X1 U7 ( .A(n355), .B(n329), .Y(n5) );
  MUX2X1 U27 ( .B(n765), .A(n797), .S(n9), .Y(\cacheDataIn<0> ) );
  MUX2X1 U30 ( .B(n766), .A(n796), .S(n11), .Y(\cacheDataIn<1> ) );
  MUX2X1 U32 ( .B(n767), .A(n795), .S(n740), .Y(\cacheDataIn<2> ) );
  MUX2X1 U33 ( .B(n768), .A(n794), .S(n740), .Y(\cacheDataIn<3> ) );
  MUX2X1 U34 ( .B(n769), .A(n793), .S(n740), .Y(\cacheDataIn<4> ) );
  MUX2X1 U35 ( .B(n770), .A(n792), .S(n740), .Y(\cacheDataIn<5> ) );
  MUX2X1 U36 ( .B(n771), .A(n791), .S(n740), .Y(\cacheDataIn<6> ) );
  MUX2X1 U37 ( .B(n772), .A(n790), .S(n740), .Y(\cacheDataIn<7> ) );
  MUX2X1 U38 ( .B(n773), .A(n789), .S(n740), .Y(\cacheDataIn<8> ) );
  MUX2X1 U39 ( .B(n774), .A(n788), .S(n740), .Y(\cacheDataIn<9> ) );
  MUX2X1 U40 ( .B(n775), .A(n787), .S(n740), .Y(\cacheDataIn<10> ) );
  MUX2X1 U41 ( .B(n776), .A(n786), .S(n740), .Y(\cacheDataIn<11> ) );
  MUX2X1 U42 ( .B(n777), .A(n785), .S(n740), .Y(\cacheDataIn<12> ) );
  MUX2X1 U43 ( .B(n778), .A(n784), .S(n740), .Y(\cacheDataIn<13> ) );
  MUX2X1 U44 ( .B(n779), .A(n783), .S(n740), .Y(\cacheDataIn<14> ) );
  MUX2X1 U45 ( .B(n780), .A(n782), .S(n740), .Y(\cacheDataIn<15> ) );
  AND2X2 U109 ( .A(valid), .B(cacheHit), .Y(waitCacheHit_in) );
  AND2X2 U123 ( .A(\Addr<0> ), .B(n591), .Y(\cacheOff<0> ) );
  NAND3X1 U230 ( .A(n741), .B(n781), .C(\Addr<1> ), .Y(n192) );
  AOI21X1 U262 ( .A(\Addr<2> ), .B(n596), .C(n742), .Y(n230) );
  AOI22X1 U269 ( .A(\Addr<15> ), .B(n478), .C(\tagOut<4> ), .D(n480), .Y(n242)
         );
  AOI22X1 U270 ( .A(\Addr<14> ), .B(n478), .C(\tagOut<3> ), .D(n480), .Y(n245)
         );
  AOI22X1 U271 ( .A(\Addr<13> ), .B(n478), .C(\tagOut<2> ), .D(n480), .Y(n246)
         );
  AOI22X1 U272 ( .A(\Addr<12> ), .B(n478), .C(\tagOut<1> ), .D(n480), .Y(n247)
         );
  AOI22X1 U273 ( .A(\Addr<11> ), .B(n478), .C(\tagOut<0> ), .D(n480), .Y(n248)
         );
  AOI22X1 U342 ( .A(waitMem_flop), .B(\cacheDataOut_flop<9> ), .C(
        \memDataOut_flop<9> ), .D(n759), .Y(n283) );
  AOI22X1 U343 ( .A(\cacheDataOut_flop<8> ), .B(waitMem_flop), .C(
        \memDataOut_flop<8> ), .D(n759), .Y(n284) );
  AOI22X1 U344 ( .A(\cacheDataOut_flop<7> ), .B(waitMem_flop), .C(
        \memDataOut_flop<7> ), .D(n759), .Y(n285) );
  AOI22X1 U345 ( .A(\cacheDataOut_flop<6> ), .B(waitMem_flop), .C(
        \memDataOut_flop<6> ), .D(n759), .Y(n286) );
  AOI22X1 U346 ( .A(\cacheDataOut_flop<5> ), .B(waitMem_flop), .C(
        \memDataOut_flop<5> ), .D(n759), .Y(n287) );
  AOI22X1 U347 ( .A(\cacheDataOut_flop<4> ), .B(waitMem_flop), .C(
        \memDataOut_flop<4> ), .D(n759), .Y(n288) );
  AOI22X1 U348 ( .A(\cacheDataOut_flop<3> ), .B(waitMem_flop), .C(
        \memDataOut_flop<3> ), .D(n759), .Y(n289) );
  AOI22X1 U349 ( .A(\cacheDataOut_flop<2> ), .B(waitMem_flop), .C(
        \memDataOut_flop<2> ), .D(n759), .Y(n290) );
  AOI22X1 U350 ( .A(\cacheDataOut_flop<1> ), .B(waitMem_flop), .C(
        \memDataOut_flop<1> ), .D(n759), .Y(n291) );
  AOI22X1 U351 ( .A(\cacheDataOut_flop<15> ), .B(waitMem_flop), .C(
        \memDataOut_flop<15> ), .D(n759), .Y(n292) );
  AOI22X1 U352 ( .A(\cacheDataOut_flop<14> ), .B(waitMem_flop), .C(
        \memDataOut_flop<14> ), .D(n759), .Y(n293) );
  AOI22X1 U353 ( .A(\cacheDataOut_flop<13> ), .B(waitMem_flop), .C(
        \memDataOut_flop<13> ), .D(n759), .Y(n294) );
  AOI22X1 U354 ( .A(\cacheDataOut_flop<12> ), .B(waitMem_flop), .C(
        \memDataOut_flop<12> ), .D(n759), .Y(n295) );
  AOI22X1 U355 ( .A(\cacheDataOut_flop<11> ), .B(waitMem_flop), .C(
        \memDataOut_flop<11> ), .D(n759), .Y(n296) );
  AOI22X1 U356 ( .A(\cacheDataOut_flop<10> ), .B(waitMem_flop), .C(
        \memDataOut_flop<10> ), .D(n759), .Y(n297) );
  AOI22X1 U357 ( .A(\cacheDataOut_flop<0> ), .B(waitMem_flop), .C(
        \memDataOut_flop<0> ), .D(n759), .Y(n298) );
  cache_cache_id0 c0 ( .enable(n386), .clk(clk), .rst(n633), .createdump(
        createdump), .tag_in({\Addr<15> , \Addr<14> , \Addr<13> , \Addr<12> , 
        \Addr<11> }), .index({n629, n628, n627, n641, n639, n637, n331, 
        \Addr<3> }), .offset({n611, n614, \cacheOff<0> }), .data_in({
        \cacheDataIn<15> , \cacheDataIn<14> , \cacheDataIn<13> , 
        \cacheDataIn<12> , \cacheDataIn<11> , \cacheDataIn<10> , 
        \cacheDataIn<9> , \cacheDataIn<8> , \cacheDataIn<7> , \cacheDataIn<6> , 
        \cacheDataIn<5> , \cacheDataIn<4> , \cacheDataIn<3> , \cacheDataIn<2> , 
        \cacheDataIn<1> , \cacheDataIn<0> }), .comp(n357), .write(n362), 
        .valid_in(n597), .tag_out({\tagOut<4> , \tagOut<3> , \tagOut<2> , 
        \tagOut<1> , \tagOut<0> }), .data_out({\cacheDataOut<15> , 
        \cacheDataOut<14> , \cacheDataOut<13> , \cacheDataOut<12> , 
        \cacheDataOut<11> , \cacheDataOut<10> , \cacheDataOut<9> , 
        \cacheDataOut<8> , \cacheDataOut<7> , \cacheDataOut<6> , 
        \cacheDataOut<5> , \cacheDataOut<4> , \cacheDataOut<3> , 
        \cacheDataOut<2> , \cacheDataOut<1> , \cacheDataOut<0> }), .hit(
        cacheHit), .dirty(dirty), .valid(valid), .err() );
  four_bank_mem fmem ( .clk(clk), .rst(n631), .createdump(createdump), .addr({
        n764, n763, n762, n761, n760, n629, n628, n627, n641, n639, n637, n635, 
        n316, n369, n372, memAddr_0}), .data_in({\memDataIn<15> , 
        \memDataIn<14> , \memDataIn<13> , \memDataIn<12> , \memDataIn<11> , 
        \memDataIn<10> , \memDataIn<9> , \memDataIn<8> , \memDataIn<7> , 
        \memDataIn<6> , \memDataIn<5> , \memDataIn<4> , \memDataIn<3> , 
        \memDataIn<2> , \memDataIn<1> , \memDataIn<0> }), .wr(n616), .rd(n618), 
        .data_out({\memDataOut<15> , \memDataOut<14> , \memDataOut<13> , 
        \memDataOut<12> , \memDataOut<11> , \memDataOut<10> , \memDataOut<9> , 
        \memDataOut<8> , \memDataOut<7> , \memDataOut<6> , \memDataOut<5> , 
        \memDataOut<4> , \memDataOut<3> , \memDataOut<2> , \memDataOut<1> , 
        \memDataOut<0> }), .stall(memStall), .busy(), .err() );
  dff_264 waitStall ( .q(Stall), .d(n358), .clk(clk), .rst(n632) );
  dff_263 waitDone ( .q(Done), .d(doneWait_in), .clk(clk), .rst(n633) );
  dff_245 \memDataOutWait[0]  ( .q(\memDataOut_flop<0> ), .d(\memDataOut<0> ), 
        .clk(clk), .rst(n632) );
  dff_246 \memDataOutWait[1]  ( .q(\memDataOut_flop<1> ), .d(\memDataOut<1> ), 
        .clk(clk), .rst(n633) );
  dff_247 \memDataOutWait[2]  ( .q(\memDataOut_flop<2> ), .d(\memDataOut<2> ), 
        .clk(clk), .rst(n631) );
  dff_248 \memDataOutWait[3]  ( .q(\memDataOut_flop<3> ), .d(\memDataOut<3> ), 
        .clk(clk), .rst(n631) );
  dff_249 \memDataOutWait[4]  ( .q(\memDataOut_flop<4> ), .d(\memDataOut<4> ), 
        .clk(clk), .rst(n632) );
  dff_250 \memDataOutWait[5]  ( .q(\memDataOut_flop<5> ), .d(\memDataOut<5> ), 
        .clk(clk), .rst(n633) );
  dff_251 \memDataOutWait[6]  ( .q(\memDataOut_flop<6> ), .d(\memDataOut<6> ), 
        .clk(clk), .rst(n631) );
  dff_252 \memDataOutWait[7]  ( .q(\memDataOut_flop<7> ), .d(\memDataOut<7> ), 
        .clk(clk), .rst(n632) );
  dff_253 \memDataOutWait[8]  ( .q(\memDataOut_flop<8> ), .d(\memDataOut<8> ), 
        .clk(clk), .rst(n631) );
  dff_254 \memDataOutWait[9]  ( .q(\memDataOut_flop<9> ), .d(\memDataOut<9> ), 
        .clk(clk), .rst(n632) );
  dff_255 \memDataOutWait[10]  ( .q(\memDataOut_flop<10> ), .d(
        \memDataOut<10> ), .clk(clk), .rst(n633) );
  dff_256 \memDataOutWait[11]  ( .q(\memDataOut_flop<11> ), .d(
        \memDataOut<11> ), .clk(clk), .rst(n631) );
  dff_257 \memDataOutWait[12]  ( .q(\memDataOut_flop<12> ), .d(
        \memDataOut<12> ), .clk(clk), .rst(n632) );
  dff_258 \memDataOutWait[13]  ( .q(\memDataOut_flop<13> ), .d(
        \memDataOut<13> ), .clk(clk), .rst(n633) );
  dff_259 \memDataOutWait[14]  ( .q(\memDataOut_flop<14> ), .d(
        \memDataOut<14> ), .clk(clk), .rst(n631) );
  dff_260 \memDataOutWait[15]  ( .q(\memDataOut_flop<15> ), .d(
        \memDataOut<15> ), .clk(clk), .rst(n632) );
  dff_262 waitMem ( .q(waitMem_flop), .d(n419), .clk(clk), .rst(n633) );
  dff_229 \cacheDataOutWait[0]  ( .q(\cacheDataOut_flop<0> ), .d(n626), .clk(
        clk), .rst(n631) );
  dff_230 \cacheDataOutWait[1]  ( .q(\cacheDataOut_flop<1> ), .d(n625), .clk(
        clk), .rst(n632) );
  dff_231 \cacheDataOutWait[2]  ( .q(\cacheDataOut_flop<2> ), .d(n624), .clk(
        clk), .rst(n633) );
  dff_232 \cacheDataOutWait[3]  ( .q(\cacheDataOut_flop<3> ), .d(n623), .clk(
        clk), .rst(n632) );
  dff_233 \cacheDataOutWait[4]  ( .q(\cacheDataOut_flop<4> ), .d(
        \cacheDataOut<4> ), .clk(clk), .rst(n633) );
  dff_234 \cacheDataOutWait[5]  ( .q(\cacheDataOut_flop<5> ), .d(
        \cacheDataOut<5> ), .clk(clk), .rst(n631) );
  dff_235 \cacheDataOutWait[6]  ( .q(\cacheDataOut_flop<6> ), .d(
        \cacheDataOut<6> ), .clk(clk), .rst(n632) );
  dff_236 \cacheDataOutWait[7]  ( .q(\cacheDataOut_flop<7> ), .d(
        \cacheDataOut<7> ), .clk(clk), .rst(n631) );
  dff_237 \cacheDataOutWait[8]  ( .q(\cacheDataOut_flop<8> ), .d(n310), .clk(
        clk), .rst(n631) );
  dff_238 \cacheDataOutWait[9]  ( .q(\cacheDataOut_flop<9> ), .d(
        \cacheDataOut<9> ), .clk(clk), .rst(n632) );
  dff_239 \cacheDataOutWait[10]  ( .q(\cacheDataOut_flop<10> ), .d(
        \cacheDataOut<10> ), .clk(clk), .rst(n633) );
  dff_240 \cacheDataOutWait[11]  ( .q(\cacheDataOut_flop<11> ), .d(
        \cacheDataOut<11> ), .clk(clk), .rst(n631) );
  dff_241 \cacheDataOutWait[12]  ( .q(\cacheDataOut_flop<12> ), .d(n335), 
        .clk(clk), .rst(n632) );
  dff_242 \cacheDataOutWait[13]  ( .q(\cacheDataOut_flop<13> ), .d(
        \cacheDataOut<13> ), .clk(clk), .rst(n633) );
  dff_243 \cacheDataOutWait[14]  ( .q(\cacheDataOut_flop<14> ), .d(n312), 
        .clk(clk), .rst(n631) );
  dff_244 \cacheDataOutWait[15]  ( .q(\cacheDataOut_flop<15> ), .d(n619), 
        .clk(clk), .rst(n632) );
  dff_261 waitCacheHit ( .q(CacheHit), .d(waitCacheHit_in), .clk(clk), .rst(
        n633) );
  dff_224 \stateReg[0]  ( .q(\state<0> ), .d(n495), .clk(clk), .rst(n633) );
  dff_225 \stateReg[1]  ( .q(\state<1> ), .d(\nxtState<1> ), .clk(clk), .rst(
        n631) );
  dff_226 \stateReg[2]  ( .q(\state<2> ), .d(\nxtState<2> ), .clk(clk), .rst(
        n632) );
  dff_227 \stateReg[3]  ( .q(\state<3> ), .d(n493), .clk(clk), .rst(n633) );
  dff_228 \stateReg[4]  ( .q(\state<4> ), .d(\nxtState<4> ), .clk(clk), .rst(
        n631) );
  dff_221 \wait4CycleFlop[0]  ( .q(\wait4Cycles_flop<0> ), .d(
        \wait4Cycles_in<0> ), .clk(clk), .rst(n633) );
  dff_222 \wait4CycleFlop[1]  ( .q(\wait4Cycles_in<0> ), .d(
        \wait4Cycles_in<1> ), .clk(clk), .rst(n632) );
  dff_223 \wait4CycleFlop[2]  ( .q(\wait4Cycles_in<1> ), .d(n453), .clk(clk), 
        .rst(n631) );
  dff_216 \evictWait[0]  ( .q(\nxtEvict<0> ), .d(\nextEvictState_in<0> ), 
        .clk(clk), .rst(n633) );
  dff_217 \evictWait[1]  ( .q(\nxtEvict<1> ), .d(n468), .clk(clk), .rst(n632)
         );
  dff_218 \evictWait[2]  ( .q(\nxtEvict<2> ), .d(n567), .clk(clk), .rst(n631)
         );
  dff_219 \evictWait[3]  ( .q(\nxtEvict<3> ), .d(n589), .clk(clk), .rst(n633)
         );
  dff_220 \evictWait[4]  ( .q(\nxtEvict<4> ), .d(n475), .clk(clk), .rst(n632)
         );
  INVX1 U358 ( .A(\state<1> ), .Y(n299) );
  INVX1 U359 ( .A(n299), .Y(n300) );
  AND2X1 U360 ( .A(n568), .B(n416), .Y(n615) );
  AND2X1 U361 ( .A(n388), .B(n497), .Y(n617) );
  INVX1 U362 ( .A(\DataIn<5> ), .Y(n792) );
  INVX1 U363 ( .A(\DataIn<6> ), .Y(n791) );
  INVX1 U364 ( .A(\DataIn<15> ), .Y(n782) );
  AND2X1 U365 ( .A(n412), .B(n431), .Y(n507) );
  INVX1 U366 ( .A(n345), .Y(n433) );
  AND2X1 U367 ( .A(n412), .B(n571), .Y(n578) );
  OR2X1 U368 ( .A(n446), .B(n329), .Y(n424) );
  INVX1 U369 ( .A(n738), .Y(n740) );
  INVX1 U370 ( .A(Rd), .Y(n679) );
  INVX1 U371 ( .A(n663), .Y(n665) );
  INVX1 U372 ( .A(\Addr<2> ), .Y(n781) );
  OR2X1 U373 ( .A(\wait4Cycles_in<1> ), .B(\wait4Cycles_in<0> ), .Y(n663) );
  AND2X1 U374 ( .A(n412), .B(n603), .Y(n513) );
  INVX1 U375 ( .A(n662), .Y(n681) );
  OR2X1 U376 ( .A(n576), .B(n317), .Y(n662) );
  INVX1 U377 ( .A(\DataIn<0> ), .Y(n797) );
  INVX1 U378 ( .A(\DataIn<8> ), .Y(n789) );
  INVX1 U379 ( .A(\DataIn<10> ), .Y(n787) );
  INVX1 U380 ( .A(\DataIn<11> ), .Y(n786) );
  INVX1 U381 ( .A(\DataIn<13> ), .Y(n784) );
  OR2X1 U382 ( .A(n465), .B(n510), .Y(n556) );
  INVX1 U383 ( .A(\nxtEvict<3> ), .Y(n654) );
  INVX1 U384 ( .A(n634), .Y(n631) );
  BUFX2 U385 ( .A(\Addr<8> ), .Y(n627) );
  BUFX2 U386 ( .A(\Addr<9> ), .Y(n628) );
  BUFX2 U387 ( .A(\Addr<10> ), .Y(n629) );
  INVX1 U388 ( .A(n448), .Y(n302) );
  INVX1 U389 ( .A(n448), .Y(n303) );
  INVX1 U390 ( .A(n448), .Y(n301) );
  OR2X1 U391 ( .A(n508), .B(n512), .Y(n558) );
  AND2X1 U392 ( .A(n603), .B(n440), .Y(n511) );
  AND2X1 U393 ( .A(n328), .B(n412), .Y(n467) );
  INVX1 U394 ( .A(n704), .Y(n352) );
  AND2X1 U395 ( .A(n341), .B(n420), .Y(n606) );
  INVX1 U396 ( .A(Wr), .Y(n354) );
  INVX1 U397 ( .A(n603), .Y(n650) );
  AND2X1 U398 ( .A(n329), .B(n733), .Y(n441) );
  INVX1 U399 ( .A(\memDataOut<0> ), .Y(n765) );
  INVX1 U400 ( .A(\memDataOut<1> ), .Y(n766) );
  INVX1 U401 ( .A(\memDataOut<2> ), .Y(n767) );
  INVX1 U402 ( .A(\memDataOut<3> ), .Y(n768) );
  INVX1 U403 ( .A(\memDataOut<4> ), .Y(n769) );
  INVX1 U404 ( .A(\memDataOut<5> ), .Y(n770) );
  INVX1 U405 ( .A(\memDataOut<6> ), .Y(n771) );
  INVX1 U406 ( .A(\memDataOut<7> ), .Y(n772) );
  INVX1 U407 ( .A(\memDataOut<8> ), .Y(n773) );
  INVX1 U408 ( .A(\memDataOut<9> ), .Y(n774) );
  INVX1 U409 ( .A(\memDataOut<10> ), .Y(n775) );
  INVX1 U410 ( .A(\memDataOut<11> ), .Y(n776) );
  INVX1 U411 ( .A(\memDataOut<12> ), .Y(n777) );
  INVX1 U412 ( .A(\memDataOut<13> ), .Y(n778) );
  INVX1 U413 ( .A(\memDataOut<14> ), .Y(n779) );
  INVX1 U414 ( .A(\memDataOut<15> ), .Y(n780) );
  OR2X1 U415 ( .A(n705), .B(n679), .Y(n516) );
  AND2X1 U416 ( .A(n448), .B(n496), .Y(n560) );
  AND2X1 U417 ( .A(\Addr<2> ), .B(n348), .Y(n661) );
  AND2X1 U418 ( .A(n533), .B(n381), .Y(n502) );
  INVX1 U419 ( .A(\Addr<0> ), .Y(n657) );
  INVX1 U420 ( .A(n371), .Y(n372) );
  OR2X1 U421 ( .A(n491), .B(n532), .Y(n474) );
  INVX1 U422 ( .A(\Addr<6> ), .Y(n640) );
  INVX1 U423 ( .A(\Addr<7> ), .Y(n642) );
  INVX1 U424 ( .A(\DataIn<1> ), .Y(n796) );
  INVX1 U425 ( .A(\DataIn<2> ), .Y(n795) );
  INVX1 U426 ( .A(\DataIn<3> ), .Y(n794) );
  INVX1 U427 ( .A(\DataIn<4> ), .Y(n793) );
  INVX1 U428 ( .A(\DataIn<7> ), .Y(n790) );
  INVX1 U429 ( .A(\DataIn<9> ), .Y(n788) );
  INVX1 U430 ( .A(\DataIn<12> ), .Y(n785) );
  INVX1 U431 ( .A(\DataIn<14> ), .Y(n783) );
  AND2X1 U432 ( .A(n586), .B(n601), .Y(n588) );
  AND2X1 U433 ( .A(\Addr<0> ), .B(n596), .Y(memAddr_0) );
  AND2X1 U434 ( .A(n408), .B(n598), .Y(n691) );
  MUX2X1 U435 ( .B(n315), .A(n782), .S(n301), .Y(\memDataIn<15> ) );
  MUX2X1 U436 ( .B(n727), .A(n792), .S(n302), .Y(\memDataIn<5> ) );
  MUX2X1 U437 ( .B(n724), .A(n789), .S(n447), .Y(\memDataIn<8> ) );
  INVX2 U438 ( .A(n447), .Y(n448) );
  MUX2X1 U439 ( .B(n726), .A(n791), .S(n303), .Y(\memDataIn<6> ) );
  MUX2X1 U440 ( .B(n336), .A(n797), .S(n447), .Y(\memDataIn<0> ) );
  INVX1 U441 ( .A(n355), .Y(n304) );
  INVX1 U442 ( .A(\state<1> ), .Y(n693) );
  AND2X1 U443 ( .A(n326), .B(n410), .Y(n484) );
  AND2X1 U444 ( .A(n344), .B(n341), .Y(n488) );
  AND2X1 U445 ( .A(n426), .B(n442), .Y(n486) );
  OR2X1 U446 ( .A(n504), .B(n514), .Y(n491) );
  OR2X1 U447 ( .A(\wait4Cycles_in<1> ), .B(n363), .Y(n305) );
  OR2X1 U448 ( .A(\wait4Cycles_in<0> ), .B(\wait4Cycles_flop<0> ), .Y(n306) );
  OR2X1 U449 ( .A(n314), .B(n427), .Y(n307) );
  OR2X1 U450 ( .A(n344), .B(n535), .Y(n471) );
  INVX1 U451 ( .A(\Addr<1> ), .Y(n348) );
  INVX1 U452 ( .A(n683), .Y(n741) );
  AND2X1 U453 ( .A(n327), .B(n317), .Y(n490) );
  AND2X1 U454 ( .A(n329), .B(n340), .Y(n391) );
  AND2X1 U455 ( .A(n547), .B(n593), .Y(n377) );
  OR2X2 U456 ( .A(n432), .B(n433), .Y(n308) );
  INVX2 U457 ( .A(\state<0> ), .Y(n712) );
  INVX1 U458 ( .A(rst), .Y(n634) );
  INVX1 U459 ( .A(\cacheDataOut<8> ), .Y(n309) );
  INVX1 U460 ( .A(n309), .Y(n310) );
  INVX1 U461 ( .A(\cacheDataOut<14> ), .Y(n311) );
  INVX1 U462 ( .A(n311), .Y(n312) );
  INVX1 U463 ( .A(\cacheDataOut<1> ), .Y(n313) );
  INVX1 U464 ( .A(n693), .Y(n314) );
  INVX1 U465 ( .A(\cacheDataOut<15> ), .Y(n315) );
  BUFX2 U466 ( .A(\Addr<3> ), .Y(n316) );
  OR2X1 U467 ( .A(n435), .B(n307), .Y(n317) );
  INVX1 U468 ( .A(n317), .Y(n318) );
  AND2X2 U469 ( .A(n598), .B(n390), .Y(n319) );
  AND2X2 U470 ( .A(\state<2> ), .B(n695), .Y(n320) );
  AND2X2 U471 ( .A(n709), .B(\state<3> ), .Y(n321) );
  AND2X2 U472 ( .A(n712), .B(n742), .Y(n322) );
  INVX1 U473 ( .A(n322), .Y(n323) );
  INVX1 U474 ( .A(n321), .Y(n324) );
  AND2X2 U475 ( .A(n712), .B(n441), .Y(n325) );
  INVX1 U476 ( .A(n325), .Y(n326) );
  INVX1 U477 ( .A(n325), .Y(n327) );
  INVX1 U478 ( .A(n653), .Y(n328) );
  BUFX2 U479 ( .A(\state<4> ), .Y(n329) );
  BUFX2 U480 ( .A(dirty), .Y(n330) );
  INVX1 U481 ( .A(\state<4> ), .Y(n716) );
  INVX1 U482 ( .A(n636), .Y(n331) );
  AND2X2 U483 ( .A(\state<0> ), .B(n321), .Y(n332) );
  AND2X2 U484 ( .A(n351), .B(n319), .Y(n595) );
  OR2X2 U485 ( .A(\state<4> ), .B(\state<1> ), .Y(n644) );
  BUFX2 U486 ( .A(n599), .Y(n333) );
  INVX1 U487 ( .A(\cacheDataOut<12> ), .Y(n334) );
  INVX1 U488 ( .A(n334), .Y(n335) );
  INVX1 U489 ( .A(\cacheDataOut<0> ), .Y(n336) );
  INVX1 U490 ( .A(\Addr<4> ), .Y(n636) );
  INVX2 U491 ( .A(\Addr<5> ), .Y(n638) );
  INVX1 U492 ( .A(\cacheDataOut<3> ), .Y(n337) );
  INVX1 U493 ( .A(\cacheDataOut<2> ), .Y(n338) );
  BUFX2 U494 ( .A(n695), .Y(n339) );
  INVX1 U495 ( .A(n695), .Y(n340) );
  INVX1 U496 ( .A(n433), .Y(n341) );
  AND2X2 U497 ( .A(n428), .B(n713), .Y(n569) );
  INVX1 U498 ( .A(n320), .Y(n342) );
  INVX1 U499 ( .A(n342), .Y(n343) );
  INVX1 U500 ( .A(n342), .Y(n344) );
  INVX1 U501 ( .A(n644), .Y(n345) );
  INVX1 U502 ( .A(n644), .Y(n698) );
  NOR3X1 U503 ( .A(n365), .B(n352), .C(n401), .Y(n346) );
  OAI21X1 U504 ( .A(n348), .B(n595), .C(n578), .Y(n347) );
  INVX1 U505 ( .A(n347), .Y(n235) );
  OAI21X1 U506 ( .A(n400), .B(n399), .C(n586), .Y(n349) );
  INVX4 U507 ( .A(n586), .Y(n742) );
  AND2X2 U508 ( .A(n443), .B(n444), .Y(n602) );
  AND2X2 U509 ( .A(n713), .B(n443), .Y(n605) );
  AND2X2 U510 ( .A(n395), .B(n339), .Y(n350) );
  NOR3X1 U511 ( .A(n365), .B(n352), .C(n401), .Y(n351) );
  OR2X2 U512 ( .A(n398), .B(n471), .Y(n470) );
  OAI21X1 U513 ( .A(n354), .B(n705), .C(n377), .Y(n353) );
  INVX1 U514 ( .A(n353), .Y(n652) );
  BUFX2 U515 ( .A(\state<2> ), .Y(n355) );
  BUFX2 U516 ( .A(n376), .Y(n356) );
  INVX1 U517 ( .A(n599), .Y(n357) );
  AND2X2 U518 ( .A(n444), .B(n356), .Y(n594) );
  AND2X2 U519 ( .A(n344), .B(n443), .Y(n600) );
  AND2X2 U520 ( .A(n344), .B(n428), .Y(n483) );
  INVX1 U521 ( .A(\state<2> ), .Y(n709) );
  INVX1 U522 ( .A(n609), .Y(n696) );
  OR2X2 U523 ( .A(n360), .B(n359), .Y(n358) );
  OR2X2 U524 ( .A(n350), .B(n349), .Y(n359) );
  INVX1 U525 ( .A(n697), .Y(n360) );
  AND2X2 U526 ( .A(n702), .B(n701), .Y(n361) );
  INVX1 U527 ( .A(n361), .Y(n362) );
  OR2X1 U528 ( .A(n306), .B(n608), .Y(n363) );
  OR2X2 U529 ( .A(n434), .B(n308), .Y(n364) );
  INVX1 U530 ( .A(n364), .Y(n365) );
  OR2X2 U531 ( .A(n433), .B(n437), .Y(n366) );
  INVX1 U532 ( .A(n444), .Y(n436) );
  AND2X2 U533 ( .A(n553), .B(n368), .Y(n367) );
  AND2X2 U534 ( .A(n378), .B(n440), .Y(n368) );
  OR2X2 U535 ( .A(n587), .B(n474), .Y(n369) );
  AND2X2 U536 ( .A(n713), .B(n376), .Y(n370) );
  AND2X2 U537 ( .A(n235), .B(n482), .Y(n371) );
  AND2X2 U538 ( .A(n622), .B(n621), .Y(n373) );
  AND2X2 U539 ( .A(n321), .B(n698), .Y(n374) );
  AND2X2 U540 ( .A(n344), .B(n445), .Y(n375) );
  AND2X2 U541 ( .A(n698), .B(\state<0> ), .Y(n376) );
  AND2X2 U542 ( .A(n652), .B(n393), .Y(n378) );
  INVX1 U543 ( .A(n378), .Y(n379) );
  AND2X2 U544 ( .A(n665), .B(n664), .Y(n380) );
  INVX1 U545 ( .A(n380), .Y(n381) );
  AND2X2 U546 ( .A(n672), .B(n673), .Y(n382) );
  INVX1 U547 ( .A(n382), .Y(n383) );
  AND2X2 U548 ( .A(cacheHit), .B(dirty), .Y(n384) );
  AND2X2 U549 ( .A(n711), .B(n710), .Y(n385) );
  INVX1 U550 ( .A(n385), .Y(n386) );
  OR2X2 U551 ( .A(n742), .B(n486), .Y(n387) );
  INVX1 U552 ( .A(n387), .Y(n388) );
  OR2X1 U553 ( .A(n439), .B(n447), .Y(n389) );
  INVX1 U554 ( .A(n389), .Y(n390) );
  BUFX2 U555 ( .A(n708), .Y(n392) );
  BUFX2 U556 ( .A(n651), .Y(n393) );
  AND2X2 U557 ( .A(n429), .B(n694), .Y(n394) );
  INVX1 U558 ( .A(n394), .Y(n395) );
  AND2X2 U559 ( .A(\Addr<2> ), .B(n592), .Y(n396) );
  INVX1 U560 ( .A(n396), .Y(n397) );
  AND2X2 U561 ( .A(n716), .B(n300), .Y(n398) );
  AND2X2 U562 ( .A(n712), .B(n696), .Y(n399) );
  OR2X2 U563 ( .A(n304), .B(n329), .Y(n400) );
  OR2X2 U564 ( .A(n418), .B(n391), .Y(n401) );
  AND2X2 U565 ( .A(n660), .B(n659), .Y(n402) );
  INVX1 U566 ( .A(n402), .Y(n403) );
  AND2X2 U567 ( .A(n501), .B(n499), .Y(n404) );
  INVX1 U568 ( .A(n404), .Y(n405) );
  AND2X2 U569 ( .A(n398), .B(n332), .Y(n406) );
  INVX1 U570 ( .A(n406), .Y(n407) );
  INVX1 U571 ( .A(n406), .Y(n408) );
  AND2X2 U572 ( .A(n620), .B(n483), .Y(n409) );
  INVX1 U573 ( .A(n409), .Y(n410) );
  AND2X2 U574 ( .A(n712), .B(n569), .Y(n411) );
  INVX1 U575 ( .A(n411), .Y(n412) );
  AND2X2 U576 ( .A(n620), .B(n488), .Y(n413) );
  INVX1 U577 ( .A(n413), .Y(n414) );
  AND2X2 U578 ( .A(n716), .B(n715), .Y(n415) );
  INVX1 U579 ( .A(n415), .Y(n416) );
  AND2X2 U580 ( .A(n500), .B(n407), .Y(n417) );
  INVX1 U581 ( .A(n417), .Y(n418) );
  INVX1 U582 ( .A(n417), .Y(n419) );
  AND2X2 U583 ( .A(\state<0> ), .B(n343), .Y(n420) );
  INVX1 U584 ( .A(n420), .Y(n421) );
  OR2X2 U585 ( .A(\state<3> ), .B(\state<0> ), .Y(n422) );
  INVX1 U586 ( .A(n422), .Y(n423) );
  INVX1 U587 ( .A(n424), .Y(n425) );
  AND2X2 U588 ( .A(n432), .B(n314), .Y(n446) );
  AND2X2 U589 ( .A(\state<0> ), .B(\state<4> ), .Y(n426) );
  INVX1 U590 ( .A(n426), .Y(n427) );
  AND2X2 U591 ( .A(\state<4> ), .B(n693), .Y(n428) );
  INVX1 U592 ( .A(n428), .Y(n429) );
  AND2X2 U593 ( .A(\state<0> ), .B(n742), .Y(n430) );
  INVX1 U594 ( .A(n430), .Y(n431) );
  INVX1 U595 ( .A(n365), .Y(n705) );
  INVX1 U596 ( .A(n620), .Y(n432) );
  INVX1 U597 ( .A(n713), .Y(n434) );
  INVX4 U598 ( .A(n643), .Y(n713) );
  INVX1 U599 ( .A(n320), .Y(n435) );
  NOR2X1 U600 ( .A(\state<0> ), .B(n436), .Y(n438) );
  INVX1 U601 ( .A(n438), .Y(n437) );
  AND2X2 U602 ( .A(\state<2> ), .B(\state<3> ), .Y(n444) );
  AND2X2 U603 ( .A(n314), .B(n653), .Y(n439) );
  INVX1 U604 ( .A(n439), .Y(n440) );
  AND2X2 U605 ( .A(n300), .B(n713), .Y(n442) );
  AND2X2 U606 ( .A(\state<0> ), .B(n398), .Y(n443) );
  AND2X2 U607 ( .A(n712), .B(n398), .Y(n445) );
  INVX1 U608 ( .A(n735), .Y(n447) );
  INVX1 U609 ( .A(n370), .Y(n449) );
  OR2X2 U610 ( .A(n375), .B(n486), .Y(n450) );
  INVX1 U611 ( .A(n450), .Y(n451) );
  AND2X1 U612 ( .A(n463), .B(n461), .Y(n452) );
  INVX1 U613 ( .A(n452), .Y(n453) );
  AND2X1 U614 ( .A(n604), .B(n467), .Y(n454) );
  INVX1 U615 ( .A(n454), .Y(n455) );
  OR2X1 U616 ( .A(n577), .B(n458), .Y(n456) );
  INVX1 U617 ( .A(n456), .Y(n457) );
  OR2X1 U618 ( .A(n582), .B(n459), .Y(n458) );
  INVX1 U619 ( .A(n414), .Y(n459) );
  AND2X1 U620 ( .A(n464), .B(n538), .Y(n460) );
  INVX1 U621 ( .A(n460), .Y(n461) );
  AND2X1 U622 ( .A(n464), .B(n415), .Y(n462) );
  INVX1 U623 ( .A(n462), .Y(n463) );
  INVX1 U624 ( .A(n630), .Y(n464) );
  OR2X1 U625 ( .A(n506), .B(n466), .Y(n465) );
  OR2X1 U626 ( .A(n505), .B(n600), .Y(n466) );
  OR2X1 U627 ( .A(n533), .B(n469), .Y(n468) );
  OR2X1 U628 ( .A(n531), .B(n532), .Y(n469) );
  OR2X1 U629 ( .A(n489), .B(n473), .Y(n472) );
  OR2X1 U630 ( .A(n554), .B(n538), .Y(n473) );
  OR2X1 U631 ( .A(n485), .B(n477), .Y(n475) );
  INVX1 U632 ( .A(n475), .Y(n476) );
  OR2X1 U633 ( .A(n318), .B(n506), .Y(n477) );
  OR2X1 U634 ( .A(n567), .B(n479), .Y(n478) );
  OR2X1 U635 ( .A(n538), .B(n589), .Y(n479) );
  OR2X1 U636 ( .A(n492), .B(n481), .Y(n480) );
  OR2X1 U637 ( .A(n612), .B(n456), .Y(n481) );
  AND2X1 U638 ( .A(n572), .B(n484), .Y(n482) );
  INVX1 U639 ( .A(n484), .Y(n485) );
  INVX1 U640 ( .A(n486), .Y(n487) );
  OR2X1 U641 ( .A(n742), .B(n670), .Y(n489) );
  INVX1 U642 ( .A(n607), .Y(n670) );
  OR2X1 U643 ( .A(n574), .B(n584), .Y(n492) );
  INVX1 U644 ( .A(n367), .Y(n493) );
  INVX1 U645 ( .A(\nxtState<0> ), .Y(n494) );
  INVX1 U646 ( .A(n494), .Y(n495) );
  BUFX2 U647 ( .A(n684), .Y(n496) );
  BUFX2 U648 ( .A(n734), .Y(n497) );
  AND2X1 U649 ( .A(n666), .B(n675), .Y(n498) );
  INVX1 U650 ( .A(n498), .Y(n499) );
  INVX1 U651 ( .A(n370), .Y(n500) );
  INVX1 U652 ( .A(n502), .Y(n501) );
  AND2X2 U653 ( .A(n607), .B(n414), .Y(n503) );
  INVX1 U654 ( .A(n503), .Y(n504) );
  INVX1 U655 ( .A(n327), .Y(n505) );
  INVX1 U656 ( .A(n487), .Y(n506) );
  INVX1 U657 ( .A(n507), .Y(n508) );
  INVX1 U658 ( .A(n676), .Y(n509) );
  INVX1 U659 ( .A(n509), .Y(n510) );
  INVX1 U660 ( .A(n511), .Y(n512) );
  INVX1 U661 ( .A(n513), .Y(n514) );
  BUFX2 U662 ( .A(n645), .Y(n515) );
  INVX1 U663 ( .A(n516), .Y(n517) );
  OR2X2 U664 ( .A(n421), .B(n398), .Y(n518) );
  INVX1 U665 ( .A(n518), .Y(n519) );
  BUFX2 U666 ( .A(n649), .Y(n520) );
  INVX1 U667 ( .A(n678), .Y(n521) );
  INVX1 U668 ( .A(n521), .Y(n522) );
  INVX1 U669 ( .A(n690), .Y(n523) );
  INVX1 U670 ( .A(n523), .Y(n524) );
  OR2X1 U671 ( .A(n488), .B(n441), .Y(n525) );
  INVX1 U672 ( .A(n525), .Y(n526) );
  INVX1 U673 ( .A(n298), .Y(\DataOut<0> ) );
  INVX1 U674 ( .A(n297), .Y(\DataOut<10> ) );
  INVX1 U675 ( .A(n296), .Y(\DataOut<11> ) );
  INVX1 U676 ( .A(n295), .Y(\DataOut<12> ) );
  INVX1 U677 ( .A(n294), .Y(\DataOut<13> ) );
  INVX1 U678 ( .A(n293), .Y(\DataOut<14> ) );
  INVX1 U679 ( .A(n292), .Y(\DataOut<15> ) );
  INVX1 U680 ( .A(n291), .Y(\DataOut<1> ) );
  INVX1 U681 ( .A(n290), .Y(\DataOut<2> ) );
  INVX1 U682 ( .A(n289), .Y(\DataOut<3> ) );
  INVX1 U683 ( .A(n288), .Y(\DataOut<4> ) );
  INVX1 U684 ( .A(n287), .Y(\DataOut<5> ) );
  INVX1 U685 ( .A(n286), .Y(\DataOut<6> ) );
  INVX1 U686 ( .A(n285), .Y(\DataOut<7> ) );
  INVX1 U687 ( .A(n284), .Y(\DataOut<8> ) );
  INVX1 U688 ( .A(n283), .Y(\DataOut<9> ) );
  INVX1 U689 ( .A(waitMem_flop), .Y(n759) );
  BUFX2 U690 ( .A(n248), .Y(n527) );
  INVX1 U691 ( .A(n527), .Y(n760) );
  INVX1 U692 ( .A(n247), .Y(n761) );
  BUFX2 U693 ( .A(n246), .Y(n528) );
  INVX1 U694 ( .A(n528), .Y(n762) );
  BUFX2 U695 ( .A(n245), .Y(n529) );
  INVX1 U696 ( .A(n529), .Y(n763) );
  BUFX2 U697 ( .A(n242), .Y(n530) );
  INVX1 U698 ( .A(n530), .Y(n764) );
  INVX1 U699 ( .A(n431), .Y(n531) );
  INVX1 U700 ( .A(n490), .Y(n532) );
  INVX1 U701 ( .A(n608), .Y(n533) );
  AND2X1 U702 ( .A(n348), .B(n781), .Y(n534) );
  INVX1 U703 ( .A(n692), .Y(n535) );
  OR2X1 U704 ( .A(n650), .B(n589), .Y(n536) );
  INVX1 U705 ( .A(n536), .Y(n537) );
  INVX1 U706 ( .A(n448), .Y(n538) );
  OR2X1 U707 ( .A(n739), .B(n5), .Y(n539) );
  INVX1 U708 ( .A(n539), .Y(n540) );
  AND2X1 U709 ( .A(n484), .B(n601), .Y(n541) );
  INVX1 U710 ( .A(n541), .Y(n542) );
  OR2X1 U711 ( .A(n444), .B(n713), .Y(n543) );
  INVX1 U712 ( .A(n543), .Y(n544) );
  INVX1 U713 ( .A(n547), .Y(n545) );
  INVX1 U714 ( .A(n545), .Y(n546) );
  BUFX2 U715 ( .A(n579), .Y(n547) );
  BUFX2 U716 ( .A(n668), .Y(n548) );
  INVX1 U717 ( .A(n677), .Y(n549) );
  INVX1 U718 ( .A(n549), .Y(n550) );
  OR2X2 U719 ( .A(n366), .B(cacheHit), .Y(n551) );
  INVX1 U720 ( .A(n551), .Y(n552) );
  BUFX2 U721 ( .A(n656), .Y(n553) );
  INVX1 U722 ( .A(n555), .Y(n554) );
  BUFX2 U723 ( .A(n671), .Y(n555) );
  INVX1 U724 ( .A(n556), .Y(n557) );
  INVX1 U725 ( .A(n558), .Y(n559) );
  INVX1 U726 ( .A(n560), .Y(n561) );
  AND2X1 U727 ( .A(n607), .B(n604), .Y(n562) );
  INVX1 U728 ( .A(n562), .Y(n563) );
  AND2X1 U729 ( .A(\Addr<2> ), .B(\Addr<1> ), .Y(n564) );
  INVX1 U730 ( .A(n564), .Y(n565) );
  AND2X1 U731 ( .A(n476), .B(n608), .Y(n566) );
  INVX1 U732 ( .A(n566), .Y(n567) );
  INVX1 U733 ( .A(n569), .Y(n568) );
  AND2X1 U734 ( .A(n444), .B(n445), .Y(n570) );
  INVX1 U735 ( .A(n570), .Y(n571) );
  INVX1 U736 ( .A(n736), .Y(n572) );
  INVX1 U737 ( .A(n572), .Y(n573) );
  INVX1 U738 ( .A(n346), .Y(n574) );
  INVX1 U739 ( .A(n674), .Y(n575) );
  INVX1 U740 ( .A(n575), .Y(n576) );
  INVX1 U741 ( .A(n578), .Y(n577) );
  AOI21X1 U742 ( .A(n650), .B(n630), .C(n570), .Y(n579) );
  INVX1 U743 ( .A(n581), .Y(n580) );
  BUFX2 U744 ( .A(n192), .Y(n581) );
  AND2X1 U745 ( .A(n713), .B(n445), .Y(n582) );
  AND2X1 U746 ( .A(n603), .B(n593), .Y(n583) );
  INVX1 U747 ( .A(n583), .Y(n584) );
  INVX1 U748 ( .A(n374), .Y(n585) );
  INVX1 U749 ( .A(n374), .Y(n586) );
  INVX1 U750 ( .A(n230), .Y(n587) );
  INVX1 U751 ( .A(n588), .Y(n589) );
  INVX1 U752 ( .A(n269), .Y(n590) );
  INVX1 U753 ( .A(n590), .Y(n591) );
  INVX1 U754 ( .A(n590), .Y(n592) );
  INVX1 U755 ( .A(n500), .Y(n675) );
  INVX1 U756 ( .A(n594), .Y(n593) );
  INVX1 U757 ( .A(n703), .Y(n682) );
  INVX1 U758 ( .A(n595), .Y(n596) );
  AND2X1 U759 ( .A(n733), .B(n426), .Y(n597) );
  INVX1 U760 ( .A(n597), .Y(n598) );
  AND2X2 U761 ( .A(n366), .B(n449), .Y(n599) );
  INVX1 U762 ( .A(n600), .Y(n601) );
  INVX1 U763 ( .A(n366), .Y(n680) );
  INVX1 U764 ( .A(n602), .Y(n603) );
  INVX1 U765 ( .A(n605), .Y(n604) );
  INVX1 U766 ( .A(n606), .Y(n607) );
  INVX1 U767 ( .A(n706), .Y(n653) );
  INVX1 U768 ( .A(n375), .Y(n608) );
  INVX1 U769 ( .A(n384), .Y(n609) );
  INVX1 U770 ( .A(n384), .Y(n610) );
  BUFX2 U771 ( .A(\cacheOff<2> ), .Y(n611) );
  INVX1 U772 ( .A(n250), .Y(n612) );
  AND2X2 U773 ( .A(n392), .B(n707), .Y(n613) );
  INVX1 U774 ( .A(n613), .Y(n614) );
  INVX1 U775 ( .A(n615), .Y(n616) );
  INVX1 U776 ( .A(n617), .Y(n618) );
  INVX1 U777 ( .A(n634), .Y(n632) );
  INVX1 U778 ( .A(n717), .Y(n619) );
  INVX1 U779 ( .A(n636), .Y(n635) );
  INVX1 U780 ( .A(n699), .Y(n733) );
  NAND2X1 U781 ( .A(n712), .B(n700), .Y(n621) );
  NAND2X1 U782 ( .A(\state<0> ), .B(n699), .Y(n622) );
  INVX1 U783 ( .A(\state<0> ), .Y(n620) );
  INVX1 U784 ( .A(n729), .Y(n623) );
  INVX1 U785 ( .A(n730), .Y(n624) );
  INVX1 U786 ( .A(n731), .Y(n625) );
  INVX1 U787 ( .A(n732), .Y(n626) );
  INVX1 U788 ( .A(\state<3> ), .Y(n695) );
  INVX1 U789 ( .A(\cacheDataOut<14> ), .Y(n718) );
  INVX1 U790 ( .A(\cacheDataOut<12> ), .Y(n720) );
  INVX1 U791 ( .A(\cacheDataOut<10> ), .Y(n722) );
  INVX1 U792 ( .A(\cacheDataOut<8> ), .Y(n724) );
  INVX1 U793 ( .A(\cacheDataOut<15> ), .Y(n717) );
  INVX1 U794 ( .A(\cacheDataOut<13> ), .Y(n719) );
  INVX1 U795 ( .A(\cacheDataOut<11> ), .Y(n721) );
  INVX1 U796 ( .A(\cacheDataOut<9> ), .Y(n723) );
  INVX1 U797 ( .A(\cacheDataOut<7> ), .Y(n725) );
  INVX1 U798 ( .A(\cacheDataOut<6> ), .Y(n726) );
  INVX1 U799 ( .A(\cacheDataOut<5> ), .Y(n727) );
  INVX1 U800 ( .A(\cacheDataOut<4> ), .Y(n728) );
  INVX1 U801 ( .A(\cacheDataOut<3> ), .Y(n729) );
  INVX1 U802 ( .A(\cacheDataOut<2> ), .Y(n730) );
  INVX1 U803 ( .A(\cacheDataOut<1> ), .Y(n731) );
  INVX1 U804 ( .A(\cacheDataOut<0> ), .Y(n732) );
  BUFX4 U805 ( .A(memStall), .Y(n630) );
  INVX8 U806 ( .A(n634), .Y(n633) );
  INVX8 U807 ( .A(n638), .Y(n637) );
  INVX8 U808 ( .A(n640), .Y(n639) );
  INVX8 U809 ( .A(n642), .Y(n641) );
  NAND2X1 U810 ( .A(n300), .B(n320), .Y(n699) );
  OR2X2 U811 ( .A(\state<3> ), .B(\state<2> ), .Y(n643) );
  OAI21X1 U812 ( .A(cacheHit), .B(valid), .C(n330), .Y(n666) );
  AOI21X1 U813 ( .A(n537), .B(n305), .C(n630), .Y(n645) );
  AOI21X1 U814 ( .A(n680), .B(n666), .C(n515), .Y(n649) );
  AND2X2 U815 ( .A(\state<4> ), .B(n300), .Y(n646) );
  NAND3X1 U816 ( .A(n620), .B(n713), .C(n646), .Y(n703) );
  NAND2X1 U817 ( .A(\nxtEvict<4> ), .B(n682), .Y(n648) );
  NAND3X1 U818 ( .A(n426), .B(n713), .C(n693), .Y(n735) );
  NOR3X1 U819 ( .A(n411), .B(n538), .C(n475), .Y(n647) );
  NAND3X1 U820 ( .A(n648), .B(n520), .C(n647), .Y(\nxtState<4> ) );
  NAND3X1 U821 ( .A(valid), .B(n552), .C(dirty), .Y(n651) );
  NAND3X1 U822 ( .A(n716), .B(n321), .C(n620), .Y(n706) );
  NOR2X1 U823 ( .A(n703), .B(n654), .Y(n655) );
  AOI21X1 U824 ( .A(n630), .B(n742), .C(n655), .Y(n656) );
  NOR3X1 U825 ( .A(n459), .B(n670), .C(n379), .Y(n669) );
  OAI21X1 U826 ( .A(n663), .B(\wait4Cycles_flop<0> ), .C(n657), .Y(n683) );
  NOR3X1 U827 ( .A(n565), .B(n683), .C(n327), .Y(n658) );
  AOI21X1 U828 ( .A(n580), .B(n409), .C(n658), .Y(n668) );
  NAND2X1 U829 ( .A(\nxtEvict<2> ), .B(n682), .Y(n660) );
  MUX2X1 U830 ( .B(n605), .A(n542), .S(n630), .Y(n659) );
  AOI21X1 U831 ( .A(n741), .B(n661), .C(n630), .Y(n674) );
  NOR2X1 U832 ( .A(n630), .B(\wait4Cycles_flop<0> ), .Y(n664) );
  NOR3X1 U833 ( .A(n681), .B(n403), .C(n405), .Y(n667) );
  NAND3X1 U834 ( .A(n669), .B(n548), .C(n667), .Y(\nxtState<2> ) );
  NAND2X1 U835 ( .A(\nxtEvict<1> ), .B(n682), .Y(n673) );
  AOI21X1 U836 ( .A(n581), .B(n409), .C(n594), .Y(n671) );
  MUX2X1 U837 ( .B(n472), .A(n605), .S(n630), .Y(n672) );
  AOI21X1 U838 ( .A(n576), .B(n318), .C(n383), .Y(n678) );
  AOI21X1 U839 ( .A(n675), .B(n609), .C(n582), .Y(n677) );
  NAND3X1 U840 ( .A(n440), .B(n546), .C(n608), .Y(n676) );
  NAND3X1 U841 ( .A(n522), .B(n550), .C(n557), .Y(\nxtState<1> ) );
  AOI21X1 U842 ( .A(n680), .B(n609), .C(n517), .Y(n690) );
  AOI21X1 U843 ( .A(\nxtEvict<0> ), .B(n682), .C(n681), .Y(n689) );
  NAND3X1 U844 ( .A(n506), .B(n741), .C(n534), .Y(n684) );
  AND2X2 U845 ( .A(n601), .B(n604), .Y(n685) );
  NAND3X1 U846 ( .A(n431), .B(n685), .C(n607), .Y(n736) );
  NOR3X1 U847 ( .A(n506), .B(n573), .C(n584), .Y(n686) );
  MUX2X1 U848 ( .B(n457), .A(n686), .S(n630), .Y(n687) );
  NOR3X1 U849 ( .A(n561), .B(n687), .C(n439), .Y(n688) );
  NAND3X1 U850 ( .A(n524), .B(n689), .C(n688), .Y(\nxtState<0> ) );
  OAI21X1 U851 ( .A(n609), .B(n333), .C(n691), .Y(doneWait_in) );
  OAI21X1 U852 ( .A(Wr), .B(Rd), .C(n339), .Y(n692) );
  AOI21X1 U853 ( .A(n620), .B(n470), .C(n442), .Y(n697) );
  NAND3X1 U854 ( .A(\state<0> ), .B(n693), .C(n610), .Y(n694) );
  AND2X2 U855 ( .A(n585), .B(n706), .Y(n702) );
  NAND2X1 U856 ( .A(\state<3> ), .B(n345), .Y(n700) );
  AOI21X1 U857 ( .A(\state<4> ), .B(n343), .C(n373), .Y(n701) );
  AND2X2 U858 ( .A(n366), .B(n703), .Y(n704) );
  NAND3X1 U859 ( .A(n448), .B(n346), .C(n451), .Y(n269) );
  AOI21X1 U860 ( .A(\Addr<1> ), .B(n591), .C(n455), .Y(n708) );
  AOI21X1 U861 ( .A(n340), .B(n445), .C(n519), .Y(n707) );
  NAND3X1 U862 ( .A(n397), .B(n526), .C(n559), .Y(\cacheOff<2> ) );
  MUX2X1 U863 ( .B(n716), .A(n428), .S(n423), .Y(n711) );
  MUX2X1 U864 ( .B(n343), .A(n304), .S(n398), .Y(n710) );
  NAND3X1 U865 ( .A(n484), .B(n608), .C(n323), .Y(\nextEvictState_in<0> ) );
  AOI21X1 U866 ( .A(\state<0> ), .B(n355), .C(n344), .Y(n714) );
  MUX2X1 U867 ( .B(n714), .A(n544), .S(n314), .Y(n715) );
  MUX2X1 U868 ( .B(n718), .A(n783), .S(n538), .Y(\memDataIn<14> ) );
  MUX2X1 U869 ( .B(n719), .A(n784), .S(n538), .Y(\memDataIn<13> ) );
  MUX2X1 U870 ( .B(n720), .A(n785), .S(n538), .Y(\memDataIn<12> ) );
  MUX2X1 U871 ( .B(n721), .A(n786), .S(n538), .Y(\memDataIn<11> ) );
  MUX2X1 U872 ( .B(n722), .A(n787), .S(n538), .Y(\memDataIn<10> ) );
  MUX2X1 U873 ( .B(n723), .A(n788), .S(n538), .Y(\memDataIn<9> ) );
  MUX2X1 U874 ( .B(n725), .A(n790), .S(n538), .Y(\memDataIn<7> ) );
  MUX2X1 U875 ( .B(n728), .A(n793), .S(n538), .Y(\memDataIn<4> ) );
  MUX2X1 U876 ( .B(n337), .A(n794), .S(n538), .Y(\memDataIn<3> ) );
  MUX2X1 U877 ( .B(n338), .A(n795), .S(n538), .Y(\memDataIn<2> ) );
  MUX2X1 U878 ( .B(n313), .A(n796), .S(n538), .Y(\memDataIn<1> ) );
  AOI21X1 U879 ( .A(n733), .B(n427), .C(n483), .Y(n734) );
  NOR3X1 U880 ( .A(n563), .B(n597), .C(n439), .Y(n250) );
  NOR2X1 U881 ( .A(n329), .B(n446), .Y(n737) );
  MUX2X1 U882 ( .B(n435), .A(n324), .S(n737), .Y(n738) );
  MUX2X1 U883 ( .B(n344), .A(n321), .S(n425), .Y(n11) );
  XNOR2X1 U884 ( .A(n329), .B(n340), .Y(n739) );
  MUX2X1 U885 ( .B(n540), .A(n344), .S(n446), .Y(n9) );
endmodule

